module memory(clk,reset,address,data_in,data_out,rwn,start,ready,address_test1,address_test2,address_test3,data_test1,data_test2,data_test3);
input clk,reset,start,rwn;
input [15:0] address,address_test1,address_test2,address_test3;
output [15:0] data_test1,data_test2,data_test3;
output ready;
input [15:0] data_in;
output reg [15:0] data_out;
reg [15:0] array[65535:0],data_t;
reg state;
reg [15:0] ad_t;
reg [1:0] counter;
reg rwn_t;
assign ready=~state;
assign data_test1=array[address_test1];
assign data_test2=array[address_test2];
assign data_test3=array[address_test3];
always @(posedge clk or posedge reset)
begin
if(reset)
begin
array[0] <= 16'b0000_0000_0000_0000;
array[1] <= 16'b0000_0000_0000_0000;
array[2] <= 16'b0000_0000_0000_0000;
array[3] <= 16'b0000_0000_0000_0000;
array[4] <= 16'b0000_0000_0000_0000;
array[5] <= 16'b0000_0000_0000_0000;
array[6] <= 16'b0000_0000_0000_0000;
array[7] <= 16'b0000_0000_0000_0000;
array[8] <= 16'b0000_0000_0000_0000;
array[9] <= 16'b0000_0000_0000_0000;
array[10] <= 16'b0000_0000_0000_0000;
array[11] <= 16'b0000_0000_0000_0000;
array[12] <= 16'b0000_0000_0000_0000;
array[13] <= 16'b0000_0000_0000_0000;
array[14] <= 16'b0000_0000_0000_0000;
array[15] <= 16'b0000_0000_0000_0000;
array[16] <= 16'b0000_0000_0000_0000;
array[17] <= 16'b0000_0000_0000_0000;
array[18] <= 16'b0000_0000_0000_0000;
array[19] <= 16'b0000_0000_0000_0000;
array[20] <= 16'b0000_0000_0000_0000;
array[21] <= 16'b0000_0000_0000_0000;
array[22] <= 16'b0000_0000_0000_0000;
array[23] <= 16'b0000_0000_0000_0000;
array[24] <= 16'b0000_0000_0000_0000;
array[25] <= 16'b0000_0000_0000_0000;
array[26] <= 16'b0000_0000_0000_0000;
array[27] <= 16'b0000_0000_0000_0000;
array[28] <= 16'b0000_0000_0000_0000;
array[29] <= 16'b0000_0000_0000_0000;
array[30] <= 16'b0000_0000_0000_0000;
array[31] <= 16'b0000_0000_0000_0000;
array[32] <= 16'b0000_0000_0000_0000;
array[33] <= 16'b0000_0000_0000_0000;
array[34] <= 16'b0000_0000_0000_0000;
array[35] <= 16'b0000_0000_0000_0000;
array[36] <= 16'b0000_0000_0000_0000;
array[37] <= 16'b0000_0000_0000_0000;
array[38] <= 16'b0000_0000_0000_0000;
array[39] <= 16'b0000_0000_0000_0000;
array[40] <= 16'b0000_0000_0000_0000;
array[41] <= 16'b0000_0000_0000_0000;
array[42] <= 16'b0000_0000_0000_0000;
array[43] <= 16'b0000_0000_0000_0000;
array[44] <= 16'b0000_0000_0000_0000;
array[45] <= 16'b0000_0000_0000_0000;
array[46] <= 16'b0000_0000_0000_0000;
array[47] <= 16'b0000_0000_0000_0000;
array[48] <= 16'b0000_0000_0000_0000;
array[49] <= 16'b0000_0000_0000_0000;
array[50] <= 16'b0000_0000_0000_0000;
array[51] <= 16'b0000_0000_0000_0000;
array[52] <= 16'b0000_0000_0000_0000;
array[53] <= 16'b0000_0000_0000_0000;
array[54] <= 16'b0000_0000_0000_0000;
array[55] <= 16'b0000_0000_0000_0000;
array[56] <= 16'b0000_0000_0000_0000;
array[57] <= 16'b0000_0000_0000_0000;
array[58] <= 16'b0000_0000_0000_0000;
array[59] <= 16'b0000_0000_0000_0000;
array[60] <= 16'b0000_0000_0000_0000;
array[61] <= 16'b0000_0000_0000_0000;
array[62] <= 16'b0000_0000_0000_0000;
array[63] <= 16'b0000_0000_0000_0000;
array[64] <= 16'b0000_0000_0000_0000;
array[65] <= 16'b0000_0000_0000_0000;
array[66] <= 16'b0000_0000_0000_0000;
array[67] <= 16'b0000_0000_0000_0000;
array[68] <= 16'b0000_0000_0000_0000;
array[69] <= 16'b0000_0000_0000_0000;
array[70] <= 16'b0000_0000_0000_0000;
array[71] <= 16'b0000_0000_0000_0000;
array[72] <= 16'b0000_0000_0000_0000;
array[73] <= 16'b0000_0000_0000_0000;
array[74] <= 16'b0000_0000_0000_0000;
array[75] <= 16'b0000_0000_0000_0000;
array[76] <= 16'b0000_0000_0000_0000;
array[77] <= 16'b0000_0000_0000_0000;
array[78] <= 16'b0000_0000_0000_0000;
array[79] <= 16'b0000_0000_0000_0000;
array[80] <= 16'b0000_0000_0000_0000;
array[81] <= 16'b0000_0000_0000_0000;
array[82] <= 16'b0000_0000_0000_0000;
array[83] <= 16'b0000_0000_0000_0000;
array[84] <= 16'b0000_0000_0000_0000;
array[85] <= 16'b0000_0000_0000_0000;
array[86] <= 16'b0000_0000_0000_0000;
array[87] <= 16'b0000_0000_0000_0000;
array[88] <= 16'b0000_0000_0000_0000;
array[89] <= 16'b0000_0000_0000_0000;
array[90] <= 16'b0000_0000_0000_0000;
array[91] <= 16'b0000_0000_0000_0000;
array[92] <= 16'b0000_0000_0000_0000;
array[93] <= 16'b0000_0000_0000_0000;
array[94] <= 16'b0000_0000_0000_0000;
array[95] <= 16'b0000_0000_0000_0000;
array[96] <= 16'b0000_0000_0000_0000;
array[97] <= 16'b0000_0000_0000_0000;
array[98] <= 16'b0000_0000_0000_0000;
array[99] <= 16'b0000_0000_0000_0000;
array[100] <= 16'b0000_0000_0000_0000;
array[101] <= 16'b0000_0000_0000_0000;
array[102] <= 16'b0000_0000_0000_0000;
array[103] <= 16'b0000_0000_0000_0000;
array[104] <= 16'b0000_0000_0000_0000;
array[105] <= 16'b0000_0000_0000_0000;
array[106] <= 16'b0000_0000_0000_0000;
array[107] <= 16'b0000_0000_0000_0000;
array[108] <= 16'b0000_0000_0000_0000;
array[109] <= 16'b0000_0000_0000_0000;
array[110] <= 16'b0000_0000_0000_0000;
array[111] <= 16'b0000_0000_0000_0000;
array[112] <= 16'b0000_0000_0000_0000;
array[113] <= 16'b0000_0000_0000_0000;
array[114] <= 16'b0000_0000_0000_0000;
array[115] <= 16'b0000_0000_0000_0000;
array[116] <= 16'b0000_0000_0000_0000;
array[117] <= 16'b0000_0000_0000_0000;
array[118] <= 16'b0000_0000_0000_0000;
array[119] <= 16'b0000_0000_0000_0000;
array[120] <= 16'b0000_0000_0000_0000;
array[121] <= 16'b0000_0000_0000_0000;
array[122] <= 16'b0000_0000_0000_0000;
array[123] <= 16'b0000_0000_0000_0000;
array[124] <= 16'b0000_0000_0000_0000;
array[125] <= 16'b0000_0000_0000_0000;
array[126] <= 16'b0000_0000_0000_0000;
array[127] <= 16'b0000_0000_0000_0000;
array[128] <= 16'b0000_0000_0000_0000;
array[129] <= 16'b0000_0000_0000_0000;
array[130] <= 16'b0000_0000_0000_0000;
array[131] <= 16'b0000_0000_0000_0000;
array[132] <= 16'b0000_0000_0000_0000;
array[133] <= 16'b0000_0000_0000_0000;
array[134] <= 16'b0000_0000_0000_0000;
array[135] <= 16'b0000_0000_0000_0000;
array[136] <= 16'b0000_0000_0000_0000;
array[137] <= 16'b0000_0000_0000_0000;
array[138] <= 16'b0000_0000_0000_0000;
array[139] <= 16'b0000_0000_0000_0000;
array[140] <= 16'b0000_0000_0000_0000;
array[141] <= 16'b0000_0000_0000_0000;
array[142] <= 16'b0000_0000_0000_0000;
array[143] <= 16'b0000_0000_0000_0000;
array[144] <= 16'b0000_0000_0000_0000;
array[145] <= 16'b0000_0000_0000_0000;
array[146] <= 16'b0000_0000_0000_0000;
array[147] <= 16'b0000_0000_0000_0000;
array[148] <= 16'b0000_0000_0000_0000;
array[149] <= 16'b0000_0000_0000_0000;
array[150] <= 16'b0000_0000_0000_0000;
array[151] <= 16'b0000_0000_0000_0000;
array[152] <= 16'b0000_0000_0000_0000;
array[153] <= 16'b0000_0000_0000_0000;
array[154] <= 16'b0000_0000_0000_0000;
array[155] <= 16'b0000_0000_0000_0000;
array[156] <= 16'b0000_0000_0000_0000;
array[157] <= 16'b0000_0000_0000_0000;
array[158] <= 16'b0000_0000_0000_0000;
array[159] <= 16'b0000_0000_0000_0000;
array[160] <= 16'b0000_0000_0000_0000;
array[161] <= 16'b0000_0000_0000_0000;
array[162] <= 16'b0000_0000_0000_0000;
array[163] <= 16'b0000_0000_0000_0000;
array[164] <= 16'b0000_0000_0000_0000;
array[165] <= 16'b0000_0000_0000_0000;
array[166] <= 16'b0000_0000_0000_0000;
array[167] <= 16'b0000_0000_0000_0000;
array[168] <= 16'b0000_0000_0000_0000;
array[169] <= 16'b0000_0000_0000_0000;
array[170] <= 16'b0000_0000_0000_0000;
array[171] <= 16'b0000_0000_0000_0000;
array[172] <= 16'b0000_0000_0000_0000;
array[173] <= 16'b0000_0000_0000_0000;
array[174] <= 16'b0000_0000_0000_0000;
array[175] <= 16'b0000_0000_0000_0000;
array[176] <= 16'b0000_0000_0000_0000;
array[177] <= 16'b0000_0000_0000_0000;
array[178] <= 16'b0000_0000_0000_0000;
array[179] <= 16'b0000_0000_0000_0000;
array[180] <= 16'b0000_0000_0000_0000;
array[181] <= 16'b0000_0000_0000_0000;
array[182] <= 16'b0000_0000_0000_0000;
array[183] <= 16'b0000_0000_0000_0000;
array[184] <= 16'b0000_0000_0000_0000;
array[185] <= 16'b0000_0000_0000_0000;
array[186] <= 16'b0000_0000_0000_0000;
array[187] <= 16'b0000_0000_0000_0000;
array[188] <= 16'b0000_0000_0000_0000;
array[189] <= 16'b0000_0000_0000_0000;
array[190] <= 16'b0000_0000_0000_0000;
array[191] <= 16'b0000_0000_0000_0000;
array[192] <= 16'b0000_0000_0000_0000;
array[193] <= 16'b0000_0000_0000_0000;
array[194] <= 16'b0000_0000_0000_0000;
array[195] <= 16'b0000_0000_0000_0000;
array[196] <= 16'b0000_0000_0000_0000;
array[197] <= 16'b0000_0000_0000_0000;
array[198] <= 16'b0000_0000_0000_0000;
array[199] <= 16'b0000_0000_0000_0000;
array[200] <= 16'b0000_0000_0000_0000;
array[201] <= 16'b0000_0000_0000_0000;
array[202] <= 16'b0000_0000_0000_0000;
array[203] <= 16'b0000_0000_0000_0000;
array[204] <= 16'b0000_0000_0000_0000;
array[205] <= 16'b0000_0000_0000_0000;
array[206] <= 16'b0000_0000_0000_0000;
array[207] <= 16'b0000_0000_0000_0000;
array[208] <= 16'b0000_0000_0000_0000;
array[209] <= 16'b0000_0000_0000_0000;
array[210] <= 16'b0000_0000_0000_0000;
array[211] <= 16'b0000_0000_0000_0000;
array[212] <= 16'b0000_0000_0000_0000;
array[213] <= 16'b0000_0000_0000_0000;
array[214] <= 16'b0000_0000_0000_0000;
array[215] <= 16'b0000_0000_0000_0000;
array[216] <= 16'b0000_0000_0000_0000;
array[217] <= 16'b0000_0000_0000_0000;
array[218] <= 16'b0000_0000_0000_0000;
array[219] <= 16'b0000_0000_0000_0000;
array[220] <= 16'b0000_0000_0000_0000;
array[221] <= 16'b0000_0000_0000_0000;
array[222] <= 16'b0000_0000_0000_0000;
array[223] <= 16'b0000_0000_0000_0000;
array[224] <= 16'b0000_0000_0000_0000;
array[225] <= 16'b0000_0000_0000_0000;
array[226] <= 16'b0000_0000_0000_0000;
array[227] <= 16'b0000_0000_0000_0000;
array[228] <= 16'b0000_0000_0000_0000;
array[229] <= 16'b0000_0000_0000_0000;
array[230] <= 16'b0000_0000_0000_0000;
array[231] <= 16'b0000_0000_0000_0000;
array[232] <= 16'b0000_0000_0000_0000;
array[233] <= 16'b0000_0000_0000_0000;
array[234] <= 16'b0000_0000_0000_0000;
array[235] <= 16'b0000_0000_0000_0000;
array[236] <= 16'b0000_0000_0000_0000;
array[237] <= 16'b0000_0000_0000_0000;
array[238] <= 16'b0000_0000_0000_0000;
array[239] <= 16'b0000_0000_0000_0000;
array[240] <= 16'b0000_0000_0000_0000;
array[241] <= 16'b0000_0000_0000_0000;
array[242] <= 16'b0000_0000_0000_0000;
array[243] <= 16'b0000_0000_0000_0000;
array[244] <= 16'b0000_0000_0000_0000;
array[245] <= 16'b0000_0000_0000_0000;
array[246] <= 16'b0000_0000_0000_0000;
array[247] <= 16'b0000_0000_0000_0000;
array[248] <= 16'b0000_0000_0000_0000;
array[249] <= 16'b0000_0000_0000_0000;
array[250] <= 16'b0000_0000_0000_0000;
array[251] <= 16'b0000_0000_0000_0000;
array[252] <= 16'b0000_0000_0000_0000;
array[253] <= 16'b0000_0000_0000_0000;
array[254] <= 16'b0000_0000_0000_0000;
array[255] <= 16'b0000_0000_0000_0000;
array[256] <= 16'b0000_0000_0000_0000;
array[257] <= 16'b0000_0000_0000_0000;
array[258] <= 16'b0000_0000_0000_0000;
array[259] <= 16'b0000_0000_0000_0000;
array[260] <= 16'b0000_0000_0000_0000;
array[261] <= 16'b0000_0000_0000_0000;
array[262] <= 16'b0000_0000_0000_0000;
array[263] <= 16'b0000_0000_0000_0000;
array[264] <= 16'b0000_0000_0000_0000;
array[265] <= 16'b0000_0000_0000_0000;
array[266] <= 16'b0000_0000_0000_0000;
array[267] <= 16'b0000_0000_0000_0000;
array[268] <= 16'b0000_0000_0000_0000;
array[269] <= 16'b0000_0000_0000_0000;
array[270] <= 16'b0000_0000_0000_0000;
array[271] <= 16'b0000_0000_0000_0000;
array[272] <= 16'b0000_0000_0000_0000;
array[273] <= 16'b0000_0000_0000_0000;
array[274] <= 16'b0000_0000_0000_0000;
array[275] <= 16'b0000_0000_0000_0000;
array[276] <= 16'b0000_0000_0000_0000;
array[277] <= 16'b0000_0000_0000_0000;
array[278] <= 16'b0000_0000_0000_0000;
array[279] <= 16'b0000_0000_0000_0000;
array[280] <= 16'b0000_0000_0000_0000;
array[281] <= 16'b0000_0000_0000_0000;
array[282] <= 16'b0000_0000_0000_0000;
array[283] <= 16'b0000_0000_0000_0000;
array[284] <= 16'b0000_0000_0000_0000;
array[285] <= 16'b0000_0000_0000_0000;
array[286] <= 16'b0000_0000_0000_0000;
array[287] <= 16'b0000_0000_0000_0000;
array[288] <= 16'b0000_0000_0000_0000;
array[289] <= 16'b0000_0000_0000_0000;
array[290] <= 16'b0000_0000_0000_0000;
array[291] <= 16'b0000_0000_0000_0000;
array[292] <= 16'b0000_0000_0000_0000;
array[293] <= 16'b0000_0000_0000_0000;
array[294] <= 16'b0000_0000_0000_0000;
array[295] <= 16'b0000_0000_0000_0000;
array[296] <= 16'b0000_0000_0000_0000;
array[297] <= 16'b0000_0000_0000_0000;
array[298] <= 16'b0000_0000_0000_0000;
array[299] <= 16'b0000_0000_0000_0000;
array[300] <= 16'b0000_0000_0000_0000;
array[301] <= 16'b0000_0000_0000_0000;
array[302] <= 16'b0000_0000_0000_0000;
array[303] <= 16'b0000_0000_0000_0000;
array[304] <= 16'b0000_0000_0000_0000;
array[305] <= 16'b0000_0000_0000_0000;
array[306] <= 16'b0000_0000_0000_0000;
array[307] <= 16'b0000_0000_0000_0000;
array[308] <= 16'b0000_0000_0000_0000;
array[309] <= 16'b0000_0000_0000_0000;
array[310] <= 16'b0000_0000_0000_0000;
array[311] <= 16'b0000_0000_0000_0000;
array[312] <= 16'b0000_0000_0000_0000;
array[313] <= 16'b0000_0000_0000_0000;
array[314] <= 16'b0000_0000_0000_0000;
array[315] <= 16'b0000_0000_0000_0000;
array[316] <= 16'b0000_0000_0000_0000;
array[317] <= 16'b0000_0000_0000_0000;
array[318] <= 16'b0000_0000_0000_0000;
array[319] <= 16'b0000_0000_0000_0000;
array[320] <= 16'b0000_0000_0000_0000;
array[321] <= 16'b0000_0000_0000_0000;
array[322] <= 16'b0000_0000_0000_0000;
array[323] <= 16'b0000_0000_0000_0000;
array[324] <= 16'b0000_0000_0000_0000;
array[325] <= 16'b0000_0000_0000_0000;
array[326] <= 16'b0000_0000_0000_0000;
array[327] <= 16'b0000_0000_0000_0000;
array[328] <= 16'b0000_0000_0000_0000;
array[329] <= 16'b0000_0000_0000_0000;
array[330] <= 16'b0000_0000_0000_0000;
array[331] <= 16'b0000_0000_0000_0000;
array[332] <= 16'b0000_0000_0000_0000;
array[333] <= 16'b0000_0000_0000_0000;
array[334] <= 16'b0000_0000_0000_0000;
array[335] <= 16'b0000_0000_0000_0000;
array[336] <= 16'b0000_0000_0000_0000;
array[337] <= 16'b0000_0000_0000_0000;
array[338] <= 16'b0000_0000_0000_0000;
array[339] <= 16'b0000_0000_0000_0000;
array[340] <= 16'b0000_0000_0000_0000;
array[341] <= 16'b0000_0000_0000_0000;
array[342] <= 16'b0000_0000_0000_0000;
array[343] <= 16'b0000_0000_0000_0000;
array[344] <= 16'b0000_0000_0000_0000;
array[345] <= 16'b0000_0000_0000_0000;
array[346] <= 16'b0000_0000_0000_0000;
array[347] <= 16'b0000_0000_0000_0000;
array[348] <= 16'b0000_0000_0000_0000;
array[349] <= 16'b0000_0000_0000_0000;
array[350] <= 16'b0000_0000_0000_0000;
array[351] <= 16'b0000_0000_0000_0000;
array[352] <= 16'b0000_0000_0000_0000;
array[353] <= 16'b0000_0000_0000_0000;
array[354] <= 16'b0000_0000_0000_0000;
array[355] <= 16'b0000_0000_0000_0000;
array[356] <= 16'b0000_0000_0000_0000;
array[357] <= 16'b0000_0000_0000_0000;
array[358] <= 16'b0000_0000_0000_0000;
array[359] <= 16'b0000_0000_0000_0000;
array[360] <= 16'b0000_0000_0000_0000;
array[361] <= 16'b0000_0000_0000_0000;
array[362] <= 16'b0000_0000_0000_0000;
array[363] <= 16'b0000_0000_0000_0000;
array[364] <= 16'b0000_0000_0000_0000;
array[365] <= 16'b0000_0000_0000_0000;
array[366] <= 16'b0000_0000_0000_0000;
array[367] <= 16'b0000_0000_0000_0000;
array[368] <= 16'b0000_0000_0000_0000;
array[369] <= 16'b0000_0000_0000_0000;
array[370] <= 16'b0000_0000_0000_0000;
array[371] <= 16'b0000_0000_0000_0000;
array[372] <= 16'b0000_0000_0000_0000;
array[373] <= 16'b0000_0000_0000_0000;
array[374] <= 16'b0000_0000_0000_0000;
array[375] <= 16'b0000_0000_0000_0000;
array[376] <= 16'b0000_0000_0000_0000;
array[377] <= 16'b0000_0000_0000_0000;
array[378] <= 16'b0000_0000_0000_0000;
array[379] <= 16'b0000_0000_0000_0000;
array[380] <= 16'b0000_0000_0000_0000;
array[381] <= 16'b0000_0000_0000_0000;
array[382] <= 16'b0000_0000_0000_0000;
array[383] <= 16'b0000_0000_0000_0000;
array[384] <= 16'b0000_0000_0000_0000;
array[385] <= 16'b0000_0000_0000_0000;
array[386] <= 16'b0000_0000_0000_0000;
array[387] <= 16'b0000_0000_0000_0000;
array[388] <= 16'b0000_0000_0000_0000;
array[389] <= 16'b0000_0000_0000_0000;
array[390] <= 16'b0000_0000_0000_0000;
array[391] <= 16'b0000_0000_0000_0000;
array[392] <= 16'b0000_0000_0000_0000;
array[393] <= 16'b0000_0000_0000_0000;
array[394] <= 16'b0000_0000_0000_0000;
array[395] <= 16'b0000_0000_0000_0000;
array[396] <= 16'b0000_0000_0000_0000;
array[397] <= 16'b0000_0000_0000_0000;
array[398] <= 16'b0000_0000_0000_0000;
array[399] <= 16'b0000_0000_0000_0000;
array[400] <= 16'b0000_0000_0000_0000;
array[401] <= 16'b0000_0000_0000_0000;
array[402] <= 16'b0000_0000_0000_0000;
array[403] <= 16'b0000_0000_0000_0000;
array[404] <= 16'b0000_0000_0000_0000;
array[405] <= 16'b0000_0000_0000_0000;
array[406] <= 16'b0000_0000_0000_0000;
array[407] <= 16'b0000_0000_0000_0000;
array[408] <= 16'b0000_0000_0000_0000;
array[409] <= 16'b0000_0000_0000_0000;
array[410] <= 16'b0000_0000_0000_0000;
array[411] <= 16'b0000_0000_0000_0000;
array[412] <= 16'b0000_0000_0000_0000;
array[413] <= 16'b0000_0000_0000_0000;
array[414] <= 16'b0000_0000_0000_0000;
array[415] <= 16'b0000_0000_0000_0000;
array[416] <= 16'b0000_0000_0000_0000;
array[417] <= 16'b0000_0000_0000_0000;
array[418] <= 16'b0000_0000_0000_0000;
array[419] <= 16'b0000_0000_0000_0000;
array[420] <= 16'b0000_0000_0000_0000;
array[421] <= 16'b0000_0000_0000_0000;
array[422] <= 16'b0000_0000_0000_0000;
array[423] <= 16'b0000_0000_0000_0000;
array[424] <= 16'b0000_0000_0000_0000;
array[425] <= 16'b0000_0000_0000_0000;
array[426] <= 16'b0000_0000_0000_0000;
array[427] <= 16'b0000_0000_0000_0000;
array[428] <= 16'b0000_0000_0000_0000;
array[429] <= 16'b0000_0000_0000_0000;
array[430] <= 16'b0000_0000_0000_0000;
array[431] <= 16'b0000_0000_0000_0000;
array[432] <= 16'b0000_0000_0000_0000;
array[433] <= 16'b0000_0000_0000_0000;
array[434] <= 16'b0000_0000_0000_0000;
array[435] <= 16'b0000_0000_0000_0000;
array[436] <= 16'b0000_0000_0000_0000;
array[437] <= 16'b0000_0000_0000_0000;
array[438] <= 16'b0000_0000_0000_0000;
array[439] <= 16'b0000_0000_0000_0000;
array[440] <= 16'b0000_0000_0000_0000;
array[441] <= 16'b0000_0000_0000_0000;
array[442] <= 16'b0000_0000_0000_0000;
array[443] <= 16'b0000_0000_0000_0000;
array[444] <= 16'b0000_0000_0000_0000;
array[445] <= 16'b0000_0000_0000_0000;
array[446] <= 16'b0000_0000_0000_0000;
array[447] <= 16'b0000_0000_0000_0000;
array[448] <= 16'b0000_0000_0000_0000;
array[449] <= 16'b0000_0000_0000_0000;
array[450] <= 16'b0000_0000_0000_0000;
array[451] <= 16'b0000_0000_0000_0000;
array[452] <= 16'b0000_0000_0000_0000;
array[453] <= 16'b0000_0000_0000_0000;
array[454] <= 16'b0000_0000_0000_0000;
array[455] <= 16'b0000_0000_0000_0000;
array[456] <= 16'b0000_0000_0000_0000;
array[457] <= 16'b0000_0000_0000_0000;
array[458] <= 16'b0000_0000_0000_0000;
array[459] <= 16'b0000_0000_0000_0000;
array[460] <= 16'b0000_0000_0000_0000;
array[461] <= 16'b0000_0000_0000_0000;
array[462] <= 16'b0000_0000_0000_0000;
array[463] <= 16'b0000_0000_0000_0000;
array[464] <= 16'b0000_0000_0000_0000;
array[465] <= 16'b0000_0000_0000_0000;
array[466] <= 16'b0000_0000_0000_0000;
array[467] <= 16'b0000_0000_0000_0000;
array[468] <= 16'b0000_0000_0000_0000;
array[469] <= 16'b0000_0000_0000_0000;
array[470] <= 16'b0000_0000_0000_0000;
array[471] <= 16'b0000_0000_0000_0000;
array[472] <= 16'b0000_0000_0000_0000;
array[473] <= 16'b0000_0000_0000_0000;
array[474] <= 16'b0000_0000_0000_0000;
array[475] <= 16'b0000_0000_0000_0000;
array[476] <= 16'b0000_0000_0000_0000;
array[477] <= 16'b0000_0000_0000_0000;
array[478] <= 16'b0000_0000_0000_0000;
array[479] <= 16'b0000_0000_0000_0000;
array[480] <= 16'b0000_0000_0000_0000;
array[481] <= 16'b0000_0000_0000_0000;
array[482] <= 16'b0000_0000_0000_0000;
array[483] <= 16'b0000_0000_0000_0000;
array[484] <= 16'b0000_0000_0000_0000;
array[485] <= 16'b0000_0000_0000_0000;
array[486] <= 16'b0000_0000_0000_0000;
array[487] <= 16'b0000_0000_0000_0000;
array[488] <= 16'b0000_0000_0000_0000;
array[489] <= 16'b0000_0000_0000_0000;
array[490] <= 16'b0000_0000_0000_0000;
array[491] <= 16'b0000_0000_0000_0000;
array[492] <= 16'b0000_0000_0000_0000;
array[493] <= 16'b0000_0000_0000_0000;
array[494] <= 16'b0000_0000_0000_0000;
array[495] <= 16'b0000_0000_0000_0000;
array[496] <= 16'b0000_0000_0000_0000;
array[497] <= 16'b0000_0000_0000_0000;
array[498] <= 16'b0000_0000_0000_0000;
array[499] <= 16'b0000_0000_0000_0000;
array[500] <= 16'b0000_0000_0000_0000;
array[501] <= 16'b0000_0000_0000_0000;
array[502] <= 16'b0000_0000_0000_0000;
array[503] <= 16'b0000_0000_0000_0000;
array[504] <= 16'b0000_0000_0000_0000;
array[505] <= 16'b0000_0000_0000_0000;
array[506] <= 16'b0000_0000_0000_0000;
array[507] <= 16'b0000_0000_0000_0000;
array[508] <= 16'b0000_0000_0000_0000;
array[509] <= 16'b0000_0000_0000_0000;
array[510] <= 16'b0000_0000_0000_0000;
array[511] <= 16'b0000_0000_0000_0000;
array[512] <= 16'b0000_0000_0000_0000;
array[513] <= 16'b0000_0000_0000_0000;
array[514] <= 16'b0000_0000_0000_0000;
array[515] <= 16'b0000_0000_0000_0000;
array[516] <= 16'b0000_0000_0000_0000;
array[517] <= 16'b0000_0000_0000_0000;
array[518] <= 16'b0000_0000_0000_0000;
array[519] <= 16'b0000_0000_0000_0000;
array[520] <= 16'b0000_0000_0000_0000;
array[521] <= 16'b0000_0000_0000_0000;
array[522] <= 16'b0000_0000_0000_0000;
array[523] <= 16'b0000_0000_0000_0000;
array[524] <= 16'b0000_0000_0000_0000;
array[525] <= 16'b0000_0000_0000_0000;
array[526] <= 16'b0000_0000_0000_0000;
array[527] <= 16'b0000_0000_0000_0000;
array[528] <= 16'b0000_0000_0000_0000;
array[529] <= 16'b0000_0000_0000_0000;
array[530] <= 16'b0000_0000_0000_0000;
array[531] <= 16'b0000_0000_0000_0000;
array[532] <= 16'b0000_0000_0000_0000;
array[533] <= 16'b0000_0000_0000_0000;
array[534] <= 16'b0000_0000_0000_0000;
array[535] <= 16'b0000_0000_0000_0000;
array[536] <= 16'b0000_0000_0000_0000;
array[537] <= 16'b0000_0000_0000_0000;
array[538] <= 16'b0000_0000_0000_0000;
array[539] <= 16'b0000_0000_0000_0000;
array[540] <= 16'b0000_0000_0000_0000;
array[541] <= 16'b0000_0000_0000_0000;
array[542] <= 16'b0000_0000_0000_0000;
array[543] <= 16'b0000_0000_0000_0000;
array[544] <= 16'b0000_0000_0000_0000;
array[545] <= 16'b0000_0000_0000_0000;
array[546] <= 16'b0000_0000_0000_0000;
array[547] <= 16'b0000_0000_0000_0000;
array[548] <= 16'b0000_0000_0000_0000;
array[549] <= 16'b0000_0000_0000_0000;
array[550] <= 16'b0000_0000_0000_0000;
array[551] <= 16'b0000_0000_0000_0000;
array[552] <= 16'b0000_0000_0000_0000;
array[553] <= 16'b0000_0000_0000_0000;
array[554] <= 16'b0000_0000_0000_0000;
array[555] <= 16'b0000_0000_0000_0000;
array[556] <= 16'b0000_0000_0000_0000;
array[557] <= 16'b0000_0000_0000_0000;
array[558] <= 16'b0000_0000_0000_0000;
array[559] <= 16'b0000_0000_0000_0000;
array[560] <= 16'b0000_0000_0000_0000;
array[561] <= 16'b0000_0000_0000_0000;
array[562] <= 16'b0000_0000_0000_0000;
array[563] <= 16'b0000_0000_0000_0000;
array[564] <= 16'b0000_0000_0000_0000;
array[565] <= 16'b0000_0000_0000_0000;
array[566] <= 16'b0000_0000_0000_0000;
array[567] <= 16'b0000_0000_0000_0000;
array[568] <= 16'b0000_0000_0000_0000;
array[569] <= 16'b0000_0000_0000_0000;
array[570] <= 16'b0000_0000_0000_0000;
array[571] <= 16'b0000_0000_0000_0000;
array[572] <= 16'b0000_0000_0000_0000;
array[573] <= 16'b0000_0000_0000_0000;
array[574] <= 16'b0000_0000_0000_0000;
array[575] <= 16'b0000_0000_0000_0000;
array[576] <= 16'b0000_0000_0000_0000;
array[577] <= 16'b0000_0000_0000_0000;
array[578] <= 16'b0000_0000_0000_0000;
array[579] <= 16'b0000_0000_0000_0000;
array[580] <= 16'b0000_0000_0000_0000;
array[581] <= 16'b0000_0000_0000_0000;
array[582] <= 16'b0000_0000_0000_0000;
array[583] <= 16'b0000_0000_0000_0000;
array[584] <= 16'b0000_0000_0000_0000;
array[585] <= 16'b0000_0000_0000_0000;
array[586] <= 16'b0000_0000_0000_0000;
array[587] <= 16'b0000_0000_0000_0000;
array[588] <= 16'b0000_0000_0000_0000;
array[589] <= 16'b0000_0000_0000_0000;
array[590] <= 16'b0000_0000_0000_0000;
array[591] <= 16'b0000_0000_0000_0000;
array[592] <= 16'b0000_0000_0000_0000;
array[593] <= 16'b0000_0000_0000_0000;
array[594] <= 16'b0000_0000_0000_0000;
array[595] <= 16'b0000_0000_0000_0000;
array[596] <= 16'b0000_0000_0000_0000;
array[597] <= 16'b0000_0000_0000_0000;
array[598] <= 16'b0000_0000_0000_0000;
array[599] <= 16'b0000_0000_0000_0000;
array[600] <= 16'b0000_0000_0000_0000;
array[601] <= 16'b0000_0000_0000_0000;
array[602] <= 16'b0000_0000_0000_0000;
array[603] <= 16'b0000_0000_0000_0000;
array[604] <= 16'b0000_0000_0000_0000;
array[605] <= 16'b0000_0000_0000_0000;
array[606] <= 16'b0000_0000_0000_0000;
array[607] <= 16'b0000_0000_0000_0000;
array[608] <= 16'b0000_0000_0000_0000;
array[609] <= 16'b0000_0000_0000_0000;
array[610] <= 16'b0000_0000_0000_0000;
array[611] <= 16'b0000_0000_0000_0000;
array[612] <= 16'b0000_0000_0000_0000;
array[613] <= 16'b0000_0000_0000_0000;
array[614] <= 16'b0000_0000_0000_0000;
array[615] <= 16'b0000_0000_0000_0000;
array[616] <= 16'b0000_0000_0000_0000;
array[617] <= 16'b0000_0000_0000_0000;
array[618] <= 16'b0000_0000_0000_0000;
array[619] <= 16'b0000_0000_0000_0000;
array[620] <= 16'b0000_0000_0000_0000;
array[621] <= 16'b0000_0000_0000_0000;
array[622] <= 16'b0000_0000_0000_0000;
array[623] <= 16'b0000_0000_0000_0000;
array[624] <= 16'b0000_0000_0000_0000;
array[625] <= 16'b0000_0000_0000_0000;
array[626] <= 16'b0000_0000_0000_0000;
array[627] <= 16'b0000_0000_0000_0000;
array[628] <= 16'b0000_0000_0000_0000;
array[629] <= 16'b0000_0000_0000_0000;
array[630] <= 16'b0000_0000_0000_0000;
array[631] <= 16'b0000_0000_0000_0000;
array[632] <= 16'b0000_0000_0000_0000;
array[633] <= 16'b0000_0000_0000_0000;
array[634] <= 16'b0000_0000_0000_0000;
array[635] <= 16'b0000_0000_0000_0000;
array[636] <= 16'b0000_0000_0000_0000;
array[637] <= 16'b0000_0000_0000_0000;
array[638] <= 16'b0000_0000_0000_0000;
array[639] <= 16'b0000_0000_0000_0000;
array[640] <= 16'b0000_0000_0000_0000;
array[641] <= 16'b0000_0000_0000_0000;
array[642] <= 16'b0000_0000_0000_0000;
array[643] <= 16'b0000_0000_0000_0000;
array[644] <= 16'b0000_0000_0000_0000;
array[645] <= 16'b0000_0000_0000_0000;
array[646] <= 16'b0000_0000_0000_0000;
array[647] <= 16'b0000_0000_0000_0000;
array[648] <= 16'b0000_0000_0000_0000;
array[649] <= 16'b0000_0000_0000_0000;
array[650] <= 16'b0000_0000_0000_0000;
array[651] <= 16'b0000_0000_0000_0000;
array[652] <= 16'b0000_0000_0000_0000;
array[653] <= 16'b0000_0000_0000_0000;
array[654] <= 16'b0000_0000_0000_0000;
array[655] <= 16'b0000_0000_0000_0000;
array[656] <= 16'b0000_0000_0000_0000;
array[657] <= 16'b0000_0000_0000_0000;
array[658] <= 16'b0000_0000_0000_0000;
array[659] <= 16'b0000_0000_0000_0000;
array[660] <= 16'b0000_0000_0000_0000;
array[661] <= 16'b0000_0000_0000_0000;
array[662] <= 16'b0000_0000_0000_0000;
array[663] <= 16'b0000_0000_0000_0000;
array[664] <= 16'b0000_0000_0000_0000;
array[665] <= 16'b0000_0000_0000_0000;
array[666] <= 16'b0000_0000_0000_0000;
array[667] <= 16'b0000_0000_0000_0000;
array[668] <= 16'b0000_0000_0000_0000;
array[669] <= 16'b0000_0000_0000_0000;
array[670] <= 16'b0000_0000_0000_0000;
array[671] <= 16'b0000_0000_0000_0000;
array[672] <= 16'b0000_0000_0000_0000;
array[673] <= 16'b0000_0000_0000_0000;
array[674] <= 16'b0000_0000_0000_0000;
array[675] <= 16'b0000_0000_0000_0000;
array[676] <= 16'b0000_0000_0000_0000;
array[677] <= 16'b0000_0000_0000_0000;
array[678] <= 16'b0000_0000_0000_0000;
array[679] <= 16'b0000_0000_0000_0000;
array[680] <= 16'b0000_0000_0000_0000;
array[681] <= 16'b0000_0000_0000_0000;
array[682] <= 16'b0000_0000_0000_0000;
array[683] <= 16'b0000_0000_0000_0000;
array[684] <= 16'b0000_0000_0000_0000;
array[685] <= 16'b0000_0000_0000_0000;
array[686] <= 16'b0000_0000_0000_0000;
array[687] <= 16'b0000_0000_0000_0000;
array[688] <= 16'b0000_0000_0000_0000;
array[689] <= 16'b0000_0000_0000_0000;
array[690] <= 16'b0000_0000_0000_0000;
array[691] <= 16'b0000_0000_0000_0000;
array[692] <= 16'b0000_0000_0000_0000;
array[693] <= 16'b0000_0000_0000_0000;
array[694] <= 16'b0000_0000_0000_0000;
array[695] <= 16'b0000_0000_0000_0000;
array[696] <= 16'b0000_0000_0000_0000;
array[697] <= 16'b0000_0000_0000_0000;
array[698] <= 16'b0000_0000_0000_0000;
array[699] <= 16'b0000_0000_0000_0000;
array[700] <= 16'b0000_0000_0000_0000;
array[701] <= 16'b0000_0000_0000_0000;
array[702] <= 16'b0000_0000_0000_0000;
array[703] <= 16'b0000_0000_0000_0000;
array[704] <= 16'b0000_0000_0000_0000;
array[705] <= 16'b0000_0000_0000_0000;
array[706] <= 16'b0000_0000_0000_0000;
array[707] <= 16'b0000_0000_0000_0000;
array[708] <= 16'b0000_0000_0000_0000;
array[709] <= 16'b0000_0000_0000_0000;
array[710] <= 16'b0000_0000_0000_0000;
array[711] <= 16'b0000_0000_0000_0000;
array[712] <= 16'b0000_0000_0000_0000;
array[713] <= 16'b0000_0000_0000_0000;
array[714] <= 16'b0000_0000_0000_0000;
array[715] <= 16'b0000_0000_0000_0000;
array[716] <= 16'b0000_0000_0000_0000;
array[717] <= 16'b0000_0000_0000_0000;
array[718] <= 16'b0000_0000_0000_0000;
array[719] <= 16'b0000_0000_0000_0000;
array[720] <= 16'b0000_0000_0000_0000;
array[721] <= 16'b0000_0000_0000_0000;
array[722] <= 16'b0000_0000_0000_0000;
array[723] <= 16'b0000_0000_0000_0000;
array[724] <= 16'b0000_0000_0000_0000;
array[725] <= 16'b0000_0000_0000_0000;
array[726] <= 16'b0000_0000_0000_0000;
array[727] <= 16'b0000_0000_0000_0000;
array[728] <= 16'b0000_0000_0000_0000;
array[729] <= 16'b0000_0000_0000_0000;
array[730] <= 16'b0000_0000_0000_0000;
array[731] <= 16'b0000_0000_0000_0000;
array[732] <= 16'b0000_0000_0000_0000;
array[733] <= 16'b0000_0000_0000_0000;
array[734] <= 16'b0000_0000_0000_0000;
array[735] <= 16'b0000_0000_0000_0000;
array[736] <= 16'b0000_0000_0000_0000;
array[737] <= 16'b0000_0000_0000_0000;
array[738] <= 16'b0000_0000_0000_0000;
array[739] <= 16'b0000_0000_0000_0000;
array[740] <= 16'b0000_0000_0000_0000;
array[741] <= 16'b0000_0000_0000_0000;
array[742] <= 16'b0000_0000_0000_0000;
array[743] <= 16'b0000_0000_0000_0000;
array[744] <= 16'b0000_0000_0000_0000;
array[745] <= 16'b0000_0000_0000_0000;
array[746] <= 16'b0000_0000_0000_0000;
array[747] <= 16'b0000_0000_0000_0000;
array[748] <= 16'b0000_0000_0000_0000;
array[749] <= 16'b0000_0000_0000_0000;
array[750] <= 16'b0000_0000_0000_0000;
array[751] <= 16'b0000_0000_0000_0000;
array[752] <= 16'b0000_0000_0000_0000;
array[753] <= 16'b0000_0000_0000_0000;
array[754] <= 16'b0000_0000_0000_0000;
array[755] <= 16'b0000_0000_0000_0000;
array[756] <= 16'b0000_0000_0000_0000;
array[757] <= 16'b0000_0000_0000_0000;
array[758] <= 16'b0000_0000_0000_0000;
array[759] <= 16'b0000_0000_0000_0000;
array[760] <= 16'b0000_0000_0000_0000;
array[761] <= 16'b0000_0000_0000_0000;
array[762] <= 16'b0000_0000_0000_0000;
array[763] <= 16'b0000_0000_0000_0000;
array[764] <= 16'b0000_0000_0000_0000;
array[765] <= 16'b0000_0000_0000_0000;
array[766] <= 16'b0000_0000_0000_0000;
array[767] <= 16'b0000_0000_0000_0000;
array[768] <= 16'b0000_0000_0000_0000;
array[769] <= 16'b0000_0000_0000_0000;
array[770] <= 16'b0000_0000_0000_0000;
array[771] <= 16'b0000_0000_0000_0000;
array[772] <= 16'b0000_0000_0000_0000;
array[773] <= 16'b0000_0000_0000_0000;
array[774] <= 16'b0000_0000_0000_0000;
array[775] <= 16'b0000_0000_0000_0000;
array[776] <= 16'b0000_0000_0000_0000;
array[777] <= 16'b0000_0000_0000_0000;
array[778] <= 16'b0000_0000_0000_0000;
array[779] <= 16'b0000_0000_0000_0000;
array[780] <= 16'b0000_0000_0000_0000;
array[781] <= 16'b0000_0000_0000_0000;
array[782] <= 16'b0000_0000_0000_0000;
array[783] <= 16'b0000_0000_0000_0000;
array[784] <= 16'b0000_0000_0000_0000;
array[785] <= 16'b0000_0000_0000_0000;
array[786] <= 16'b0000_0000_0000_0000;
array[787] <= 16'b0000_0000_0000_0000;
array[788] <= 16'b0000_0000_0000_0000;
array[789] <= 16'b0000_0000_0000_0000;
array[790] <= 16'b0000_0000_0000_0000;
array[791] <= 16'b0000_0000_0000_0000;
array[792] <= 16'b0000_0000_0000_0000;
array[793] <= 16'b0000_0000_0000_0000;
array[794] <= 16'b0000_0000_0000_0000;
array[795] <= 16'b0000_0000_0000_0000;
array[796] <= 16'b0000_0000_0000_0000;
array[797] <= 16'b0000_0000_0000_0000;
array[798] <= 16'b0000_0000_0000_0000;
array[799] <= 16'b0000_0000_0000_0000;
array[800] <= 16'b0000_0000_0000_0000;
array[801] <= 16'b0000_0000_0000_0000;
array[802] <= 16'b0000_0000_0000_0000;
array[803] <= 16'b0000_0000_0000_0000;
array[804] <= 16'b0000_0000_0000_0000;
array[805] <= 16'b0000_0000_0000_0000;
array[806] <= 16'b0000_0000_0000_0000;
array[807] <= 16'b0000_0000_0000_0000;
array[808] <= 16'b0000_0000_0000_0000;
array[809] <= 16'b0000_0000_0000_0000;
array[810] <= 16'b0000_0000_0000_0000;
array[811] <= 16'b0000_0000_0000_0000;
array[812] <= 16'b0000_0000_0000_0000;
array[813] <= 16'b0000_0000_0000_0000;
array[814] <= 16'b0000_0000_0000_0000;
array[815] <= 16'b0000_0000_0000_0000;
array[816] <= 16'b0000_0000_0000_0000;
array[817] <= 16'b0000_0000_0000_0000;
array[818] <= 16'b0000_0000_0000_0000;
array[819] <= 16'b0000_0000_0000_0000;
array[820] <= 16'b0000_0000_0000_0000;
array[821] <= 16'b0000_0000_0000_0000;
array[822] <= 16'b0000_0000_0000_0000;
array[823] <= 16'b0000_0000_0000_0000;
array[824] <= 16'b0000_0000_0000_0000;
array[825] <= 16'b0000_0000_0000_0000;
array[826] <= 16'b0000_0000_0000_0000;
array[827] <= 16'b0000_0000_0000_0000;
array[828] <= 16'b0000_0000_0000_0000;
array[829] <= 16'b0000_0000_0000_0000;
array[830] <= 16'b0000_0000_0000_0000;
array[831] <= 16'b0000_0000_0000_0000;
array[832] <= 16'b0000_0000_0000_0000;
array[833] <= 16'b0000_0000_0000_0000;
array[834] <= 16'b0000_0000_0000_0000;
array[835] <= 16'b0000_0000_0000_0000;
array[836] <= 16'b0000_0000_0000_0000;
array[837] <= 16'b0000_0000_0000_0000;
array[838] <= 16'b0000_0000_0000_0000;
array[839] <= 16'b0000_0000_0000_0000;
array[840] <= 16'b0000_0000_0000_0000;
array[841] <= 16'b0000_0000_0000_0000;
array[842] <= 16'b0000_0000_0000_0000;
array[843] <= 16'b0000_0000_0000_0000;
array[844] <= 16'b0000_0000_0000_0000;
array[845] <= 16'b0000_0000_0000_0000;
array[846] <= 16'b0000_0000_0000_0000;
array[847] <= 16'b0000_0000_0000_0000;
array[848] <= 16'b0000_0000_0000_0000;
array[849] <= 16'b0000_0000_0000_0000;
array[850] <= 16'b0000_0000_0000_0000;
array[851] <= 16'b0000_0000_0000_0000;
array[852] <= 16'b0000_0000_0000_0000;
array[853] <= 16'b0000_0000_0000_0000;
array[854] <= 16'b0000_0000_0000_0000;
array[855] <= 16'b0000_0000_0000_0000;
array[856] <= 16'b0000_0000_0000_0000;
array[857] <= 16'b0000_0000_0000_0000;
array[858] <= 16'b0000_0000_0000_0000;
array[859] <= 16'b0000_0000_0000_0000;
array[860] <= 16'b0000_0000_0000_0000;
array[861] <= 16'b0000_0000_0000_0000;
array[862] <= 16'b0000_0000_0000_0000;
array[863] <= 16'b0000_0000_0000_0000;
array[864] <= 16'b0000_0000_0000_0000;
array[865] <= 16'b0000_0000_0000_0000;
array[866] <= 16'b0000_0000_0000_0000;
array[867] <= 16'b0000_0000_0000_0000;
array[868] <= 16'b0000_0000_0000_0000;
array[869] <= 16'b0000_0000_0000_0000;
array[870] <= 16'b0000_0000_0000_0000;
array[871] <= 16'b0000_0000_0000_0000;
array[872] <= 16'b0000_0000_0000_0000;
array[873] <= 16'b0000_0000_0000_0000;
array[874] <= 16'b0000_0000_0000_0000;
array[875] <= 16'b0000_0000_0000_0000;
array[876] <= 16'b0000_0000_0000_0000;
array[877] <= 16'b0000_0000_0000_0000;
array[878] <= 16'b0000_0000_0000_0000;
array[879] <= 16'b0000_0000_0000_0000;
array[880] <= 16'b0000_0000_0000_0000;
array[881] <= 16'b0000_0000_0000_0000;
array[882] <= 16'b0000_0000_0000_0000;
array[883] <= 16'b0000_0000_0000_0000;
array[884] <= 16'b0000_0000_0000_0000;
array[885] <= 16'b0000_0000_0000_0000;
array[886] <= 16'b0000_0000_0000_0000;
array[887] <= 16'b0000_0000_0000_0000;
array[888] <= 16'b0000_0000_0000_0000;
array[889] <= 16'b0000_0000_0000_0000;
array[890] <= 16'b0000_0000_0000_0000;
array[891] <= 16'b0000_0000_0000_0000;
array[892] <= 16'b0000_0000_0000_0000;
array[893] <= 16'b0000_0000_0000_0000;
array[894] <= 16'b0000_0000_0000_0000;
array[895] <= 16'b0000_0000_0000_0000;
array[896] <= 16'b0000_0000_0000_0000;
array[897] <= 16'b0000_0000_0000_0000;
array[898] <= 16'b0000_0000_0000_0000;
array[899] <= 16'b0000_0000_0000_0000;
array[900] <= 16'b0000_0000_0000_0000;
array[901] <= 16'b0000_0000_0000_0000;
array[902] <= 16'b0000_0000_0000_0000;
array[903] <= 16'b0000_0000_0000_0000;
array[904] <= 16'b0000_0000_0000_0000;
array[905] <= 16'b0000_0000_0000_0000;
array[906] <= 16'b0000_0000_0000_0000;
array[907] <= 16'b0000_0000_0000_0000;
array[908] <= 16'b0000_0000_0000_0000;
array[909] <= 16'b0000_0000_0000_0000;
array[910] <= 16'b0000_0000_0000_0000;
array[911] <= 16'b0000_0000_0000_0000;
array[912] <= 16'b0000_0000_0000_0000;
array[913] <= 16'b0000_0000_0000_0000;
array[914] <= 16'b0000_0000_0000_0000;
array[915] <= 16'b0000_0000_0000_0000;
array[916] <= 16'b0000_0000_0000_0000;
array[917] <= 16'b0000_0000_0000_0000;
array[918] <= 16'b0000_0000_0000_0000;
array[919] <= 16'b0000_0000_0000_0000;
array[920] <= 16'b0000_0000_0000_0000;
array[921] <= 16'b0000_0000_0000_0000;
array[922] <= 16'b0000_0000_0000_0000;
array[923] <= 16'b0000_0000_0000_0000;
array[924] <= 16'b0000_0000_0000_0000;
array[925] <= 16'b0000_0000_0000_0000;
array[926] <= 16'b0000_0000_0000_0000;
array[927] <= 16'b0000_0000_0000_0000;
array[928] <= 16'b0000_0000_0000_0000;
array[929] <= 16'b0000_0000_0000_0000;
array[930] <= 16'b0000_0000_0000_0000;
array[931] <= 16'b0000_0000_0000_0000;
array[932] <= 16'b0000_0000_0000_0000;
array[933] <= 16'b0000_0000_0000_0000;
array[934] <= 16'b0000_0000_0000_0000;
array[935] <= 16'b0000_0000_0000_0000;
array[936] <= 16'b0000_0000_0000_0000;
array[937] <= 16'b0000_0000_0000_0000;
array[938] <= 16'b0000_0000_0000_0000;
array[939] <= 16'b0000_0000_0000_0000;
array[940] <= 16'b0000_0000_0000_0000;
array[941] <= 16'b0000_0000_0000_0000;
array[942] <= 16'b0000_0000_0000_0000;
array[943] <= 16'b0000_0000_0000_0000;
array[944] <= 16'b0000_0000_0000_0000;
array[945] <= 16'b0000_0000_0000_0000;
array[946] <= 16'b0000_0000_0000_0000;
array[947] <= 16'b0000_0000_0000_0000;
array[948] <= 16'b0000_0000_0000_0000;
array[949] <= 16'b0000_0000_0000_0000;
array[950] <= 16'b0000_0000_0000_0000;
array[951] <= 16'b0000_0000_0000_0000;
array[952] <= 16'b0000_0000_0000_0000;
array[953] <= 16'b0000_0000_0000_0000;
array[954] <= 16'b0000_0000_0000_0000;
array[955] <= 16'b0000_0000_0000_0000;
array[956] <= 16'b0000_0000_0000_0000;
array[957] <= 16'b0000_0000_0000_0000;
array[958] <= 16'b0000_0000_0000_0000;
array[959] <= 16'b0000_0000_0000_0000;
array[960] <= 16'b0000_0000_0000_0000;
array[961] <= 16'b0000_0000_0000_0000;
array[962] <= 16'b0000_0000_0000_0000;
array[963] <= 16'b0000_0000_0000_0000;
array[964] <= 16'b0000_0000_0000_0000;
array[965] <= 16'b0000_0000_0000_0000;
array[966] <= 16'b0000_0000_0000_0000;
array[967] <= 16'b0000_0000_0000_0000;
array[968] <= 16'b0000_0000_0000_0000;
array[969] <= 16'b0000_0000_0000_0000;
array[970] <= 16'b0000_0000_0000_0000;
array[971] <= 16'b0000_0000_0000_0000;
array[972] <= 16'b0000_0000_0000_0000;
array[973] <= 16'b0000_0000_0000_0000;
array[974] <= 16'b0000_0000_0000_0000;
array[975] <= 16'b0000_0000_0000_0000;
array[976] <= 16'b0000_0000_0000_0000;
array[977] <= 16'b0000_0000_0000_0000;
array[978] <= 16'b0000_0000_0000_0000;
array[979] <= 16'b0000_0000_0000_0000;
array[980] <= 16'b0000_0000_0000_0000;
array[981] <= 16'b0000_0000_0000_0000;
array[982] <= 16'b0000_0000_0000_0000;
array[983] <= 16'b0000_0000_0000_0000;
array[984] <= 16'b0000_0000_0000_0000;
array[985] <= 16'b0000_0000_0000_0000;
array[986] <= 16'b0000_0000_0000_0000;
array[987] <= 16'b0000_0000_0000_0000;
array[988] <= 16'b0000_0000_0000_0000;
array[989] <= 16'b0000_0000_0000_0000;
array[990] <= 16'b0000_0000_0000_0000;
array[991] <= 16'b0000_0000_0000_0000;
array[992] <= 16'b0000_0000_0000_0000;
array[993] <= 16'b0000_0000_0000_0000;
array[994] <= 16'b0000_0000_0000_0000;
array[995] <= 16'b0000_0000_0000_0000;
array[996] <= 16'b0000_0000_0000_0000;
array[997] <= 16'b0000_0000_0000_0000;
array[998] <= 16'b0000_0000_0000_0000;
array[999] <= 16'b0000_0000_0000_0000;
array[1000] <= 16'b0000_0000_0000_0000;
array[1001] <= 16'b0000_0000_0000_0000;
array[1002] <= 16'b0000_0000_0000_0000;
array[1003] <= 16'b0000_0000_0000_0000;
array[1004] <= 16'b0000_0000_0000_0000;
array[1005] <= 16'b0000_0000_0000_0000;
array[1006] <= 16'b0000_0000_0000_0000;
array[1007] <= 16'b0000_0000_0000_0000;
array[1008] <= 16'b0000_0000_0000_0000;
array[1009] <= 16'b0000_0000_0000_0000;
array[1010] <= 16'b0000_0000_0000_0000;
array[1011] <= 16'b0000_0000_0000_0000;
array[1012] <= 16'b0000_0000_0000_0000;
array[1013] <= 16'b0000_0000_0000_0000;
array[1014] <= 16'b0000_0000_0000_0000;
array[1015] <= 16'b0000_0000_0000_0000;
array[1016] <= 16'b0000_0000_0000_0000;
array[1017] <= 16'b0000_0000_0000_0000;
array[1018] <= 16'b0000_0000_0000_0000;
array[1019] <= 16'b0000_0000_0000_0000;
array[1020] <= 16'b0000_0000_0000_0000;
array[1021] <= 16'b0000_0000_0000_0000;
array[1022] <= 16'b0000_0000_0000_0000;
array[1023] <= 16'b0000_0000_0000_0000;
array[1024] <= 16'b0000_0000_0000_0000;
array[1025] <= 16'b0000_0000_0000_0000;
array[1026] <= 16'b0000_0000_0000_0000;
array[1027] <= 16'b0000_0000_0000_0000;
array[1028] <= 16'b0000_0000_0000_0000;
array[1029] <= 16'b0000_0000_0000_0000;
array[1030] <= 16'b0000_0000_0000_0000;
array[1031] <= 16'b0000_0000_0000_0000;
array[1032] <= 16'b0000_0000_0000_0000;
array[1033] <= 16'b0000_0000_0000_0000;
array[1034] <= 16'b0000_0000_0000_0000;
array[1035] <= 16'b0000_0000_0000_0000;
array[1036] <= 16'b0000_0000_0000_0000;
array[1037] <= 16'b0000_0000_0000_0000;
array[1038] <= 16'b0000_0000_0000_0000;
array[1039] <= 16'b0000_0000_0000_0000;
array[1040] <= 16'b0000_0000_0000_0000;
array[1041] <= 16'b0000_0000_0000_0000;
array[1042] <= 16'b0000_0000_0000_0000;
array[1043] <= 16'b0000_0000_0000_0000;
array[1044] <= 16'b0000_0000_0000_0000;
array[1045] <= 16'b0000_0000_0000_0000;
array[1046] <= 16'b0000_0000_0000_0000;
array[1047] <= 16'b0000_0000_0000_0000;
array[1048] <= 16'b0000_0000_0000_0000;
array[1049] <= 16'b0000_0000_0000_0000;
array[1050] <= 16'b0000_0000_0000_0000;
array[1051] <= 16'b0000_0000_0000_0000;
array[1052] <= 16'b0000_0000_0000_0000;
array[1053] <= 16'b0000_0000_0000_0000;
array[1054] <= 16'b0000_0000_0000_0000;
array[1055] <= 16'b0000_0000_0000_0000;
array[1056] <= 16'b0000_0000_0000_0000;
array[1057] <= 16'b0000_0000_0000_0000;
array[1058] <= 16'b0000_0000_0000_0000;
array[1059] <= 16'b0000_0000_0000_0000;
array[1060] <= 16'b0000_0000_0000_0000;
array[1061] <= 16'b0000_0000_0000_0000;
array[1062] <= 16'b0000_0000_0000_0000;
array[1063] <= 16'b0000_0000_0000_0000;
array[1064] <= 16'b0000_0000_0000_0000;
array[1065] <= 16'b0000_0000_0000_0000;
array[1066] <= 16'b0000_0000_0000_0000;
array[1067] <= 16'b0000_0000_0000_0000;
array[1068] <= 16'b0000_0000_0000_0000;
array[1069] <= 16'b0000_0000_0000_0000;
array[1070] <= 16'b0000_0000_0000_0000;
array[1071] <= 16'b0000_0000_0000_0000;
array[1072] <= 16'b0000_0000_0000_0000;
array[1073] <= 16'b0000_0000_0000_0000;
array[1074] <= 16'b0000_0000_0000_0000;
array[1075] <= 16'b0000_0000_0000_0000;
array[1076] <= 16'b0000_0000_0000_0000;
array[1077] <= 16'b0000_0000_0000_0000;
array[1078] <= 16'b0000_0000_0000_0000;
array[1079] <= 16'b0000_0000_0000_0000;
array[1080] <= 16'b0000_0000_0000_0000;
array[1081] <= 16'b0000_0000_0000_0000;
array[1082] <= 16'b0000_0000_0000_0000;
array[1083] <= 16'b0000_0000_0000_0000;
array[1084] <= 16'b0000_0000_0000_0000;
array[1085] <= 16'b0000_0000_0000_0000;
array[1086] <= 16'b0000_0000_0000_0000;
array[1087] <= 16'b0000_0000_0000_0000;
array[1088] <= 16'b0000_0000_0000_0000;
array[1089] <= 16'b0000_0000_0000_0000;
array[1090] <= 16'b0000_0000_0000_0000;
array[1091] <= 16'b0000_0000_0000_0000;
array[1092] <= 16'b0000_0000_0000_0000;
array[1093] <= 16'b0000_0000_0000_0000;
array[1094] <= 16'b0000_0000_0000_0000;
array[1095] <= 16'b0000_0000_0000_0000;
array[1096] <= 16'b0000_0000_0000_0000;
array[1097] <= 16'b0000_0000_0000_0000;
array[1098] <= 16'b0000_0000_0000_0000;
array[1099] <= 16'b0000_0000_0000_0000;
array[1100] <= 16'b0000_0000_0000_0000;
array[1101] <= 16'b0000_0000_0000_0000;
array[1102] <= 16'b0000_0000_0000_0000;
array[1103] <= 16'b0000_0000_0000_0000;
array[1104] <= 16'b0000_0000_0000_0000;
array[1105] <= 16'b0000_0000_0000_0000;
array[1106] <= 16'b0000_0000_0000_0000;
array[1107] <= 16'b0000_0000_0000_0000;
array[1108] <= 16'b0000_0000_0000_0000;
array[1109] <= 16'b0000_0000_0000_0000;
array[1110] <= 16'b0000_0000_0000_0000;
array[1111] <= 16'b0000_0000_0000_0000;
array[1112] <= 16'b0000_0000_0000_0000;
array[1113] <= 16'b0000_0000_0000_0000;
array[1114] <= 16'b0000_0000_0000_0000;
array[1115] <= 16'b0000_0000_0000_0000;
array[1116] <= 16'b0000_0000_0000_0000;
array[1117] <= 16'b0000_0000_0000_0000;
array[1118] <= 16'b0000_0000_0000_0000;
array[1119] <= 16'b0000_0000_0000_0000;
array[1120] <= 16'b0000_0000_0000_0000;
array[1121] <= 16'b0000_0000_0000_0000;
array[1122] <= 16'b0000_0000_0000_0000;
array[1123] <= 16'b0000_0000_0000_0000;
array[1124] <= 16'b0000_0000_0000_0000;
array[1125] <= 16'b0000_0000_0000_0000;
array[1126] <= 16'b0000_0000_0000_0000;
array[1127] <= 16'b0000_0000_0000_0000;
array[1128] <= 16'b0000_0000_0000_0000;
array[1129] <= 16'b0000_0000_0000_0000;
array[1130] <= 16'b0000_0000_0000_0000;
array[1131] <= 16'b0000_0000_0000_0000;
array[1132] <= 16'b0000_0000_0000_0000;
array[1133] <= 16'b0000_0000_0000_0000;
array[1134] <= 16'b0000_0000_0000_0000;
array[1135] <= 16'b0000_0000_0000_0000;
array[1136] <= 16'b0000_0000_0000_0000;
array[1137] <= 16'b0000_0000_0000_0000;
array[1138] <= 16'b0000_0000_0000_0000;
array[1139] <= 16'b0000_0000_0000_0000;
array[1140] <= 16'b0000_0000_0000_0000;
array[1141] <= 16'b0000_0000_0000_0000;
array[1142] <= 16'b0000_0000_0000_0000;
array[1143] <= 16'b0000_0000_0000_0000;
array[1144] <= 16'b0000_0000_0000_0000;
array[1145] <= 16'b0000_0000_0000_0000;
array[1146] <= 16'b0000_0000_0000_0000;
array[1147] <= 16'b0000_0000_0000_0000;
array[1148] <= 16'b0000_0000_0000_0000;
array[1149] <= 16'b0000_0000_0000_0000;
array[1150] <= 16'b0000_0000_0000_0000;
array[1151] <= 16'b0000_0000_0000_0000;
array[1152] <= 16'b0000_0000_0000_0000;
array[1153] <= 16'b0000_0000_0000_0000;
array[1154] <= 16'b0000_0000_0000_0000;
array[1155] <= 16'b0000_0000_0000_0000;
array[1156] <= 16'b0000_0000_0000_0000;
array[1157] <= 16'b0000_0000_0000_0000;
array[1158] <= 16'b0000_0000_0000_0000;
array[1159] <= 16'b0000_0000_0000_0000;
array[1160] <= 16'b0000_0000_0000_0000;
array[1161] <= 16'b0000_0000_0000_0000;
array[1162] <= 16'b0000_0000_0000_0000;
array[1163] <= 16'b0000_0000_0000_0000;
array[1164] <= 16'b0000_0000_0000_0000;
array[1165] <= 16'b0000_0000_0000_0000;
array[1166] <= 16'b0000_0000_0000_0000;
array[1167] <= 16'b0000_0000_0000_0000;
array[1168] <= 16'b0000_0000_0000_0000;
array[1169] <= 16'b0000_0000_0000_0000;
array[1170] <= 16'b0000_0000_0000_0000;
array[1171] <= 16'b0000_0000_0000_0000;
array[1172] <= 16'b0000_0000_0000_0000;
array[1173] <= 16'b0000_0000_0000_0000;
array[1174] <= 16'b0000_0000_0000_0000;
array[1175] <= 16'b0000_0000_0000_0000;
array[1176] <= 16'b0000_0000_0000_0000;
array[1177] <= 16'b0000_0000_0000_0000;
array[1178] <= 16'b0000_0000_0000_0000;
array[1179] <= 16'b0000_0000_0000_0000;
array[1180] <= 16'b0000_0000_0000_0000;
array[1181] <= 16'b0000_0000_0000_0000;
array[1182] <= 16'b0000_0000_0000_0000;
array[1183] <= 16'b0000_0000_0000_0000;
array[1184] <= 16'b0000_0000_0000_0000;
array[1185] <= 16'b0000_0000_0000_0000;
array[1186] <= 16'b0000_0000_0000_0000;
array[1187] <= 16'b0000_0000_0000_0000;
array[1188] <= 16'b0000_0000_0000_0000;
array[1189] <= 16'b0000_0000_0000_0000;
array[1190] <= 16'b0000_0000_0000_0000;
array[1191] <= 16'b0000_0000_0000_0000;
array[1192] <= 16'b0000_0000_0000_0000;
array[1193] <= 16'b0000_0000_0000_0000;
array[1194] <= 16'b0000_0000_0000_0000;
array[1195] <= 16'b0000_0000_0000_0000;
array[1196] <= 16'b0000_0000_0000_0000;
array[1197] <= 16'b0000_0000_0000_0000;
array[1198] <= 16'b0000_0000_0000_0000;
array[1199] <= 16'b0000_0000_0000_0000;
array[1200] <= 16'b0000_0000_0000_0000;
array[1201] <= 16'b0000_0000_0000_0000;
array[1202] <= 16'b0000_0000_0000_0000;
array[1203] <= 16'b0000_0000_0000_0000;
array[1204] <= 16'b0000_0000_0000_0000;
array[1205] <= 16'b0000_0000_0000_0000;
array[1206] <= 16'b0000_0000_0000_0000;
array[1207] <= 16'b0000_0000_0000_0000;
array[1208] <= 16'b0000_0000_0000_0000;
array[1209] <= 16'b0000_0000_0000_0000;
array[1210] <= 16'b0000_0000_0000_0000;
array[1211] <= 16'b0000_0000_0000_0000;
array[1212] <= 16'b0000_0000_0000_0000;
array[1213] <= 16'b0000_0000_0000_0000;
array[1214] <= 16'b0000_0000_0000_0000;
array[1215] <= 16'b0000_0000_0000_0000;
array[1216] <= 16'b0000_0000_0000_0000;
array[1217] <= 16'b0000_0000_0000_0000;
array[1218] <= 16'b0000_0000_0000_0000;
array[1219] <= 16'b0000_0000_0000_0000;
array[1220] <= 16'b0000_0000_0000_0000;
array[1221] <= 16'b0000_0000_0000_0000;
array[1222] <= 16'b0000_0000_0000_0000;
array[1223] <= 16'b0000_0000_0000_0000;
array[1224] <= 16'b0000_0000_0000_0000;
array[1225] <= 16'b0000_0000_0000_0000;
array[1226] <= 16'b0000_0000_0000_0000;
array[1227] <= 16'b0000_0000_0000_0000;
array[1228] <= 16'b0000_0000_0000_0000;
array[1229] <= 16'b0000_0000_0000_0000;
array[1230] <= 16'b0000_0000_0000_0000;
array[1231] <= 16'b0000_0000_0000_0000;
array[1232] <= 16'b0000_0000_0000_0000;
array[1233] <= 16'b0000_0000_0000_0000;
array[1234] <= 16'b0000_0000_0000_0000;
array[1235] <= 16'b0000_0000_0000_0000;
array[1236] <= 16'b0000_0000_0000_0000;
array[1237] <= 16'b0000_0000_0000_0000;
array[1238] <= 16'b0000_0000_0000_0000;
array[1239] <= 16'b0000_0000_0000_0000;
array[1240] <= 16'b0000_0000_0000_0000;
array[1241] <= 16'b0000_0000_0000_0000;
array[1242] <= 16'b0000_0000_0000_0000;
array[1243] <= 16'b0000_0000_0000_0000;
array[1244] <= 16'b0000_0000_0000_0000;
array[1245] <= 16'b0000_0000_0000_0000;
array[1246] <= 16'b0000_0000_0000_0000;
array[1247] <= 16'b0000_0000_0000_0000;
array[1248] <= 16'b0000_0000_0000_0000;
array[1249] <= 16'b0000_0000_0000_0000;
array[1250] <= 16'b0000_0000_0000_0000;
array[1251] <= 16'b0000_0000_0000_0000;
array[1252] <= 16'b0000_0000_0000_0000;
array[1253] <= 16'b0000_0000_0000_0000;
array[1254] <= 16'b0000_0000_0000_0000;
array[1255] <= 16'b0000_0000_0000_0000;
array[1256] <= 16'b0000_0000_0000_0000;
array[1257] <= 16'b0000_0000_0000_0000;
array[1258] <= 16'b0000_0000_0000_0000;
array[1259] <= 16'b0000_0000_0000_0000;
array[1260] <= 16'b0000_0000_0000_0000;
array[1261] <= 16'b0000_0000_0000_0000;
array[1262] <= 16'b0000_0000_0000_0000;
array[1263] <= 16'b0000_0000_0000_0000;
array[1264] <= 16'b0000_0000_0000_0000;
array[1265] <= 16'b0000_0000_0000_0000;
array[1266] <= 16'b0000_0000_0000_0000;
array[1267] <= 16'b0000_0000_0000_0000;
array[1268] <= 16'b0000_0000_0000_0000;
array[1269] <= 16'b0000_0000_0000_0000;
array[1270] <= 16'b0000_0000_0000_0000;
array[1271] <= 16'b0000_0000_0000_0000;
array[1272] <= 16'b0000_0000_0000_0000;
array[1273] <= 16'b0000_0000_0000_0000;
array[1274] <= 16'b0000_0000_0000_0000;
array[1275] <= 16'b0000_0000_0000_0000;
array[1276] <= 16'b0000_0000_0000_0000;
array[1277] <= 16'b0000_0000_0000_0000;
array[1278] <= 16'b0000_0000_0000_0000;
array[1279] <= 16'b0000_0000_0000_0000;
array[1280] <= 16'b0000_0000_0000_0000;
array[1281] <= 16'b0000_0000_0000_0000;
array[1282] <= 16'b0000_0000_0000_0000;
array[1283] <= 16'b0000_0000_0000_0000;
array[1284] <= 16'b0000_0000_0000_0000;
array[1285] <= 16'b0000_0000_0000_0000;
array[1286] <= 16'b0000_0000_0000_0000;
array[1287] <= 16'b0000_0000_0000_0000;
array[1288] <= 16'b0000_0000_0000_0000;
array[1289] <= 16'b0000_0000_0000_0000;
array[1290] <= 16'b0000_0000_0000_0000;
array[1291] <= 16'b0000_0000_0000_0000;
array[1292] <= 16'b0000_0000_0000_0000;
array[1293] <= 16'b0000_0000_0000_0000;
array[1294] <= 16'b0000_0000_0000_0000;
array[1295] <= 16'b0000_0000_0000_0000;
array[1296] <= 16'b0000_0000_0000_0000;
array[1297] <= 16'b0000_0000_0000_0000;
array[1298] <= 16'b0000_0000_0000_0000;
array[1299] <= 16'b0000_0000_0000_0000;
array[1300] <= 16'b0000_0000_0000_0000;
array[1301] <= 16'b0000_0000_0000_0000;
array[1302] <= 16'b0000_0000_0000_0000;
array[1303] <= 16'b0000_0000_0000_0000;
array[1304] <= 16'b0000_0000_0000_0000;
array[1305] <= 16'b0000_0000_0000_0000;
array[1306] <= 16'b0000_0000_0000_0000;
array[1307] <= 16'b0000_0000_0000_0000;
array[1308] <= 16'b0000_0000_0000_0000;
array[1309] <= 16'b0000_0000_0000_0000;
array[1310] <= 16'b0000_0000_0000_0000;
array[1311] <= 16'b0000_0000_0000_0000;
array[1312] <= 16'b0000_0000_0000_0000;
array[1313] <= 16'b0000_0000_0000_0000;
array[1314] <= 16'b0000_0000_0000_0000;
array[1315] <= 16'b0000_0000_0000_0000;
array[1316] <= 16'b0000_0000_0000_0000;
array[1317] <= 16'b0000_0000_0000_0000;
array[1318] <= 16'b0000_0000_0000_0000;
array[1319] <= 16'b0000_0000_0000_0000;
array[1320] <= 16'b0000_0000_0000_0000;
array[1321] <= 16'b0000_0000_0000_0000;
array[1322] <= 16'b0000_0000_0000_0000;
array[1323] <= 16'b0000_0000_0000_0000;
array[1324] <= 16'b0000_0000_0000_0000;
array[1325] <= 16'b0000_0000_0000_0000;
array[1326] <= 16'b0000_0000_0000_0000;
array[1327] <= 16'b0000_0000_0000_0000;
array[1328] <= 16'b0000_0000_0000_0000;
array[1329] <= 16'b0000_0000_0000_0000;
array[1330] <= 16'b0000_0000_0000_0000;
array[1331] <= 16'b0000_0000_0000_0000;
array[1332] <= 16'b0000_0000_0000_0000;
array[1333] <= 16'b0000_0000_0000_0000;
array[1334] <= 16'b0000_0000_0000_0000;
array[1335] <= 16'b0000_0000_0000_0000;
array[1336] <= 16'b0000_0000_0000_0000;
array[1337] <= 16'b0000_0000_0000_0000;
array[1338] <= 16'b0000_0000_0000_0000;
array[1339] <= 16'b0000_0000_0000_0000;
array[1340] <= 16'b0000_0000_0000_0000;
array[1341] <= 16'b0000_0000_0000_0000;
array[1342] <= 16'b0000_0000_0000_0000;
array[1343] <= 16'b0000_0000_0000_0000;
array[1344] <= 16'b0000_0000_0000_0000;
array[1345] <= 16'b0000_0000_0000_0000;
array[1346] <= 16'b0000_0000_0000_0000;
array[1347] <= 16'b0000_0000_0000_0000;
array[1348] <= 16'b0000_0000_0000_0000;
array[1349] <= 16'b0000_0000_0000_0000;
array[1350] <= 16'b0000_0000_0000_0000;
array[1351] <= 16'b0000_0000_0000_0000;
array[1352] <= 16'b0000_0000_0000_0000;
array[1353] <= 16'b0000_0000_0000_0000;
array[1354] <= 16'b0000_0000_0000_0000;
array[1355] <= 16'b0000_0000_0000_0000;
array[1356] <= 16'b0000_0000_0000_0000;
array[1357] <= 16'b0000_0000_0000_0000;
array[1358] <= 16'b0000_0000_0000_0000;
array[1359] <= 16'b0000_0000_0000_0000;
array[1360] <= 16'b0000_0000_0000_0000;
array[1361] <= 16'b0000_0000_0000_0000;
array[1362] <= 16'b0000_0000_0000_0000;
array[1363] <= 16'b0000_0000_0000_0000;
array[1364] <= 16'b0000_0000_0000_0000;
array[1365] <= 16'b0000_0000_0000_0000;
array[1366] <= 16'b0000_0000_0000_0000;
array[1367] <= 16'b0000_0000_0000_0000;
array[1368] <= 16'b0000_0000_0000_0000;
array[1369] <= 16'b0000_0000_0000_0000;
array[1370] <= 16'b0000_0000_0000_0000;
array[1371] <= 16'b0000_0000_0000_0000;
array[1372] <= 16'b0000_0000_0000_0000;
array[1373] <= 16'b0000_0000_0000_0000;
array[1374] <= 16'b0000_0000_0000_0000;
array[1375] <= 16'b0000_0000_0000_0000;
array[1376] <= 16'b0000_0000_0000_0000;
array[1377] <= 16'b0000_0000_0000_0000;
array[1378] <= 16'b0000_0000_0000_0000;
array[1379] <= 16'b0000_0000_0000_0000;
array[1380] <= 16'b0000_0000_0000_0000;
array[1381] <= 16'b0000_0000_0000_0000;
array[1382] <= 16'b0000_0000_0000_0000;
array[1383] <= 16'b0000_0000_0000_0000;
array[1384] <= 16'b0000_0000_0000_0000;
array[1385] <= 16'b0000_0000_0000_0000;
array[1386] <= 16'b0000_0000_0000_0000;
array[1387] <= 16'b0000_0000_0000_0000;
array[1388] <= 16'b0000_0000_0000_0000;
array[1389] <= 16'b0000_0000_0000_0000;
array[1390] <= 16'b0000_0000_0000_0000;
array[1391] <= 16'b0000_0000_0000_0000;
array[1392] <= 16'b0000_0000_0000_0000;
array[1393] <= 16'b0000_0000_0000_0000;
array[1394] <= 16'b0000_0000_0000_0000;
array[1395] <= 16'b0000_0000_0000_0000;
array[1396] <= 16'b0000_0000_0000_0000;
array[1397] <= 16'b0000_0000_0000_0000;
array[1398] <= 16'b0000_0000_0000_0000;
array[1399] <= 16'b0000_0000_0000_0000;
array[1400] <= 16'b0000_0000_0000_0000;
array[1401] <= 16'b0000_0000_0000_0000;
array[1402] <= 16'b0000_0000_0000_0000;
array[1403] <= 16'b0000_0000_0000_0000;
array[1404] <= 16'b0000_0000_0000_0000;
array[1405] <= 16'b0000_0000_0000_0000;
array[1406] <= 16'b0000_0000_0000_0000;
array[1407] <= 16'b0000_0000_0000_0000;
array[1408] <= 16'b0000_0000_0000_0000;
array[1409] <= 16'b0000_0000_0000_0000;
array[1410] <= 16'b0000_0000_0000_0000;
array[1411] <= 16'b0000_0000_0000_0000;
array[1412] <= 16'b0000_0000_0000_0000;
array[1413] <= 16'b0000_0000_0000_0000;
array[1414] <= 16'b0000_0000_0000_0000;
array[1415] <= 16'b0000_0000_0000_0000;
array[1416] <= 16'b0000_0000_0000_0000;
array[1417] <= 16'b0000_0000_0000_0000;
array[1418] <= 16'b0000_0000_0000_0000;
array[1419] <= 16'b0000_0000_0000_0000;
array[1420] <= 16'b0000_0000_0000_0000;
array[1421] <= 16'b0000_0000_0000_0000;
array[1422] <= 16'b0000_0000_0000_0000;
array[1423] <= 16'b0000_0000_0000_0000;
array[1424] <= 16'b0000_0000_0000_0000;
array[1425] <= 16'b0000_0000_0000_0000;
array[1426] <= 16'b0000_0000_0000_0000;
array[1427] <= 16'b0000_0000_0000_0000;
array[1428] <= 16'b0000_0000_0000_0000;
array[1429] <= 16'b0000_0000_0000_0000;
array[1430] <= 16'b0000_0000_0000_0000;
array[1431] <= 16'b0000_0000_0000_0000;
array[1432] <= 16'b0000_0000_0000_0000;
array[1433] <= 16'b0000_0000_0000_0000;
array[1434] <= 16'b0000_0000_0000_0000;
array[1435] <= 16'b0000_0000_0000_0000;
array[1436] <= 16'b0000_0000_0000_0000;
array[1437] <= 16'b0000_0000_0000_0000;
array[1438] <= 16'b0000_0000_0000_0000;
array[1439] <= 16'b0000_0000_0000_0000;
array[1440] <= 16'b0000_0000_0000_0000;
array[1441] <= 16'b0000_0000_0000_0000;
array[1442] <= 16'b0000_0000_0000_0000;
array[1443] <= 16'b0000_0000_0000_0000;
array[1444] <= 16'b0000_0000_0000_0000;
array[1445] <= 16'b0000_0000_0000_0000;
array[1446] <= 16'b0000_0000_0000_0000;
array[1447] <= 16'b0000_0000_0000_0000;
array[1448] <= 16'b0000_0000_0000_0000;
array[1449] <= 16'b0000_0000_0000_0000;
array[1450] <= 16'b0000_0000_0000_0000;
array[1451] <= 16'b0000_0000_0000_0000;
array[1452] <= 16'b0000_0000_0000_0000;
array[1453] <= 16'b0000_0000_0000_0000;
array[1454] <= 16'b0000_0000_0000_0000;
array[1455] <= 16'b0000_0000_0000_0000;
array[1456] <= 16'b0000_0000_0000_0000;
array[1457] <= 16'b0000_0000_0000_0000;
array[1458] <= 16'b0000_0000_0000_0000;
array[1459] <= 16'b0000_0000_0000_0000;
array[1460] <= 16'b0000_0000_0000_0000;
array[1461] <= 16'b0000_0000_0000_0000;
array[1462] <= 16'b0000_0000_0000_0000;
array[1463] <= 16'b0000_0000_0000_0000;
array[1464] <= 16'b0000_0000_0000_0000;
array[1465] <= 16'b0000_0000_0000_0000;
array[1466] <= 16'b0000_0000_0000_0000;
array[1467] <= 16'b0000_0000_0000_0000;
array[1468] <= 16'b0000_0000_0000_0000;
array[1469] <= 16'b0000_0000_0000_0000;
array[1470] <= 16'b0000_0000_0000_0000;
array[1471] <= 16'b0000_0000_0000_0000;
array[1472] <= 16'b0000_0000_0000_0000;
array[1473] <= 16'b0000_0000_0000_0000;
array[1474] <= 16'b0000_0000_0000_0000;
array[1475] <= 16'b0000_0000_0000_0000;
array[1476] <= 16'b0000_0000_0000_0000;
array[1477] <= 16'b0000_0000_0000_0000;
array[1478] <= 16'b0000_0000_0000_0000;
array[1479] <= 16'b0000_0000_0000_0000;
array[1480] <= 16'b0000_0000_0000_0000;
array[1481] <= 16'b0000_0000_0000_0000;
array[1482] <= 16'b0000_0000_0000_0000;
array[1483] <= 16'b0000_0000_0000_0000;
array[1484] <= 16'b0000_0000_0000_0000;
array[1485] <= 16'b0000_0000_0000_0000;
array[1486] <= 16'b0000_0000_0000_0000;
array[1487] <= 16'b0000_0000_0000_0000;
array[1488] <= 16'b0000_0000_0000_0000;
array[1489] <= 16'b0000_0000_0000_0000;
array[1490] <= 16'b0000_0000_0000_0000;
array[1491] <= 16'b0000_0000_0000_0000;
array[1492] <= 16'b0000_0000_0000_0000;
array[1493] <= 16'b0000_0000_0000_0000;
array[1494] <= 16'b0000_0000_0000_0000;
array[1495] <= 16'b0000_0000_0000_0000;
array[1496] <= 16'b0000_0000_0000_0000;
array[1497] <= 16'b0000_0000_0000_0000;
array[1498] <= 16'b0000_0000_0000_0000;
array[1499] <= 16'b0000_0000_0000_0000;
array[1500] <= 16'b0000_0000_0000_0000;
array[1501] <= 16'b0000_0000_0000_0000;
array[1502] <= 16'b0000_0000_0000_0000;
array[1503] <= 16'b0000_0000_0000_0000;
array[1504] <= 16'b0000_0000_0000_0000;
array[1505] <= 16'b0000_0000_0000_0000;
array[1506] <= 16'b0000_0000_0000_0000;
array[1507] <= 16'b0000_0000_0000_0000;
array[1508] <= 16'b0000_0000_0000_0000;
array[1509] <= 16'b0000_0000_0000_0000;
array[1510] <= 16'b0000_0000_0000_0000;
array[1511] <= 16'b0000_0000_0000_0000;
array[1512] <= 16'b0000_0000_0000_0000;
array[1513] <= 16'b0000_0000_0000_0000;
array[1514] <= 16'b0000_0000_0000_0000;
array[1515] <= 16'b0000_0000_0000_0000;
array[1516] <= 16'b0000_0000_0000_0000;
array[1517] <= 16'b0000_0000_0000_0000;
array[1518] <= 16'b0000_0000_0000_0000;
array[1519] <= 16'b0000_0000_0000_0000;
array[1520] <= 16'b0000_0000_0000_0000;
array[1521] <= 16'b0000_0000_0000_0000;
array[1522] <= 16'b0000_0000_0000_0000;
array[1523] <= 16'b0000_0000_0000_0000;
array[1524] <= 16'b0000_0000_0000_0000;
array[1525] <= 16'b0000_0000_0000_0000;
array[1526] <= 16'b0000_0000_0000_0000;
array[1527] <= 16'b0000_0000_0000_0000;
array[1528] <= 16'b0000_0000_0000_0000;
array[1529] <= 16'b0000_0000_0000_0000;
array[1530] <= 16'b0000_0000_0000_0000;
array[1531] <= 16'b0000_0000_0000_0000;
array[1532] <= 16'b0000_0000_0000_0000;
array[1533] <= 16'b0000_0000_0000_0000;
array[1534] <= 16'b0000_0000_0000_0000;
array[1535] <= 16'b0000_0000_0000_0000;
array[1536] <= 16'b0000_0000_0000_0000;
array[1537] <= 16'b0000_0000_0000_0000;
array[1538] <= 16'b0000_0000_0000_0000;
array[1539] <= 16'b0000_0000_0000_0000;
array[1540] <= 16'b0000_0000_0000_0000;
array[1541] <= 16'b0000_0000_0000_0000;
array[1542] <= 16'b0000_0000_0000_0000;
array[1543] <= 16'b0000_0000_0000_0000;
array[1544] <= 16'b0000_0000_0000_0000;
array[1545] <= 16'b0000_0000_0000_0000;
array[1546] <= 16'b0000_0000_0000_0000;
array[1547] <= 16'b0000_0000_0000_0000;
array[1548] <= 16'b0000_0000_0000_0000;
array[1549] <= 16'b0000_0000_0000_0000;
array[1550] <= 16'b0000_0000_0000_0000;
array[1551] <= 16'b0000_0000_0000_0000;
array[1552] <= 16'b0000_0000_0000_0000;
array[1553] <= 16'b0000_0000_0000_0000;
array[1554] <= 16'b0000_0000_0000_0000;
array[1555] <= 16'b0000_0000_0000_0000;
array[1556] <= 16'b0000_0000_0000_0000;
array[1557] <= 16'b0000_0000_0000_0000;
array[1558] <= 16'b0000_0000_0000_0000;
array[1559] <= 16'b0000_0000_0000_0000;
array[1560] <= 16'b0000_0000_0000_0000;
array[1561] <= 16'b0000_0000_0000_0000;
array[1562] <= 16'b0000_0000_0000_0000;
array[1563] <= 16'b0000_0000_0000_0000;
array[1564] <= 16'b0000_0000_0000_0000;
array[1565] <= 16'b0000_0000_0000_0000;
array[1566] <= 16'b0000_0000_0000_0000;
array[1567] <= 16'b0000_0000_0000_0000;
array[1568] <= 16'b0000_0000_0000_0000;
array[1569] <= 16'b0000_0000_0000_0000;
array[1570] <= 16'b0000_0000_0000_0000;
array[1571] <= 16'b0000_0000_0000_0000;
array[1572] <= 16'b0000_0000_0000_0000;
array[1573] <= 16'b0000_0000_0000_0000;
array[1574] <= 16'b0000_0000_0000_0000;
array[1575] <= 16'b0000_0000_0000_0000;
array[1576] <= 16'b0000_0000_0000_0000;
array[1577] <= 16'b0000_0000_0000_0000;
array[1578] <= 16'b0000_0000_0000_0000;
array[1579] <= 16'b0000_0000_0000_0000;
array[1580] <= 16'b0000_0000_0000_0000;
array[1581] <= 16'b0000_0000_0000_0000;
array[1582] <= 16'b0000_0000_0000_0000;
array[1583] <= 16'b0000_0000_0000_0000;
array[1584] <= 16'b0000_0000_0000_0000;
array[1585] <= 16'b0000_0000_0000_0000;
array[1586] <= 16'b0000_0000_0000_0000;
array[1587] <= 16'b0000_0000_0000_0000;
array[1588] <= 16'b0000_0000_0000_0000;
array[1589] <= 16'b0000_0000_0000_0000;
array[1590] <= 16'b0000_0000_0000_0000;
array[1591] <= 16'b0000_0000_0000_0000;
array[1592] <= 16'b0000_0000_0000_0000;
array[1593] <= 16'b0000_0000_0000_0000;
array[1594] <= 16'b0000_0000_0000_0000;
array[1595] <= 16'b0000_0000_0000_0000;
array[1596] <= 16'b0000_0000_0000_0000;
array[1597] <= 16'b0000_0000_0000_0000;
array[1598] <= 16'b0000_0000_0000_0000;
array[1599] <= 16'b0000_0000_0000_0000;
array[1600] <= 16'b0000_0000_0000_0000;
array[1601] <= 16'b0000_0000_0000_0000;
array[1602] <= 16'b0000_0000_0000_0000;
array[1603] <= 16'b0000_0000_0000_0000;
array[1604] <= 16'b0000_0000_0000_0000;
array[1605] <= 16'b0000_0000_0000_0000;
array[1606] <= 16'b0000_0000_0000_0000;
array[1607] <= 16'b0000_0000_0000_0000;
array[1608] <= 16'b0000_0000_0000_0000;
array[1609] <= 16'b0000_0000_0000_0000;
array[1610] <= 16'b0000_0000_0000_0000;
array[1611] <= 16'b0000_0000_0000_0000;
array[1612] <= 16'b0000_0000_0000_0000;
array[1613] <= 16'b0000_0000_0000_0000;
array[1614] <= 16'b0000_0000_0000_0000;
array[1615] <= 16'b0000_0000_0000_0000;
array[1616] <= 16'b0000_0000_0000_0000;
array[1617] <= 16'b0000_0000_0000_0000;
array[1618] <= 16'b0000_0000_0000_0000;
array[1619] <= 16'b0000_0000_0000_0000;
array[1620] <= 16'b0000_0000_0000_0000;
array[1621] <= 16'b0000_0000_0000_0000;
array[1622] <= 16'b0000_0000_0000_0000;
array[1623] <= 16'b0000_0000_0000_0000;
array[1624] <= 16'b0000_0000_0000_0000;
array[1625] <= 16'b0000_0000_0000_0000;
array[1626] <= 16'b0000_0000_0000_0000;
array[1627] <= 16'b0000_0000_0000_0000;
array[1628] <= 16'b0000_0000_0000_0000;
array[1629] <= 16'b0000_0000_0000_0000;
array[1630] <= 16'b0000_0000_0000_0000;
array[1631] <= 16'b0000_0000_0000_0000;
array[1632] <= 16'b0000_0000_0000_0000;
array[1633] <= 16'b0000_0000_0000_0000;
array[1634] <= 16'b0000_0000_0000_0000;
array[1635] <= 16'b0000_0000_0000_0000;
array[1636] <= 16'b0000_0000_0000_0000;
array[1637] <= 16'b0000_0000_0000_0000;
array[1638] <= 16'b0000_0000_0000_0000;
array[1639] <= 16'b0000_0000_0000_0000;
array[1640] <= 16'b0000_0000_0000_0000;
array[1641] <= 16'b0000_0000_0000_0000;
array[1642] <= 16'b0000_0000_0000_0000;
array[1643] <= 16'b0000_0000_0000_0000;
array[1644] <= 16'b0000_0000_0000_0000;
array[1645] <= 16'b0000_0000_0000_0000;
array[1646] <= 16'b0000_0000_0000_0000;
array[1647] <= 16'b0000_0000_0000_0000;
array[1648] <= 16'b0000_0000_0000_0000;
array[1649] <= 16'b0000_0000_0000_0000;
array[1650] <= 16'b0000_0000_0000_0000;
array[1651] <= 16'b0000_0000_0000_0000;
array[1652] <= 16'b0000_0000_0000_0000;
array[1653] <= 16'b0000_0000_0000_0000;
array[1654] <= 16'b0000_0000_0000_0000;
array[1655] <= 16'b0000_0000_0000_0000;
array[1656] <= 16'b0000_0000_0000_0000;
array[1657] <= 16'b0000_0000_0000_0000;
array[1658] <= 16'b0000_0000_0000_0000;
array[1659] <= 16'b0000_0000_0000_0000;
array[1660] <= 16'b0000_0000_0000_0000;
array[1661] <= 16'b0000_0000_0000_0000;
array[1662] <= 16'b0000_0000_0000_0000;
array[1663] <= 16'b0000_0000_0000_0000;
array[1664] <= 16'b0000_0000_0000_0000;
array[1665] <= 16'b0000_0000_0000_0000;
array[1666] <= 16'b0000_0000_0000_0000;
array[1667] <= 16'b0000_0000_0000_0000;
array[1668] <= 16'b0000_0000_0000_0000;
array[1669] <= 16'b0000_0000_0000_0000;
array[1670] <= 16'b0000_0000_0000_0000;
array[1671] <= 16'b0000_0000_0000_0000;
array[1672] <= 16'b0000_0000_0000_0000;
array[1673] <= 16'b0000_0000_0000_0000;
array[1674] <= 16'b0000_0000_0000_0000;
array[1675] <= 16'b0000_0000_0000_0000;
array[1676] <= 16'b0000_0000_0000_0000;
array[1677] <= 16'b0000_0000_0000_0000;
array[1678] <= 16'b0000_0000_0000_0000;
array[1679] <= 16'b0000_0000_0000_0000;
array[1680] <= 16'b0000_0000_0000_0000;
array[1681] <= 16'b0000_0000_0000_0000;
array[1682] <= 16'b0000_0000_0000_0000;
array[1683] <= 16'b0000_0000_0000_0000;
array[1684] <= 16'b0000_0000_0000_0000;
array[1685] <= 16'b0000_0000_0000_0000;
array[1686] <= 16'b0000_0000_0000_0000;
array[1687] <= 16'b0000_0000_0000_0000;
array[1688] <= 16'b0000_0000_0000_0000;
array[1689] <= 16'b0000_0000_0000_0000;
array[1690] <= 16'b0000_0000_0000_0000;
array[1691] <= 16'b0000_0000_0000_0000;
array[1692] <= 16'b0000_0000_0000_0000;
array[1693] <= 16'b0000_0000_0000_0000;
array[1694] <= 16'b0000_0000_0000_0000;
array[1695] <= 16'b0000_0000_0000_0000;
array[1696] <= 16'b0000_0000_0000_0000;
array[1697] <= 16'b0000_0000_0000_0000;
array[1698] <= 16'b0000_0000_0000_0000;
array[1699] <= 16'b0000_0000_0000_0000;
array[1700] <= 16'b0000_0000_0000_0000;
array[1701] <= 16'b0000_0000_0000_0000;
array[1702] <= 16'b0000_0000_0000_0000;
array[1703] <= 16'b0000_0000_0000_0000;
array[1704] <= 16'b0000_0000_0000_0000;
array[1705] <= 16'b0000_0000_0000_0000;
array[1706] <= 16'b0000_0000_0000_0000;
array[1707] <= 16'b0000_0000_0000_0000;
array[1708] <= 16'b0000_0000_0000_0000;
array[1709] <= 16'b0000_0000_0000_0000;
array[1710] <= 16'b0000_0000_0000_0000;
array[1711] <= 16'b0000_0000_0000_0000;
array[1712] <= 16'b0000_0000_0000_0000;
array[1713] <= 16'b0000_0000_0000_0000;
array[1714] <= 16'b0000_0000_0000_0000;
array[1715] <= 16'b0000_0000_0000_0000;
array[1716] <= 16'b0000_0000_0000_0000;
array[1717] <= 16'b0000_0000_0000_0000;
array[1718] <= 16'b0000_0000_0000_0000;
array[1719] <= 16'b0000_0000_0000_0000;
array[1720] <= 16'b0000_0000_0000_0000;
array[1721] <= 16'b0000_0000_0000_0000;
array[1722] <= 16'b0000_0000_0000_0000;
array[1723] <= 16'b0000_0000_0000_0000;
array[1724] <= 16'b0000_0000_0000_0000;
array[1725] <= 16'b0000_0000_0000_0000;
array[1726] <= 16'b0000_0000_0000_0000;
array[1727] <= 16'b0000_0000_0000_0000;
array[1728] <= 16'b0000_0000_0000_0000;
array[1729] <= 16'b0000_0000_0000_0000;
array[1730] <= 16'b0000_0000_0000_0000;
array[1731] <= 16'b0000_0000_0000_0000;
array[1732] <= 16'b0000_0000_0000_0000;
array[1733] <= 16'b0000_0000_0000_0000;
array[1734] <= 16'b0000_0000_0000_0000;
array[1735] <= 16'b0000_0000_0000_0000;
array[1736] <= 16'b0000_0000_0000_0000;
array[1737] <= 16'b0000_0000_0000_0000;
array[1738] <= 16'b0000_0000_0000_0000;
array[1739] <= 16'b0000_0000_0000_0000;
array[1740] <= 16'b0000_0000_0000_0000;
array[1741] <= 16'b0000_0000_0000_0000;
array[1742] <= 16'b0000_0000_0000_0000;
array[1743] <= 16'b0000_0000_0000_0000;
array[1744] <= 16'b0000_0000_0000_0000;
array[1745] <= 16'b0000_0000_0000_0000;
array[1746] <= 16'b0000_0000_0000_0000;
array[1747] <= 16'b0000_0000_0000_0000;
array[1748] <= 16'b0000_0000_0000_0000;
array[1749] <= 16'b0000_0000_0000_0000;
array[1750] <= 16'b0000_0000_0000_0000;
array[1751] <= 16'b0000_0000_0000_0000;
array[1752] <= 16'b0000_0000_0000_0000;
array[1753] <= 16'b0000_0000_0000_0000;
array[1754] <= 16'b0000_0000_0000_0000;
array[1755] <= 16'b0000_0000_0000_0000;
array[1756] <= 16'b0000_0000_0000_0000;
array[1757] <= 16'b0000_0000_0000_0000;
array[1758] <= 16'b0000_0000_0000_0000;
array[1759] <= 16'b0000_0000_0000_0000;
array[1760] <= 16'b0000_0000_0000_0000;
array[1761] <= 16'b0000_0000_0000_0000;
array[1762] <= 16'b0000_0000_0000_0000;
array[1763] <= 16'b0000_0000_0000_0000;
array[1764] <= 16'b0000_0000_0000_0000;
array[1765] <= 16'b0000_0000_0000_0000;
array[1766] <= 16'b0000_0000_0000_0000;
array[1767] <= 16'b0000_0000_0000_0000;
array[1768] <= 16'b0000_0000_0000_0000;
array[1769] <= 16'b0000_0000_0000_0000;
array[1770] <= 16'b0000_0000_0000_0000;
array[1771] <= 16'b0000_0000_0000_0000;
array[1772] <= 16'b0000_0000_0000_0000;
array[1773] <= 16'b0000_0000_0000_0000;
array[1774] <= 16'b0000_0000_0000_0000;
array[1775] <= 16'b0000_0000_0000_0000;
array[1776] <= 16'b0000_0000_0000_0000;
array[1777] <= 16'b0000_0000_0000_0000;
array[1778] <= 16'b0000_0000_0000_0000;
array[1779] <= 16'b0000_0000_0000_0000;
array[1780] <= 16'b0000_0000_0000_0000;
array[1781] <= 16'b0000_0000_0000_0000;
array[1782] <= 16'b0000_0000_0000_0000;
array[1783] <= 16'b0000_0000_0000_0000;
array[1784] <= 16'b0000_0000_0000_0000;
array[1785] <= 16'b0000_0000_0000_0000;
array[1786] <= 16'b0000_0000_0000_0000;
array[1787] <= 16'b0000_0000_0000_0000;
array[1788] <= 16'b0000_0000_0000_0000;
array[1789] <= 16'b0000_0000_0000_0000;
array[1790] <= 16'b0000_0000_0000_0000;
array[1791] <= 16'b0000_0000_0000_0000;
array[1792] <= 16'b0000_0000_0000_0000;
array[1793] <= 16'b0000_0000_0000_0000;
array[1794] <= 16'b0000_0000_0000_0000;
array[1795] <= 16'b0000_0000_0000_0000;
array[1796] <= 16'b0000_0000_0000_0000;
array[1797] <= 16'b0000_0000_0000_0000;
array[1798] <= 16'b0000_0000_0000_0000;
array[1799] <= 16'b0000_0000_0000_0000;
array[1800] <= 16'b0000_0000_0000_0000;
array[1801] <= 16'b0000_0000_0000_0000;
array[1802] <= 16'b0000_0000_0000_0000;
array[1803] <= 16'b0000_0000_0000_0000;
array[1804] <= 16'b0000_0000_0000_0000;
array[1805] <= 16'b0000_0000_0000_0000;
array[1806] <= 16'b0000_0000_0000_0000;
array[1807] <= 16'b0000_0000_0000_0000;
array[1808] <= 16'b0000_0000_0000_0000;
array[1809] <= 16'b0000_0000_0000_0000;
array[1810] <= 16'b0000_0000_0000_0000;
array[1811] <= 16'b0000_0000_0000_0000;
array[1812] <= 16'b0000_0000_0000_0000;
array[1813] <= 16'b0000_0000_0000_0000;
array[1814] <= 16'b0000_0000_0000_0000;
array[1815] <= 16'b0000_0000_0000_0000;
array[1816] <= 16'b0000_0000_0000_0000;
array[1817] <= 16'b0000_0000_0000_0000;
array[1818] <= 16'b0000_0000_0000_0000;
array[1819] <= 16'b0000_0000_0000_0000;
array[1820] <= 16'b0000_0000_0000_0000;
array[1821] <= 16'b0000_0000_0000_0000;
array[1822] <= 16'b0000_0000_0000_0000;
array[1823] <= 16'b0000_0000_0000_0000;
array[1824] <= 16'b0000_0000_0000_0000;
array[1825] <= 16'b0000_0000_0000_0000;
array[1826] <= 16'b0000_0000_0000_0000;
array[1827] <= 16'b0000_0000_0000_0000;
array[1828] <= 16'b0000_0000_0000_0000;
array[1829] <= 16'b0000_0000_0000_0000;
array[1830] <= 16'b0000_0000_0000_0000;
array[1831] <= 16'b0000_0000_0000_0000;
array[1832] <= 16'b0000_0000_0000_0000;
array[1833] <= 16'b0000_0000_0000_0000;
array[1834] <= 16'b0000_0000_0000_0000;
array[1835] <= 16'b0000_0000_0000_0000;
array[1836] <= 16'b0000_0000_0000_0000;
array[1837] <= 16'b0000_0000_0000_0000;
array[1838] <= 16'b0000_0000_0000_0000;
array[1839] <= 16'b0000_0000_0000_0000;
array[1840] <= 16'b0000_0000_0000_0000;
array[1841] <= 16'b0000_0000_0000_0000;
array[1842] <= 16'b0000_0000_0000_0000;
array[1843] <= 16'b0000_0000_0000_0000;
array[1844] <= 16'b0000_0000_0000_0000;
array[1845] <= 16'b0000_0000_0000_0000;
array[1846] <= 16'b0000_0000_0000_0000;
array[1847] <= 16'b0000_0000_0000_0000;
array[1848] <= 16'b0000_0000_0000_0000;
array[1849] <= 16'b0000_0000_0000_0000;
array[1850] <= 16'b0000_0000_0000_0000;
array[1851] <= 16'b0000_0000_0000_0000;
array[1852] <= 16'b0000_0000_0000_0000;
array[1853] <= 16'b0000_0000_0000_0000;
array[1854] <= 16'b0000_0000_0000_0000;
array[1855] <= 16'b0000_0000_0000_0000;
array[1856] <= 16'b0000_0000_0000_0000;
array[1857] <= 16'b0000_0000_0000_0000;
array[1858] <= 16'b0000_0000_0000_0000;
array[1859] <= 16'b0000_0000_0000_0000;
array[1860] <= 16'b0000_0000_0000_0000;
array[1861] <= 16'b0000_0000_0000_0000;
array[1862] <= 16'b0000_0000_0000_0000;
array[1863] <= 16'b0000_0000_0000_0000;
array[1864] <= 16'b0000_0000_0000_0000;
array[1865] <= 16'b0000_0000_0000_0000;
array[1866] <= 16'b0000_0000_0000_0000;
array[1867] <= 16'b0000_0000_0000_0000;
array[1868] <= 16'b0000_0000_0000_0000;
array[1869] <= 16'b0000_0000_0000_0000;
array[1870] <= 16'b0000_0000_0000_0000;
array[1871] <= 16'b0000_0000_0000_0000;
array[1872] <= 16'b0000_0000_0000_0000;
array[1873] <= 16'b0000_0000_0000_0000;
array[1874] <= 16'b0000_0000_0000_0000;
array[1875] <= 16'b0000_0000_0000_0000;
array[1876] <= 16'b0000_0000_0000_0000;
array[1877] <= 16'b0000_0000_0000_0000;
array[1878] <= 16'b0000_0000_0000_0000;
array[1879] <= 16'b0000_0000_0000_0000;
array[1880] <= 16'b0000_0000_0000_0000;
array[1881] <= 16'b0000_0000_0000_0000;
array[1882] <= 16'b0000_0000_0000_0000;
array[1883] <= 16'b0000_0000_0000_0000;
array[1884] <= 16'b0000_0000_0000_0000;
array[1885] <= 16'b0000_0000_0000_0000;
array[1886] <= 16'b0000_0000_0000_0000;
array[1887] <= 16'b0000_0000_0000_0000;
array[1888] <= 16'b0000_0000_0000_0000;
array[1889] <= 16'b0000_0000_0000_0000;
array[1890] <= 16'b0000_0000_0000_0000;
array[1891] <= 16'b0000_0000_0000_0000;
array[1892] <= 16'b0000_0000_0000_0000;
array[1893] <= 16'b0000_0000_0000_0000;
array[1894] <= 16'b0000_0000_0000_0000;
array[1895] <= 16'b0000_0000_0000_0000;
array[1896] <= 16'b0000_0000_0000_0000;
array[1897] <= 16'b0000_0000_0000_0000;
array[1898] <= 16'b0000_0000_0000_0000;
array[1899] <= 16'b0000_0000_0000_0000;
array[1900] <= 16'b0000_0000_0000_0000;
array[1901] <= 16'b0000_0000_0000_0000;
array[1902] <= 16'b0000_0000_0000_0000;
array[1903] <= 16'b0000_0000_0000_0000;
array[1904] <= 16'b0000_0000_0000_0000;
array[1905] <= 16'b0000_0000_0000_0000;
array[1906] <= 16'b0000_0000_0000_0000;
array[1907] <= 16'b0000_0000_0000_0000;
array[1908] <= 16'b0000_0000_0000_0000;
array[1909] <= 16'b0000_0000_0000_0000;
array[1910] <= 16'b0000_0000_0000_0000;
array[1911] <= 16'b0000_0000_0000_0000;
array[1912] <= 16'b0000_0000_0000_0000;
array[1913] <= 16'b0000_0000_0000_0000;
array[1914] <= 16'b0000_0000_0000_0000;
array[1915] <= 16'b0000_0000_0000_0000;
array[1916] <= 16'b0000_0000_0000_0000;
array[1917] <= 16'b0000_0000_0000_0000;
array[1918] <= 16'b0000_0000_0000_0000;
array[1919] <= 16'b0000_0000_0000_0000;
array[1920] <= 16'b0000_0000_0000_0000;
array[1921] <= 16'b0000_0000_0000_0000;
array[1922] <= 16'b0000_0000_0000_0000;
array[1923] <= 16'b0000_0000_0000_0000;
array[1924] <= 16'b0000_0000_0000_0000;
array[1925] <= 16'b0000_0000_0000_0000;
array[1926] <= 16'b0000_0000_0000_0000;
array[1927] <= 16'b0000_0000_0000_0000;
array[1928] <= 16'b0000_0000_0000_0000;
array[1929] <= 16'b0000_0000_0000_0000;
array[1930] <= 16'b0000_0000_0000_0000;
array[1931] <= 16'b0000_0000_0000_0000;
array[1932] <= 16'b0000_0000_0000_0000;
array[1933] <= 16'b0000_0000_0000_0000;
array[1934] <= 16'b0000_0000_0000_0000;
array[1935] <= 16'b0000_0000_0000_0000;
array[1936] <= 16'b0000_0000_0000_0000;
array[1937] <= 16'b0000_0000_0000_0000;
array[1938] <= 16'b0000_0000_0000_0000;
array[1939] <= 16'b0000_0000_0000_0000;
array[1940] <= 16'b0000_0000_0000_0000;
array[1941] <= 16'b0000_0000_0000_0000;
array[1942] <= 16'b0000_0000_0000_0000;
array[1943] <= 16'b0000_0000_0000_0000;
array[1944] <= 16'b0000_0000_0000_0000;
array[1945] <= 16'b0000_0000_0000_0000;
array[1946] <= 16'b0000_0000_0000_0000;
array[1947] <= 16'b0000_0000_0000_0000;
array[1948] <= 16'b0000_0000_0000_0000;
array[1949] <= 16'b0000_0000_0000_0000;
array[1950] <= 16'b0000_0000_0000_0000;
array[1951] <= 16'b0000_0000_0000_0000;
array[1952] <= 16'b0000_0000_0000_0000;
array[1953] <= 16'b0000_0000_0000_0000;
array[1954] <= 16'b0000_0000_0000_0000;
array[1955] <= 16'b0000_0000_0000_0000;
array[1956] <= 16'b0000_0000_0000_0000;
array[1957] <= 16'b0000_0000_0000_0000;
array[1958] <= 16'b0000_0000_0000_0000;
array[1959] <= 16'b0000_0000_0000_0000;
array[1960] <= 16'b0000_0000_0000_0000;
array[1961] <= 16'b0000_0000_0000_0000;
array[1962] <= 16'b0000_0000_0000_0000;
array[1963] <= 16'b0000_0000_0000_0000;
array[1964] <= 16'b0000_0000_0000_0000;
array[1965] <= 16'b0000_0000_0000_0000;
array[1966] <= 16'b0000_0000_0000_0000;
array[1967] <= 16'b0000_0000_0000_0000;
array[1968] <= 16'b0000_0000_0000_0000;
array[1969] <= 16'b0000_0000_0000_0000;
array[1970] <= 16'b0000_0000_0000_0000;
array[1971] <= 16'b0000_0000_0000_0000;
array[1972] <= 16'b0000_0000_0000_0000;
array[1973] <= 16'b0000_0000_0000_0000;
array[1974] <= 16'b0000_0000_0000_0000;
array[1975] <= 16'b0000_0000_0000_0000;
array[1976] <= 16'b0000_0000_0000_0000;
array[1977] <= 16'b0000_0000_0000_0000;
array[1978] <= 16'b0000_0000_0000_0000;
array[1979] <= 16'b0000_0000_0000_0000;
array[1980] <= 16'b0000_0000_0000_0000;
array[1981] <= 16'b0000_0000_0000_0000;
array[1982] <= 16'b0000_0000_0000_0000;
array[1983] <= 16'b0000_0000_0000_0000;
array[1984] <= 16'b0000_0000_0000_0000;
array[1985] <= 16'b0000_0000_0000_0000;
array[1986] <= 16'b0000_0000_0000_0000;
array[1987] <= 16'b0000_0000_0000_0000;
array[1988] <= 16'b0000_0000_0000_0000;
array[1989] <= 16'b0000_0000_0000_0000;
array[1990] <= 16'b0000_0000_0000_0000;
array[1991] <= 16'b0000_0000_0000_0000;
array[1992] <= 16'b0000_0000_0000_0000;
array[1993] <= 16'b0000_0000_0000_0000;
array[1994] <= 16'b0000_0000_0000_0000;
array[1995] <= 16'b0000_0000_0000_0000;
array[1996] <= 16'b0000_0000_0000_0000;
array[1997] <= 16'b0000_0000_0000_0000;
array[1998] <= 16'b0000_0000_0000_0000;
array[1999] <= 16'b0000_0000_0000_0000;
array[2000] <= 16'b0000_0000_0000_0000;
array[2001] <= 16'b0000_0000_0000_0000;
array[2002] <= 16'b0000_0000_0000_0000;
array[2003] <= 16'b0000_0000_0000_0000;
array[2004] <= 16'b0000_0000_0000_0000;
array[2005] <= 16'b0000_0000_0000_0000;
array[2006] <= 16'b0000_0000_0000_0000;
array[2007] <= 16'b0000_0000_0000_0000;
array[2008] <= 16'b0000_0000_0000_0000;
array[2009] <= 16'b0000_0000_0000_0000;
array[2010] <= 16'b0000_0000_0000_0000;
array[2011] <= 16'b0000_0000_0000_0000;
array[2012] <= 16'b0000_0000_0000_0000;
array[2013] <= 16'b0000_0000_0000_0000;
array[2014] <= 16'b0000_0000_0000_0000;
array[2015] <= 16'b0000_0000_0000_0000;
array[2016] <= 16'b0000_0000_0000_0000;
array[2017] <= 16'b0000_0000_0000_0000;
array[2018] <= 16'b0000_0000_0000_0000;
array[2019] <= 16'b0000_0000_0000_0000;
array[2020] <= 16'b0000_0000_0000_0000;
array[2021] <= 16'b0000_0000_0000_0000;
array[2022] <= 16'b0000_0000_0000_0000;
array[2023] <= 16'b0000_0000_0000_0000;
array[2024] <= 16'b0000_0000_0000_0000;
array[2025] <= 16'b0000_0000_0000_0000;
array[2026] <= 16'b0000_0000_0000_0000;
array[2027] <= 16'b0000_0000_0000_0000;
array[2028] <= 16'b0000_0000_0000_0000;
array[2029] <= 16'b0000_0000_0000_0000;
array[2030] <= 16'b0000_0000_0000_0000;
array[2031] <= 16'b0000_0000_0000_0000;
array[2032] <= 16'b0000_0000_0000_0000;
array[2033] <= 16'b0000_0000_0000_0000;
array[2034] <= 16'b0000_0000_0000_0000;
array[2035] <= 16'b0000_0000_0000_0000;
array[2036] <= 16'b0000_0000_0000_0000;
array[2037] <= 16'b0000_0000_0000_0000;
array[2038] <= 16'b0000_0000_0000_0000;
array[2039] <= 16'b0000_0000_0000_0000;
array[2040] <= 16'b0000_0000_0000_0000;
array[2041] <= 16'b0000_0000_0000_0000;
array[2042] <= 16'b0000_0000_0000_0000;
array[2043] <= 16'b0000_0000_0000_0000;
array[2044] <= 16'b0000_0000_0000_0000;
array[2045] <= 16'b0000_0000_0000_0000;
array[2046] <= 16'b0000_0000_0000_0000;
array[2047] <= 16'b0000_0000_0000_0000;
array[2048] <= 16'b0000_0000_0000_0000;
array[2049] <= 16'b0000_0000_0000_0000;
array[2050] <= 16'b0000_0000_0000_0000;
array[2051] <= 16'b0000_0000_0000_0000;
array[2052] <= 16'b0000_0000_0000_0000;
array[2053] <= 16'b0000_0000_0000_0000;
array[2054] <= 16'b0000_0000_0000_0000;
array[2055] <= 16'b0000_0000_0000_0000;
array[2056] <= 16'b0000_0000_0000_0000;
array[2057] <= 16'b0000_0000_0000_0000;
array[2058] <= 16'b0000_0000_0000_0000;
array[2059] <= 16'b0000_0000_0000_0000;
array[2060] <= 16'b0000_0000_0000_0000;
array[2061] <= 16'b0000_0000_0000_0000;
array[2062] <= 16'b0000_0000_0000_0000;
array[2063] <= 16'b0000_0000_0000_0000;
array[2064] <= 16'b0000_0000_0000_0000;
array[2065] <= 16'b0000_0000_0000_0000;
array[2066] <= 16'b0000_0000_0000_0000;
array[2067] <= 16'b0000_0000_0000_0000;
array[2068] <= 16'b0000_0000_0000_0000;
array[2069] <= 16'b0000_0000_0000_0000;
array[2070] <= 16'b0000_0000_0000_0000;
array[2071] <= 16'b0000_0000_0000_0000;
array[2072] <= 16'b0000_0000_0000_0000;
array[2073] <= 16'b0000_0000_0000_0000;
array[2074] <= 16'b0000_0000_0000_0000;
array[2075] <= 16'b0000_0000_0000_0000;
array[2076] <= 16'b0000_0000_0000_0000;
array[2077] <= 16'b0000_0000_0000_0000;
array[2078] <= 16'b0000_0000_0000_0000;
array[2079] <= 16'b0000_0000_0000_0000;
array[2080] <= 16'b0000_0000_0000_0000;
array[2081] <= 16'b0000_0000_0000_0000;
array[2082] <= 16'b0000_0000_0000_0000;
array[2083] <= 16'b0000_0000_0000_0000;
array[2084] <= 16'b0000_0000_0000_0000;
array[2085] <= 16'b0000_0000_0000_0000;
array[2086] <= 16'b0000_0000_0000_0000;
array[2087] <= 16'b0000_0000_0000_0000;
array[2088] <= 16'b0000_0000_0000_0000;
array[2089] <= 16'b0000_0000_0000_0000;
array[2090] <= 16'b0000_0000_0000_0000;
array[2091] <= 16'b0000_0000_0000_0000;
array[2092] <= 16'b0000_0000_0000_0000;
array[2093] <= 16'b0000_0000_0000_0000;
array[2094] <= 16'b0000_0000_0000_0000;
array[2095] <= 16'b0000_0000_0000_0000;
array[2096] <= 16'b0000_0000_0000_0000;
array[2097] <= 16'b0000_0000_0000_0000;
array[2098] <= 16'b0000_0000_0000_0000;
array[2099] <= 16'b0000_0000_0000_0000;
array[2100] <= 16'b0000_0000_0000_0000;
array[2101] <= 16'b0000_0000_0000_0000;
array[2102] <= 16'b0000_0000_0000_0000;
array[2103] <= 16'b0000_0000_0000_0000;
array[2104] <= 16'b0000_0000_0000_0000;
array[2105] <= 16'b0000_0000_0000_0000;
array[2106] <= 16'b0000_0000_0000_0000;
array[2107] <= 16'b0000_0000_0000_0000;
array[2108] <= 16'b0000_0000_0000_0000;
array[2109] <= 16'b0000_0000_0000_0000;
array[2110] <= 16'b0000_0000_0000_0000;
array[2111] <= 16'b0000_0000_0000_0000;
array[2112] <= 16'b0000_0000_0000_0000;
array[2113] <= 16'b0000_0000_0000_0000;
array[2114] <= 16'b0000_0000_0000_0000;
array[2115] <= 16'b0000_0000_0000_0000;
array[2116] <= 16'b0000_0000_0000_0000;
array[2117] <= 16'b0000_0000_0000_0000;
array[2118] <= 16'b0000_0000_0000_0000;
array[2119] <= 16'b0000_0000_0000_0000;
array[2120] <= 16'b0000_0000_0000_0000;
array[2121] <= 16'b0000_0000_0000_0000;
array[2122] <= 16'b0000_0000_0000_0000;
array[2123] <= 16'b0000_0000_0000_0000;
array[2124] <= 16'b0000_0000_0000_0000;
array[2125] <= 16'b0000_0000_0000_0000;
array[2126] <= 16'b0000_0000_0000_0000;
array[2127] <= 16'b0000_0000_0000_0000;
array[2128] <= 16'b0000_0000_0000_0000;
array[2129] <= 16'b0000_0000_0000_0000;
array[2130] <= 16'b0000_0000_0000_0000;
array[2131] <= 16'b0000_0000_0000_0000;
array[2132] <= 16'b0000_0000_0000_0000;
array[2133] <= 16'b0000_0000_0000_0000;
array[2134] <= 16'b0000_0000_0000_0000;
array[2135] <= 16'b0000_0000_0000_0000;
array[2136] <= 16'b0000_0000_0000_0000;
array[2137] <= 16'b0000_0000_0000_0000;
array[2138] <= 16'b0000_0000_0000_0000;
array[2139] <= 16'b0000_0000_0000_0000;
array[2140] <= 16'b0000_0000_0000_0000;
array[2141] <= 16'b0000_0000_0000_0000;
array[2142] <= 16'b0000_0000_0000_0000;
array[2143] <= 16'b0000_0000_0000_0000;
array[2144] <= 16'b0000_0000_0000_0000;
array[2145] <= 16'b0000_0000_0000_0000;
array[2146] <= 16'b0000_0000_0000_0000;
array[2147] <= 16'b0000_0000_0000_0000;
array[2148] <= 16'b0000_0000_0000_0000;
array[2149] <= 16'b0000_0000_0000_0000;
array[2150] <= 16'b0000_0000_0000_0000;
array[2151] <= 16'b0000_0000_0000_0000;
array[2152] <= 16'b0000_0000_0000_0000;
array[2153] <= 16'b0000_0000_0000_0000;
array[2154] <= 16'b0000_0000_0000_0000;
array[2155] <= 16'b0000_0000_0000_0000;
array[2156] <= 16'b0000_0000_0000_0000;
array[2157] <= 16'b0000_0000_0000_0000;
array[2158] <= 16'b0000_0000_0000_0000;
array[2159] <= 16'b0000_0000_0000_0000;
array[2160] <= 16'b0000_0000_0000_0000;
array[2161] <= 16'b0000_0000_0000_0000;
array[2162] <= 16'b0000_0000_0000_0000;
array[2163] <= 16'b0000_0000_0000_0000;
array[2164] <= 16'b0000_0000_0000_0000;
array[2165] <= 16'b0000_0000_0000_0000;
array[2166] <= 16'b0000_0000_0000_0000;
array[2167] <= 16'b0000_0000_0000_0000;
array[2168] <= 16'b0000_0000_0000_0000;
array[2169] <= 16'b0000_0000_0000_0000;
array[2170] <= 16'b0000_0000_0000_0000;
array[2171] <= 16'b0000_0000_0000_0000;
array[2172] <= 16'b0000_0000_0000_0000;
array[2173] <= 16'b0000_0000_0000_0000;
array[2174] <= 16'b0000_0000_0000_0000;
array[2175] <= 16'b0000_0000_0000_0000;
array[2176] <= 16'b0000_0000_0000_0000;
array[2177] <= 16'b0000_0000_0000_0000;
array[2178] <= 16'b0000_0000_0000_0000;
array[2179] <= 16'b0000_0000_0000_0000;
array[2180] <= 16'b0000_0000_0000_0000;
array[2181] <= 16'b0000_0000_0000_0000;
array[2182] <= 16'b0000_0000_0000_0000;
array[2183] <= 16'b0000_0000_0000_0000;
array[2184] <= 16'b0000_0000_0000_0000;
array[2185] <= 16'b0000_0000_0000_0000;
array[2186] <= 16'b0000_0000_0000_0000;
array[2187] <= 16'b0000_0000_0000_0000;
array[2188] <= 16'b0000_0000_0000_0000;
array[2189] <= 16'b0000_0000_0000_0000;
array[2190] <= 16'b0000_0000_0000_0000;
array[2191] <= 16'b0000_0000_0000_0000;
array[2192] <= 16'b0000_0000_0000_0000;
array[2193] <= 16'b0000_0000_0000_0000;
array[2194] <= 16'b0000_0000_0000_0000;
array[2195] <= 16'b0000_0000_0000_0000;
array[2196] <= 16'b0000_0000_0000_0000;
array[2197] <= 16'b0000_0000_0000_0000;
array[2198] <= 16'b0000_0000_0000_0000;
array[2199] <= 16'b0000_0000_0000_0000;
array[2200] <= 16'b0000_0000_0000_0000;
array[2201] <= 16'b0000_0000_0000_0000;
array[2202] <= 16'b0000_0000_0000_0000;
array[2203] <= 16'b0000_0000_0000_0000;
array[2204] <= 16'b0000_0000_0000_0000;
array[2205] <= 16'b0000_0000_0000_0000;
array[2206] <= 16'b0000_0000_0000_0000;
array[2207] <= 16'b0000_0000_0000_0000;
array[2208] <= 16'b0000_0000_0000_0000;
array[2209] <= 16'b0000_0000_0000_0000;
array[2210] <= 16'b0000_0000_0000_0000;
array[2211] <= 16'b0000_0000_0000_0000;
array[2212] <= 16'b0000_0000_0000_0000;
array[2213] <= 16'b0000_0000_0000_0000;
array[2214] <= 16'b0000_0000_0000_0000;
array[2215] <= 16'b0000_0000_0000_0000;
array[2216] <= 16'b0000_0000_0000_0000;
array[2217] <= 16'b0000_0000_0000_0000;
array[2218] <= 16'b0000_0000_0000_0000;
array[2219] <= 16'b0000_0000_0000_0000;
array[2220] <= 16'b0000_0000_0000_0000;
array[2221] <= 16'b0000_0000_0000_0000;
array[2222] <= 16'b0000_0000_0000_0000;
array[2223] <= 16'b0000_0000_0000_0000;
array[2224] <= 16'b0000_0000_0000_0000;
array[2225] <= 16'b0000_0000_0000_0000;
array[2226] <= 16'b0000_0000_0000_0000;
array[2227] <= 16'b0000_0000_0000_0000;
array[2228] <= 16'b0000_0000_0000_0000;
array[2229] <= 16'b0000_0000_0000_0000;
array[2230] <= 16'b0000_0000_0000_0000;
array[2231] <= 16'b0000_0000_0000_0000;
array[2232] <= 16'b0000_0000_0000_0000;
array[2233] <= 16'b0000_0000_0000_0000;
array[2234] <= 16'b0000_0000_0000_0000;
array[2235] <= 16'b0000_0000_0000_0000;
array[2236] <= 16'b0000_0000_0000_0000;
array[2237] <= 16'b0000_0000_0000_0000;
array[2238] <= 16'b0000_0000_0000_0000;
array[2239] <= 16'b0000_0000_0000_0000;
array[2240] <= 16'b0000_0000_0000_0000;
array[2241] <= 16'b0000_0000_0000_0000;
array[2242] <= 16'b0000_0000_0000_0000;
array[2243] <= 16'b0000_0000_0000_0000;
array[2244] <= 16'b0000_0000_0000_0000;
array[2245] <= 16'b0000_0000_0000_0000;
array[2246] <= 16'b0000_0000_0000_0000;
array[2247] <= 16'b0000_0000_0000_0000;
array[2248] <= 16'b0000_0000_0000_0000;
array[2249] <= 16'b0000_0000_0000_0000;
array[2250] <= 16'b0000_0000_0000_0000;
array[2251] <= 16'b0000_0000_0000_0000;
array[2252] <= 16'b0000_0000_0000_0000;
array[2253] <= 16'b0000_0000_0000_0000;
array[2254] <= 16'b0000_0000_0000_0000;
array[2255] <= 16'b0000_0000_0000_0000;
array[2256] <= 16'b0000_0000_0000_0000;
array[2257] <= 16'b0000_0000_0000_0000;
array[2258] <= 16'b0000_0000_0000_0000;
array[2259] <= 16'b0000_0000_0000_0000;
array[2260] <= 16'b0000_0000_0000_0000;
array[2261] <= 16'b0000_0000_0000_0000;
array[2262] <= 16'b0000_0000_0000_0000;
array[2263] <= 16'b0000_0000_0000_0000;
array[2264] <= 16'b0000_0000_0000_0000;
array[2265] <= 16'b0000_0000_0000_0000;
array[2266] <= 16'b0000_0000_0000_0000;
array[2267] <= 16'b0000_0000_0000_0000;
array[2268] <= 16'b0000_0000_0000_0000;
array[2269] <= 16'b0000_0000_0000_0000;
array[2270] <= 16'b0000_0000_0000_0000;
array[2271] <= 16'b0000_0000_0000_0000;
array[2272] <= 16'b0000_0000_0000_0000;
array[2273] <= 16'b0000_0000_0000_0000;
array[2274] <= 16'b0000_0000_0000_0000;
array[2275] <= 16'b0000_0000_0000_0000;
array[2276] <= 16'b0000_0000_0000_0000;
array[2277] <= 16'b0000_0000_0000_0000;
array[2278] <= 16'b0000_0000_0000_0000;
array[2279] <= 16'b0000_0000_0000_0000;
array[2280] <= 16'b0000_0000_0000_0000;
array[2281] <= 16'b0000_0000_0000_0000;
array[2282] <= 16'b0000_0000_0000_0000;
array[2283] <= 16'b0000_0000_0000_0000;
array[2284] <= 16'b0000_0000_0000_0000;
array[2285] <= 16'b0000_0000_0000_0000;
array[2286] <= 16'b0000_0000_0000_0000;
array[2287] <= 16'b0000_0000_0000_0000;
array[2288] <= 16'b0000_0000_0000_0000;
array[2289] <= 16'b0000_0000_0000_0000;
array[2290] <= 16'b0000_0000_0000_0000;
array[2291] <= 16'b0000_0000_0000_0000;
array[2292] <= 16'b0000_0000_0000_0000;
array[2293] <= 16'b0000_0000_0000_0000;
array[2294] <= 16'b0000_0000_0000_0000;
array[2295] <= 16'b0000_0000_0000_0000;
array[2296] <= 16'b0000_0000_0000_0000;
array[2297] <= 16'b0000_0000_0000_0000;
array[2298] <= 16'b0000_0000_0000_0000;
array[2299] <= 16'b0000_0000_0000_0000;
array[2300] <= 16'b0000_0000_0000_0000;
array[2301] <= 16'b0000_0000_0000_0000;
array[2302] <= 16'b0000_0000_0000_0000;
array[2303] <= 16'b0000_0000_0000_0000;
array[2304] <= 16'b0000_0000_0000_0000;
array[2305] <= 16'b0000_0000_0000_0000;
array[2306] <= 16'b0000_0000_0000_0000;
array[2307] <= 16'b0000_0000_0000_0000;
array[2308] <= 16'b0000_0000_0000_0000;
array[2309] <= 16'b0000_0000_0000_0000;
array[2310] <= 16'b0000_0000_0000_0000;
array[2311] <= 16'b0000_0000_0000_0000;
array[2312] <= 16'b0000_0000_0000_0000;
array[2313] <= 16'b0000_0000_0000_0000;
array[2314] <= 16'b0000_0000_0000_0000;
array[2315] <= 16'b0000_0000_0000_0000;
array[2316] <= 16'b0000_0000_0000_0000;
array[2317] <= 16'b0000_0000_0000_0000;
array[2318] <= 16'b0000_0000_0000_0000;
array[2319] <= 16'b0000_0000_0000_0000;
array[2320] <= 16'b0000_0000_0000_0000;
array[2321] <= 16'b0000_0000_0000_0000;
array[2322] <= 16'b0000_0000_0000_0000;
array[2323] <= 16'b0000_0000_0000_0000;
array[2324] <= 16'b0000_0000_0000_0000;
array[2325] <= 16'b0000_0000_0000_0000;
array[2326] <= 16'b0000_0000_0000_0000;
array[2327] <= 16'b0000_0000_0000_0000;
array[2328] <= 16'b0000_0000_0000_0000;
array[2329] <= 16'b0000_0000_0000_0000;
array[2330] <= 16'b0000_0000_0000_0000;
array[2331] <= 16'b0000_0000_0000_0000;
array[2332] <= 16'b0000_0000_0000_0000;
array[2333] <= 16'b0000_0000_0000_0000;
array[2334] <= 16'b0000_0000_0000_0000;
array[2335] <= 16'b0000_0000_0000_0000;
array[2336] <= 16'b0000_0000_0000_0000;
array[2337] <= 16'b0000_0000_0000_0000;
array[2338] <= 16'b0000_0000_0000_0000;
array[2339] <= 16'b0000_0000_0000_0000;
array[2340] <= 16'b0000_0000_0000_0000;
array[2341] <= 16'b0000_0000_0000_0000;
array[2342] <= 16'b0000_0000_0000_0000;
array[2343] <= 16'b0000_0000_0000_0000;
array[2344] <= 16'b0000_0000_0000_0000;
array[2345] <= 16'b0000_0000_0000_0000;
array[2346] <= 16'b0000_0000_0000_0000;
array[2347] <= 16'b0000_0000_0000_0000;
array[2348] <= 16'b0000_0000_0000_0000;
array[2349] <= 16'b0000_0000_0000_0000;
array[2350] <= 16'b0000_0000_0000_0000;
array[2351] <= 16'b0000_0000_0000_0000;
array[2352] <= 16'b0000_0000_0000_0000;
array[2353] <= 16'b0000_0000_0000_0000;
array[2354] <= 16'b0000_0000_0000_0000;
array[2355] <= 16'b0000_0000_0000_0000;
array[2356] <= 16'b0000_0000_0000_0000;
array[2357] <= 16'b0000_0000_0000_0000;
array[2358] <= 16'b0000_0000_0000_0000;
array[2359] <= 16'b0000_0000_0000_0000;
array[2360] <= 16'b0000_0000_0000_0000;
array[2361] <= 16'b0000_0000_0000_0000;
array[2362] <= 16'b0000_0000_0000_0000;
array[2363] <= 16'b0000_0000_0000_0000;
array[2364] <= 16'b0000_0000_0000_0000;
array[2365] <= 16'b0000_0000_0000_0000;
array[2366] <= 16'b0000_0000_0000_0000;
array[2367] <= 16'b0000_0000_0000_0000;
array[2368] <= 16'b0000_0000_0000_0000;
array[2369] <= 16'b0000_0000_0000_0000;
array[2370] <= 16'b0000_0000_0000_0000;
array[2371] <= 16'b0000_0000_0000_0000;
array[2372] <= 16'b0000_0000_0000_0000;
array[2373] <= 16'b0000_0000_0000_0000;
array[2374] <= 16'b0000_0000_0000_0000;
array[2375] <= 16'b0000_0000_0000_0000;
array[2376] <= 16'b0000_0000_0000_0000;
array[2377] <= 16'b0000_0000_0000_0000;
array[2378] <= 16'b0000_0000_0000_0000;
array[2379] <= 16'b0000_0000_0000_0000;
array[2380] <= 16'b0000_0000_0000_0000;
array[2381] <= 16'b0000_0000_0000_0000;
array[2382] <= 16'b0000_0000_0000_0000;
array[2383] <= 16'b0000_0000_0000_0000;
array[2384] <= 16'b0000_0000_0000_0000;
array[2385] <= 16'b0000_0000_0000_0000;
array[2386] <= 16'b0000_0000_0000_0000;
array[2387] <= 16'b0000_0000_0000_0000;
array[2388] <= 16'b0000_0000_0000_0000;
array[2389] <= 16'b0000_0000_0000_0000;
array[2390] <= 16'b0000_0000_0000_0000;
array[2391] <= 16'b0000_0000_0000_0000;
array[2392] <= 16'b0000_0000_0000_0000;
array[2393] <= 16'b0000_0000_0000_0000;
array[2394] <= 16'b0000_0000_0000_0000;
array[2395] <= 16'b0000_0000_0000_0000;
array[2396] <= 16'b0000_0000_0000_0000;
array[2397] <= 16'b0000_0000_0000_0000;
array[2398] <= 16'b0000_0000_0000_0000;
array[2399] <= 16'b0000_0000_0000_0000;
array[2400] <= 16'b0000_0000_0000_0000;
array[2401] <= 16'b0000_0000_0000_0000;
array[2402] <= 16'b0000_0000_0000_0000;
array[2403] <= 16'b0000_0000_0000_0000;
array[2404] <= 16'b0000_0000_0000_0000;
array[2405] <= 16'b0000_0000_0000_0000;
array[2406] <= 16'b0000_0000_0000_0000;
array[2407] <= 16'b0000_0000_0000_0000;
array[2408] <= 16'b0000_0000_0000_0000;
array[2409] <= 16'b0000_0000_0000_0000;
array[2410] <= 16'b0000_0000_0000_0000;
array[2411] <= 16'b0000_0000_0000_0000;
array[2412] <= 16'b0000_0000_0000_0000;
array[2413] <= 16'b0000_0000_0000_0000;
array[2414] <= 16'b0000_0000_0000_0000;
array[2415] <= 16'b0000_0000_0000_0000;
array[2416] <= 16'b0000_0000_0000_0000;
array[2417] <= 16'b0000_0000_0000_0000;
array[2418] <= 16'b0000_0000_0000_0000;
array[2419] <= 16'b0000_0000_0000_0000;
array[2420] <= 16'b0000_0000_0000_0000;
array[2421] <= 16'b0000_0000_0000_0000;
array[2422] <= 16'b0000_0000_0000_0000;
array[2423] <= 16'b0000_0000_0000_0000;
array[2424] <= 16'b0000_0000_0000_0000;
array[2425] <= 16'b0000_0000_0000_0000;
array[2426] <= 16'b0000_0000_0000_0000;
array[2427] <= 16'b0000_0000_0000_0000;
array[2428] <= 16'b0000_0000_0000_0000;
array[2429] <= 16'b0000_0000_0000_0000;
array[2430] <= 16'b0000_0000_0000_0000;
array[2431] <= 16'b0000_0000_0000_0000;
array[2432] <= 16'b0000_0000_0000_0000;
array[2433] <= 16'b0000_0000_0000_0000;
array[2434] <= 16'b0000_0000_0000_0000;
array[2435] <= 16'b0000_0000_0000_0000;
array[2436] <= 16'b0000_0000_0000_0000;
array[2437] <= 16'b0000_0000_0000_0000;
array[2438] <= 16'b0000_0000_0000_0000;
array[2439] <= 16'b0000_0000_0000_0000;
array[2440] <= 16'b0000_0000_0000_0000;
array[2441] <= 16'b0000_0000_0000_0000;
array[2442] <= 16'b0000_0000_0000_0000;
array[2443] <= 16'b0000_0000_0000_0000;
array[2444] <= 16'b0000_0000_0000_0000;
array[2445] <= 16'b0000_0000_0000_0000;
array[2446] <= 16'b0000_0000_0000_0000;
array[2447] <= 16'b0000_0000_0000_0000;
array[2448] <= 16'b0000_0000_0000_0000;
array[2449] <= 16'b0000_0000_0000_0000;
array[2450] <= 16'b0000_0000_0000_0000;
array[2451] <= 16'b0000_0000_0000_0000;
array[2452] <= 16'b0000_0000_0000_0000;
array[2453] <= 16'b0000_0000_0000_0000;
array[2454] <= 16'b0000_0000_0000_0000;
array[2455] <= 16'b0000_0000_0000_0000;
array[2456] <= 16'b0000_0000_0000_0000;
array[2457] <= 16'b0000_0000_0000_0000;
array[2458] <= 16'b0000_0000_0000_0000;
array[2459] <= 16'b0000_0000_0000_0000;
array[2460] <= 16'b0000_0000_0000_0000;
array[2461] <= 16'b0000_0000_0000_0000;
array[2462] <= 16'b0000_0000_0000_0000;
array[2463] <= 16'b0000_0000_0000_0000;
array[2464] <= 16'b0000_0000_0000_0000;
array[2465] <= 16'b0000_0000_0000_0000;
array[2466] <= 16'b0000_0000_0000_0000;
array[2467] <= 16'b0000_0000_0000_0000;
array[2468] <= 16'b0000_0000_0000_0000;
array[2469] <= 16'b0000_0000_0000_0000;
array[2470] <= 16'b0000_0000_0000_0000;
array[2471] <= 16'b0000_0000_0000_0000;
array[2472] <= 16'b0000_0000_0000_0000;
array[2473] <= 16'b0000_0000_0000_0000;
array[2474] <= 16'b0000_0000_0000_0000;
array[2475] <= 16'b0000_0000_0000_0000;
array[2476] <= 16'b0000_0000_0000_0000;
array[2477] <= 16'b0000_0000_0000_0000;
array[2478] <= 16'b0000_0000_0000_0000;
array[2479] <= 16'b0000_0000_0000_0000;
array[2480] <= 16'b0000_0000_0000_0000;
array[2481] <= 16'b0000_0000_0000_0000;
array[2482] <= 16'b0000_0000_0000_0000;
array[2483] <= 16'b0000_0000_0000_0000;
array[2484] <= 16'b0000_0000_0000_0000;
array[2485] <= 16'b0000_0000_0000_0000;
array[2486] <= 16'b0000_0000_0000_0000;
array[2487] <= 16'b0000_0000_0000_0000;
array[2488] <= 16'b0000_0000_0000_0000;
array[2489] <= 16'b0000_0000_0000_0000;
array[2490] <= 16'b0000_0000_0000_0000;
array[2491] <= 16'b0000_0000_0000_0000;
array[2492] <= 16'b0000_0000_0000_0000;
array[2493] <= 16'b0000_0000_0000_0000;
array[2494] <= 16'b0000_0000_0000_0000;
array[2495] <= 16'b0000_0000_0000_0000;
array[2496] <= 16'b0000_0000_0000_0000;
array[2497] <= 16'b0000_0000_0000_0000;
array[2498] <= 16'b0000_0000_0000_0000;
array[2499] <= 16'b0000_0000_0000_0000;
array[2500] <= 16'b0000_0000_0000_0000;
array[2501] <= 16'b0000_0000_0000_0000;
array[2502] <= 16'b0000_0000_0000_0000;
array[2503] <= 16'b0000_0000_0000_0000;
array[2504] <= 16'b0000_0000_0000_0000;
array[2505] <= 16'b0000_0000_0000_0000;
array[2506] <= 16'b0000_0000_0000_0000;
array[2507] <= 16'b0000_0000_0000_0000;
array[2508] <= 16'b0000_0000_0000_0000;
array[2509] <= 16'b0000_0000_0000_0000;
array[2510] <= 16'b0000_0000_0000_0000;
array[2511] <= 16'b0000_0000_0000_0000;
array[2512] <= 16'b0000_0000_0000_0000;
array[2513] <= 16'b0000_0000_0000_0000;
array[2514] <= 16'b0000_0000_0000_0000;
array[2515] <= 16'b0000_0000_0000_0000;
array[2516] <= 16'b0000_0000_0000_0000;
array[2517] <= 16'b0000_0000_0000_0000;
array[2518] <= 16'b0000_0000_0000_0000;
array[2519] <= 16'b0000_0000_0000_0000;
array[2520] <= 16'b0000_0000_0000_0000;
array[2521] <= 16'b0000_0000_0000_0000;
array[2522] <= 16'b0000_0000_0000_0000;
array[2523] <= 16'b0000_0000_0000_0000;
array[2524] <= 16'b0000_0000_0000_0000;
array[2525] <= 16'b0000_0000_0000_0000;
array[2526] <= 16'b0000_0000_0000_0000;
array[2527] <= 16'b0000_0000_0000_0000;
array[2528] <= 16'b0000_0000_0000_0000;
array[2529] <= 16'b0000_0000_0000_0000;
array[2530] <= 16'b0000_0000_0000_0000;
array[2531] <= 16'b0000_0000_0000_0000;
array[2532] <= 16'b0000_0000_0000_0000;
array[2533] <= 16'b0000_0000_0000_0000;
array[2534] <= 16'b0000_0000_0000_0000;
array[2535] <= 16'b0000_0000_0000_0000;
array[2536] <= 16'b0000_0000_0000_0000;
array[2537] <= 16'b0000_0000_0000_0000;
array[2538] <= 16'b0000_0000_0000_0000;
array[2539] <= 16'b0000_0000_0000_0000;
array[2540] <= 16'b0000_0000_0000_0000;
array[2541] <= 16'b0000_0000_0000_0000;
array[2542] <= 16'b0000_0000_0000_0000;
array[2543] <= 16'b0000_0000_0000_0000;
array[2544] <= 16'b0000_0000_0000_0000;
array[2545] <= 16'b0000_0000_0000_0000;
array[2546] <= 16'b0000_0000_0000_0000;
array[2547] <= 16'b0000_0000_0000_0000;
array[2548] <= 16'b0000_0000_0000_0000;
array[2549] <= 16'b0000_0000_0000_0000;
array[2550] <= 16'b0000_0000_0000_0000;
array[2551] <= 16'b0000_0000_0000_0000;
array[2552] <= 16'b0000_0000_0000_0000;
array[2553] <= 16'b0000_0000_0000_0000;
array[2554] <= 16'b0000_0000_0000_0000;
array[2555] <= 16'b0000_0000_0000_0000;
array[2556] <= 16'b0000_0000_0000_0000;
array[2557] <= 16'b0000_0000_0000_0000;
array[2558] <= 16'b0000_0000_0000_0000;
array[2559] <= 16'b0000_0000_0000_0000;
array[2560] <= 16'b0000_0000_0000_0000;
array[2561] <= 16'b0000_0000_0000_0000;
array[2562] <= 16'b0000_0000_0000_0000;
array[2563] <= 16'b0000_0000_0000_0000;
array[2564] <= 16'b0000_0000_0000_0000;
array[2565] <= 16'b0000_0000_0000_0000;
array[2566] <= 16'b0000_0000_0000_0000;
array[2567] <= 16'b0000_0000_0000_0000;
array[2568] <= 16'b0000_0000_0000_0000;
array[2569] <= 16'b0000_0000_0000_0000;
array[2570] <= 16'b0000_0000_0000_0000;
array[2571] <= 16'b0000_0000_0000_0000;
array[2572] <= 16'b0000_0000_0000_0000;
array[2573] <= 16'b0000_0000_0000_0000;
array[2574] <= 16'b0000_0000_0000_0000;
array[2575] <= 16'b0000_0000_0000_0000;
array[2576] <= 16'b0000_0000_0000_0000;
array[2577] <= 16'b0000_0000_0000_0000;
array[2578] <= 16'b0000_0000_0000_0000;
array[2579] <= 16'b0000_0000_0000_0000;
array[2580] <= 16'b0000_0000_0000_0000;
array[2581] <= 16'b0000_0000_0000_0000;
array[2582] <= 16'b0000_0000_0000_0000;
array[2583] <= 16'b0000_0000_0000_0000;
array[2584] <= 16'b0000_0000_0000_0000;
array[2585] <= 16'b0000_0000_0000_0000;
array[2586] <= 16'b0000_0000_0000_0000;
array[2587] <= 16'b0000_0000_0000_0000;
array[2588] <= 16'b0000_0000_0000_0000;
array[2589] <= 16'b0000_0000_0000_0000;
array[2590] <= 16'b0000_0000_0000_0000;
array[2591] <= 16'b0000_0000_0000_0000;
array[2592] <= 16'b0000_0000_0000_0000;
array[2593] <= 16'b0000_0000_0000_0000;
array[2594] <= 16'b0000_0000_0000_0000;
array[2595] <= 16'b0000_0000_0000_0000;
array[2596] <= 16'b0000_0000_0000_0000;
array[2597] <= 16'b0000_0000_0000_0000;
array[2598] <= 16'b0000_0000_0000_0000;
array[2599] <= 16'b0000_0000_0000_0000;
array[2600] <= 16'b0000_0000_0000_0000;
array[2601] <= 16'b0000_0000_0000_0000;
array[2602] <= 16'b0000_0000_0000_0000;
array[2603] <= 16'b0000_0000_0000_0000;
array[2604] <= 16'b0000_0000_0000_0000;
array[2605] <= 16'b0000_0000_0000_0000;
array[2606] <= 16'b0000_0000_0000_0000;
array[2607] <= 16'b0000_0000_0000_0000;
array[2608] <= 16'b0000_0000_0000_0000;
array[2609] <= 16'b0000_0000_0000_0000;
array[2610] <= 16'b0000_0000_0000_0000;
array[2611] <= 16'b0000_0000_0000_0000;
array[2612] <= 16'b0000_0000_0000_0000;
array[2613] <= 16'b0000_0000_0000_0000;
array[2614] <= 16'b0000_0000_0000_0000;
array[2615] <= 16'b0000_0000_0000_0000;
array[2616] <= 16'b0000_0000_0000_0000;
array[2617] <= 16'b0000_0000_0000_0000;
array[2618] <= 16'b0000_0000_0000_0000;
array[2619] <= 16'b0000_0000_0000_0000;
array[2620] <= 16'b0000_0000_0000_0000;
array[2621] <= 16'b0000_0000_0000_0000;
array[2622] <= 16'b0000_0000_0000_0000;
array[2623] <= 16'b0000_0000_0000_0000;
array[2624] <= 16'b0000_0000_0000_0000;
array[2625] <= 16'b0000_0000_0000_0000;
array[2626] <= 16'b0000_0000_0000_0000;
array[2627] <= 16'b0000_0000_0000_0000;
array[2628] <= 16'b0000_0000_0000_0000;
array[2629] <= 16'b0000_0000_0000_0000;
array[2630] <= 16'b0000_0000_0000_0000;
array[2631] <= 16'b0000_0000_0000_0000;
array[2632] <= 16'b0000_0000_0000_0000;
array[2633] <= 16'b0000_0000_0000_0000;
array[2634] <= 16'b0000_0000_0000_0000;
array[2635] <= 16'b0000_0000_0000_0000;
array[2636] <= 16'b0000_0000_0000_0000;
array[2637] <= 16'b0000_0000_0000_0000;
array[2638] <= 16'b0000_0000_0000_0000;
array[2639] <= 16'b0000_0000_0000_0000;
array[2640] <= 16'b0000_0000_0000_0000;
array[2641] <= 16'b0000_0000_0000_0000;
array[2642] <= 16'b0000_0000_0000_0000;
array[2643] <= 16'b0000_0000_0000_0000;
array[2644] <= 16'b0000_0000_0000_0000;
array[2645] <= 16'b0000_0000_0000_0000;
array[2646] <= 16'b0000_0000_0000_0000;
array[2647] <= 16'b0000_0000_0000_0000;
array[2648] <= 16'b0000_0000_0000_0000;
array[2649] <= 16'b0000_0000_0000_0000;
array[2650] <= 16'b0000_0000_0000_0000;
array[2651] <= 16'b0000_0000_0000_0000;
array[2652] <= 16'b0000_0000_0000_0000;
array[2653] <= 16'b0000_0000_0000_0000;
array[2654] <= 16'b0000_0000_0000_0000;
array[2655] <= 16'b0000_0000_0000_0000;
array[2656] <= 16'b0000_0000_0000_0000;
array[2657] <= 16'b0000_0000_0000_0000;
array[2658] <= 16'b0000_0000_0000_0000;
array[2659] <= 16'b0000_0000_0000_0000;
array[2660] <= 16'b0000_0000_0000_0000;
array[2661] <= 16'b0000_0000_0000_0000;
array[2662] <= 16'b0000_0000_0000_0000;
array[2663] <= 16'b0000_0000_0000_0000;
array[2664] <= 16'b0000_0000_0000_0000;
array[2665] <= 16'b0000_0000_0000_0000;
array[2666] <= 16'b0000_0000_0000_0000;
array[2667] <= 16'b0000_0000_0000_0000;
array[2668] <= 16'b0000_0000_0000_0000;
array[2669] <= 16'b0000_0000_0000_0000;
array[2670] <= 16'b0000_0000_0000_0000;
array[2671] <= 16'b0000_0000_0000_0000;
array[2672] <= 16'b0000_0000_0000_0000;
array[2673] <= 16'b0000_0000_0000_0000;
array[2674] <= 16'b0000_0000_0000_0000;
array[2675] <= 16'b0000_0000_0000_0000;
array[2676] <= 16'b0000_0000_0000_0000;
array[2677] <= 16'b0000_0000_0000_0000;
array[2678] <= 16'b0000_0000_0000_0000;
array[2679] <= 16'b0000_0000_0000_0000;
array[2680] <= 16'b0000_0000_0000_0000;
array[2681] <= 16'b0000_0000_0000_0000;
array[2682] <= 16'b0000_0000_0000_0000;
array[2683] <= 16'b0000_0000_0000_0000;
array[2684] <= 16'b0000_0000_0000_0000;
array[2685] <= 16'b0000_0000_0000_0000;
array[2686] <= 16'b0000_0000_0000_0000;
array[2687] <= 16'b0000_0000_0000_0000;
array[2688] <= 16'b0000_0000_0000_0000;
array[2689] <= 16'b0000_0000_0000_0000;
array[2690] <= 16'b0000_0000_0000_0000;
array[2691] <= 16'b0000_0000_0000_0000;
array[2692] <= 16'b0000_0000_0000_0000;
array[2693] <= 16'b0000_0000_0000_0000;
array[2694] <= 16'b0000_0000_0000_0000;
array[2695] <= 16'b0000_0000_0000_0000;
array[2696] <= 16'b0000_0000_0000_0000;
array[2697] <= 16'b0000_0000_0000_0000;
array[2698] <= 16'b0000_0000_0000_0000;
array[2699] <= 16'b0000_0000_0000_0000;
array[2700] <= 16'b0000_0000_0000_0000;
array[2701] <= 16'b0000_0000_0000_0000;
array[2702] <= 16'b0000_0000_0000_0000;
array[2703] <= 16'b0000_0000_0000_0000;
array[2704] <= 16'b0000_0000_0000_0000;
array[2705] <= 16'b0000_0000_0000_0000;
array[2706] <= 16'b0000_0000_0000_0000;
array[2707] <= 16'b0000_0000_0000_0000;
array[2708] <= 16'b0000_0000_0000_0000;
array[2709] <= 16'b0000_0000_0000_0000;
array[2710] <= 16'b0000_0000_0000_0000;
array[2711] <= 16'b0000_0000_0000_0000;
array[2712] <= 16'b0000_0000_0000_0000;
array[2713] <= 16'b0000_0000_0000_0000;
array[2714] <= 16'b0000_0000_0000_0000;
array[2715] <= 16'b0000_0000_0000_0000;
array[2716] <= 16'b0000_0000_0000_0000;
array[2717] <= 16'b0000_0000_0000_0000;
array[2718] <= 16'b0000_0000_0000_0000;
array[2719] <= 16'b0000_0000_0000_0000;
array[2720] <= 16'b0000_0000_0000_0000;
array[2721] <= 16'b0000_0000_0000_0000;
array[2722] <= 16'b0000_0000_0000_0000;
array[2723] <= 16'b0000_0000_0000_0000;
array[2724] <= 16'b0000_0000_0000_0000;
array[2725] <= 16'b0000_0000_0000_0000;
array[2726] <= 16'b0000_0000_0000_0000;
array[2727] <= 16'b0000_0000_0000_0000;
array[2728] <= 16'b0000_0000_0000_0000;
array[2729] <= 16'b0000_0000_0000_0000;
array[2730] <= 16'b0000_0000_0000_0000;
array[2731] <= 16'b0000_0000_0000_0000;
array[2732] <= 16'b0000_0000_0000_0000;
array[2733] <= 16'b0000_0000_0000_0000;
array[2734] <= 16'b0000_0000_0000_0000;
array[2735] <= 16'b0000_0000_0000_0000;
array[2736] <= 16'b0000_0000_0000_0000;
array[2737] <= 16'b0000_0000_0000_0000;
array[2738] <= 16'b0000_0000_0000_0000;
array[2739] <= 16'b0000_0000_0000_0000;
array[2740] <= 16'b0000_0000_0000_0000;
array[2741] <= 16'b0000_0000_0000_0000;
array[2742] <= 16'b0000_0000_0000_0000;
array[2743] <= 16'b0000_0000_0000_0000;
array[2744] <= 16'b0000_0000_0000_0000;
array[2745] <= 16'b0000_0000_0000_0000;
array[2746] <= 16'b0000_0000_0000_0000;
array[2747] <= 16'b0000_0000_0000_0000;
array[2748] <= 16'b0000_0000_0000_0000;
array[2749] <= 16'b0000_0000_0000_0000;
array[2750] <= 16'b0000_0000_0000_0000;
array[2751] <= 16'b0000_0000_0000_0000;
array[2752] <= 16'b0000_0000_0000_0000;
array[2753] <= 16'b0000_0000_0000_0000;
array[2754] <= 16'b0000_0000_0000_0000;
array[2755] <= 16'b0000_0000_0000_0000;
array[2756] <= 16'b0000_0000_0000_0000;
array[2757] <= 16'b0000_0000_0000_0000;
array[2758] <= 16'b0000_0000_0000_0000;
array[2759] <= 16'b0000_0000_0000_0000;
array[2760] <= 16'b0000_0000_0000_0000;
array[2761] <= 16'b0000_0000_0000_0000;
array[2762] <= 16'b0000_0000_0000_0000;
array[2763] <= 16'b0000_0000_0000_0000;
array[2764] <= 16'b0000_0000_0000_0000;
array[2765] <= 16'b0000_0000_0000_0000;
array[2766] <= 16'b0000_0000_0000_0000;
array[2767] <= 16'b0000_0000_0000_0000;
array[2768] <= 16'b0000_0000_0000_0000;
array[2769] <= 16'b0000_0000_0000_0000;
array[2770] <= 16'b0000_0000_0000_0000;
array[2771] <= 16'b0000_0000_0000_0000;
array[2772] <= 16'b0000_0000_0000_0000;
array[2773] <= 16'b0000_0000_0000_0000;
array[2774] <= 16'b0000_0000_0000_0000;
array[2775] <= 16'b0000_0000_0000_0000;
array[2776] <= 16'b0000_0000_0000_0000;
array[2777] <= 16'b0000_0000_0000_0000;
array[2778] <= 16'b0000_0000_0000_0000;
array[2779] <= 16'b0000_0000_0000_0000;
array[2780] <= 16'b0000_0000_0000_0000;
array[2781] <= 16'b0000_0000_0000_0000;
array[2782] <= 16'b0000_0000_0000_0000;
array[2783] <= 16'b0000_0000_0000_0000;
array[2784] <= 16'b0000_0000_0000_0000;
array[2785] <= 16'b0000_0000_0000_0000;
array[2786] <= 16'b0000_0000_0000_0000;
array[2787] <= 16'b0000_0000_0000_0000;
array[2788] <= 16'b0000_0000_0000_0000;
array[2789] <= 16'b0000_0000_0000_0000;
array[2790] <= 16'b0000_0000_0000_0000;
array[2791] <= 16'b0000_0000_0000_0000;
array[2792] <= 16'b0000_0000_0000_0000;
array[2793] <= 16'b0000_0000_0000_0000;
array[2794] <= 16'b0000_0000_0000_0000;
array[2795] <= 16'b0000_0000_0000_0000;
array[2796] <= 16'b0000_0000_0000_0000;
array[2797] <= 16'b0000_0000_0000_0000;
array[2798] <= 16'b0000_0000_0000_0000;
array[2799] <= 16'b0000_0000_0000_0000;
array[2800] <= 16'b0000_0000_0000_0000;
array[2801] <= 16'b0000_0000_0000_0000;
array[2802] <= 16'b0000_0000_0000_0000;
array[2803] <= 16'b0000_0000_0000_0000;
array[2804] <= 16'b0000_0000_0000_0000;
array[2805] <= 16'b0000_0000_0000_0000;
array[2806] <= 16'b0000_0000_0000_0000;
array[2807] <= 16'b0000_0000_0000_0000;
array[2808] <= 16'b0000_0000_0000_0000;
array[2809] <= 16'b0000_0000_0000_0000;
array[2810] <= 16'b0000_0000_0000_0000;
array[2811] <= 16'b0000_0000_0000_0000;
array[2812] <= 16'b0000_0000_0000_0000;
array[2813] <= 16'b0000_0000_0000_0000;
array[2814] <= 16'b0000_0000_0000_0000;
array[2815] <= 16'b0000_0000_0000_0000;
array[2816] <= 16'b0000_0000_0000_0000;
array[2817] <= 16'b0000_0000_0000_0000;
array[2818] <= 16'b0000_0000_0000_0000;
array[2819] <= 16'b0000_0000_0000_0000;
array[2820] <= 16'b0000_0000_0000_0000;
array[2821] <= 16'b0000_0000_0000_0000;
array[2822] <= 16'b0000_0000_0000_0000;
array[2823] <= 16'b0000_0000_0000_0000;
array[2824] <= 16'b0000_0000_0000_0000;
array[2825] <= 16'b0000_0000_0000_0000;
array[2826] <= 16'b0000_0000_0000_0000;
array[2827] <= 16'b0000_0000_0000_0000;
array[2828] <= 16'b0000_0000_0000_0000;
array[2829] <= 16'b0000_0000_0000_0000;
array[2830] <= 16'b0000_0000_0000_0000;
array[2831] <= 16'b0000_0000_0000_0000;
array[2832] <= 16'b0000_0000_0000_0000;
array[2833] <= 16'b0000_0000_0000_0000;
array[2834] <= 16'b0000_0000_0000_0000;
array[2835] <= 16'b0000_0000_0000_0000;
array[2836] <= 16'b0000_0000_0000_0000;
array[2837] <= 16'b0000_0000_0000_0000;
array[2838] <= 16'b0000_0000_0000_0000;
array[2839] <= 16'b0000_0000_0000_0000;
array[2840] <= 16'b0000_0000_0000_0000;
array[2841] <= 16'b0000_0000_0000_0000;
array[2842] <= 16'b0000_0000_0000_0000;
array[2843] <= 16'b0000_0000_0000_0000;
array[2844] <= 16'b0000_0000_0000_0000;
array[2845] <= 16'b0000_0000_0000_0000;
array[2846] <= 16'b0000_0000_0000_0000;
array[2847] <= 16'b0000_0000_0000_0000;
array[2848] <= 16'b0000_0000_0000_0000;
array[2849] <= 16'b0000_0000_0000_0000;
array[2850] <= 16'b0000_0000_0000_0000;
array[2851] <= 16'b0000_0000_0000_0000;
array[2852] <= 16'b0000_0000_0000_0000;
array[2853] <= 16'b0000_0000_0000_0000;
array[2854] <= 16'b0000_0000_0000_0000;
array[2855] <= 16'b0000_0000_0000_0000;
array[2856] <= 16'b0000_0000_0000_0000;
array[2857] <= 16'b0000_0000_0000_0000;
array[2858] <= 16'b0000_0000_0000_0000;
array[2859] <= 16'b0000_0000_0000_0000;
array[2860] <= 16'b0000_0000_0000_0000;
array[2861] <= 16'b0000_0000_0000_0000;
array[2862] <= 16'b0000_0000_0000_0000;
array[2863] <= 16'b0000_0000_0000_0000;
array[2864] <= 16'b0000_0000_0000_0000;
array[2865] <= 16'b0000_0000_0000_0000;
array[2866] <= 16'b0000_0000_0000_0000;
array[2867] <= 16'b0000_0000_0000_0000;
array[2868] <= 16'b0000_0000_0000_0000;
array[2869] <= 16'b0000_0000_0000_0000;
array[2870] <= 16'b0000_0000_0000_0000;
array[2871] <= 16'b0000_0000_0000_0000;
array[2872] <= 16'b0000_0000_0000_0000;
array[2873] <= 16'b0000_0000_0000_0000;
array[2874] <= 16'b0000_0000_0000_0000;
array[2875] <= 16'b0000_0000_0000_0000;
array[2876] <= 16'b0000_0000_0000_0000;
array[2877] <= 16'b0000_0000_0000_0000;
array[2878] <= 16'b0000_0000_0000_0000;
array[2879] <= 16'b0000_0000_0000_0000;
array[2880] <= 16'b0000_0000_0000_0000;
array[2881] <= 16'b0000_0000_0000_0000;
array[2882] <= 16'b0000_0000_0000_0000;
array[2883] <= 16'b0000_0000_0000_0000;
array[2884] <= 16'b0000_0000_0000_0000;
array[2885] <= 16'b0000_0000_0000_0000;
array[2886] <= 16'b0000_0000_0000_0000;
array[2887] <= 16'b0000_0000_0000_0000;
array[2888] <= 16'b0000_0000_0000_0000;
array[2889] <= 16'b0000_0000_0000_0000;
array[2890] <= 16'b0000_0000_0000_0000;
array[2891] <= 16'b0000_0000_0000_0000;
array[2892] <= 16'b0000_0000_0000_0000;
array[2893] <= 16'b0000_0000_0000_0000;
array[2894] <= 16'b0000_0000_0000_0000;
array[2895] <= 16'b0000_0000_0000_0000;
array[2896] <= 16'b0000_0000_0000_0000;
array[2897] <= 16'b0000_0000_0000_0000;
array[2898] <= 16'b0000_0000_0000_0000;
array[2899] <= 16'b0000_0000_0000_0000;
array[2900] <= 16'b0000_0000_0000_0000;
array[2901] <= 16'b0000_0000_0000_0000;
array[2902] <= 16'b0000_0000_0000_0000;
array[2903] <= 16'b0000_0000_0000_0000;
array[2904] <= 16'b0000_0000_0000_0000;
array[2905] <= 16'b0000_0000_0000_0000;
array[2906] <= 16'b0000_0000_0000_0000;
array[2907] <= 16'b0000_0000_0000_0000;
array[2908] <= 16'b0000_0000_0000_0000;
array[2909] <= 16'b0000_0000_0000_0000;
array[2910] <= 16'b0000_0000_0000_0000;
array[2911] <= 16'b0000_0000_0000_0000;
array[2912] <= 16'b0000_0000_0000_0000;
array[2913] <= 16'b0000_0000_0000_0000;
array[2914] <= 16'b0000_0000_0000_0000;
array[2915] <= 16'b0000_0000_0000_0000;
array[2916] <= 16'b0000_0000_0000_0000;
array[2917] <= 16'b0000_0000_0000_0000;
array[2918] <= 16'b0000_0000_0000_0000;
array[2919] <= 16'b0000_0000_0000_0000;
array[2920] <= 16'b0000_0000_0000_0000;
array[2921] <= 16'b0000_0000_0000_0000;
array[2922] <= 16'b0000_0000_0000_0000;
array[2923] <= 16'b0000_0000_0000_0000;
array[2924] <= 16'b0000_0000_0000_0000;
array[2925] <= 16'b0000_0000_0000_0000;
array[2926] <= 16'b0000_0000_0000_0000;
array[2927] <= 16'b0000_0000_0000_0000;
array[2928] <= 16'b0000_0000_0000_0000;
array[2929] <= 16'b0000_0000_0000_0000;
array[2930] <= 16'b0000_0000_0000_0000;
array[2931] <= 16'b0000_0000_0000_0000;
array[2932] <= 16'b0000_0000_0000_0000;
array[2933] <= 16'b0000_0000_0000_0000;
array[2934] <= 16'b0000_0000_0000_0000;
array[2935] <= 16'b0000_0000_0000_0000;
array[2936] <= 16'b0000_0000_0000_0000;
array[2937] <= 16'b0000_0000_0000_0000;
array[2938] <= 16'b0000_0000_0000_0000;
array[2939] <= 16'b0000_0000_0000_0000;
array[2940] <= 16'b0000_0000_0000_0000;
array[2941] <= 16'b0000_0000_0000_0000;
array[2942] <= 16'b0000_0000_0000_0000;
array[2943] <= 16'b0000_0000_0000_0000;
array[2944] <= 16'b0000_0000_0000_0000;
array[2945] <= 16'b0000_0000_0000_0000;
array[2946] <= 16'b0000_0000_0000_0000;
array[2947] <= 16'b0000_0000_0000_0000;
array[2948] <= 16'b0000_0000_0000_0000;
array[2949] <= 16'b0000_0000_0000_0000;
array[2950] <= 16'b0000_0000_0000_0000;
array[2951] <= 16'b0000_0000_0000_0000;
array[2952] <= 16'b0000_0000_0000_0000;
array[2953] <= 16'b0000_0000_0000_0000;
array[2954] <= 16'b0000_0000_0000_0000;
array[2955] <= 16'b0000_0000_0000_0000;
array[2956] <= 16'b0000_0000_0000_0000;
array[2957] <= 16'b0000_0000_0000_0000;
array[2958] <= 16'b0000_0000_0000_0000;
array[2959] <= 16'b0000_0000_0000_0000;
array[2960] <= 16'b0000_0000_0000_0000;
array[2961] <= 16'b0000_0000_0000_0000;
array[2962] <= 16'b0000_0000_0000_0000;
array[2963] <= 16'b0000_0000_0000_0000;
array[2964] <= 16'b0000_0000_0000_0000;
array[2965] <= 16'b0000_0000_0000_0000;
array[2966] <= 16'b0000_0000_0000_0000;
array[2967] <= 16'b0000_0000_0000_0000;
array[2968] <= 16'b0000_0000_0000_0000;
array[2969] <= 16'b0000_0000_0000_0000;
array[2970] <= 16'b0000_0000_0000_0000;
array[2971] <= 16'b0000_0000_0000_0000;
array[2972] <= 16'b0000_0000_0000_0000;
array[2973] <= 16'b0000_0000_0000_0000;
array[2974] <= 16'b0000_0000_0000_0000;
array[2975] <= 16'b0000_0000_0000_0000;
array[2976] <= 16'b0000_0000_0000_0000;
array[2977] <= 16'b0000_0000_0000_0000;
array[2978] <= 16'b0000_0000_0000_0000;
array[2979] <= 16'b0000_0000_0000_0000;
array[2980] <= 16'b0000_0000_0000_0000;
array[2981] <= 16'b0000_0000_0000_0000;
array[2982] <= 16'b0000_0000_0000_0000;
array[2983] <= 16'b0000_0000_0000_0000;
array[2984] <= 16'b0000_0000_0000_0000;
array[2985] <= 16'b0000_0000_0000_0000;
array[2986] <= 16'b0000_0000_0000_0000;
array[2987] <= 16'b0000_0000_0000_0000;
array[2988] <= 16'b0000_0000_0000_0000;
array[2989] <= 16'b0000_0000_0000_0000;
array[2990] <= 16'b0000_0000_0000_0000;
array[2991] <= 16'b0000_0000_0000_0000;
array[2992] <= 16'b0000_0000_0000_0000;
array[2993] <= 16'b0000_0000_0000_0000;
array[2994] <= 16'b0000_0000_0000_0000;
array[2995] <= 16'b0000_0000_0000_0000;
array[2996] <= 16'b0000_0000_0000_0000;
array[2997] <= 16'b0000_0000_0000_0000;
array[2998] <= 16'b0000_0000_0000_0000;
array[2999] <= 16'b0000_0000_0000_0000;
array[3000] <= 16'b0000_0000_0000_0000;
array[3001] <= 16'b0000_0000_0000_0000;
array[3002] <= 16'b0000_0000_0000_0000;
array[3003] <= 16'b0000_0000_0000_0000;
array[3004] <= 16'b0000_0000_0000_0000;
array[3005] <= 16'b0000_0000_0000_0000;
array[3006] <= 16'b0000_0000_0000_0000;
array[3007] <= 16'b0000_0000_0000_0000;
array[3008] <= 16'b0000_0000_0000_0000;
array[3009] <= 16'b0000_0000_0000_0000;
array[3010] <= 16'b0000_0000_0000_0000;
array[3011] <= 16'b0000_0000_0000_0000;
array[3012] <= 16'b0000_0000_0000_0000;
array[3013] <= 16'b0000_0000_0000_0000;
array[3014] <= 16'b0000_0000_0000_0000;
array[3015] <= 16'b0000_0000_0000_0000;
array[3016] <= 16'b0000_0000_0000_0000;
array[3017] <= 16'b0000_0000_0000_0000;
array[3018] <= 16'b0000_0000_0000_0000;
array[3019] <= 16'b0000_0000_0000_0000;
array[3020] <= 16'b0000_0000_0000_0000;
array[3021] <= 16'b0000_0000_0000_0000;
array[3022] <= 16'b0000_0000_0000_0000;
array[3023] <= 16'b0000_0000_0000_0000;
array[3024] <= 16'b0000_0000_0000_0000;
array[3025] <= 16'b0000_0000_0000_0000;
array[3026] <= 16'b0000_0000_0000_0000;
array[3027] <= 16'b0000_0000_0000_0000;
array[3028] <= 16'b0000_0000_0000_0000;
array[3029] <= 16'b0000_0000_0000_0000;
array[3030] <= 16'b0000_0000_0000_0000;
array[3031] <= 16'b0000_0000_0000_0000;
array[3032] <= 16'b0000_0000_0000_0000;
array[3033] <= 16'b0000_0000_0000_0000;
array[3034] <= 16'b0000_0000_0000_0000;
array[3035] <= 16'b0000_0000_0000_0000;
array[3036] <= 16'b0000_0000_0000_0000;
array[3037] <= 16'b0000_0000_0000_0000;
array[3038] <= 16'b0000_0000_0000_0000;
array[3039] <= 16'b0000_0000_0000_0000;
array[3040] <= 16'b0000_0000_0000_0000;
array[3041] <= 16'b0000_0000_0000_0000;
array[3042] <= 16'b0000_0000_0000_0000;
array[3043] <= 16'b0000_0000_0000_0000;
array[3044] <= 16'b0000_0000_0000_0000;
array[3045] <= 16'b0000_0000_0000_0000;
array[3046] <= 16'b0000_0000_0000_0000;
array[3047] <= 16'b0000_0000_0000_0000;
array[3048] <= 16'b0000_0000_0000_0000;
array[3049] <= 16'b0000_0000_0000_0000;
array[3050] <= 16'b0000_0000_0000_0000;
array[3051] <= 16'b0000_0000_0000_0000;
array[3052] <= 16'b0000_0000_0000_0000;
array[3053] <= 16'b0000_0000_0000_0000;
array[3054] <= 16'b0000_0000_0000_0000;
array[3055] <= 16'b0000_0000_0000_0000;
array[3056] <= 16'b0000_0000_0000_0000;
array[3057] <= 16'b0000_0000_0000_0000;
array[3058] <= 16'b0000_0000_0000_0000;
array[3059] <= 16'b0000_0000_0000_0000;
array[3060] <= 16'b0000_0000_0000_0000;
array[3061] <= 16'b0000_0000_0000_0000;
array[3062] <= 16'b0000_0000_0000_0000;
array[3063] <= 16'b0000_0000_0000_0000;
array[3064] <= 16'b0000_0000_0000_0000;
array[3065] <= 16'b0000_0000_0000_0000;
array[3066] <= 16'b0000_0000_0000_0000;
array[3067] <= 16'b0000_0000_0000_0000;
array[3068] <= 16'b0000_0000_0000_0000;
array[3069] <= 16'b0000_0000_0000_0000;
array[3070] <= 16'b0000_0000_0000_0000;
array[3071] <= 16'b0000_0000_0000_0000;
array[3072] <= 16'b0000_0000_0000_0000;
array[3073] <= 16'b0000_0000_0000_0000;
array[3074] <= 16'b0000_0000_0000_0000;
array[3075] <= 16'b0000_0000_0000_0000;
array[3076] <= 16'b0000_0000_0000_0000;
array[3077] <= 16'b0000_0000_0000_0000;
array[3078] <= 16'b0000_0000_0000_0000;
array[3079] <= 16'b0000_0000_0000_0000;
array[3080] <= 16'b0000_0000_0000_0000;
array[3081] <= 16'b0000_0000_0000_0000;
array[3082] <= 16'b0000_0000_0000_0000;
array[3083] <= 16'b0000_0000_0000_0000;
array[3084] <= 16'b0000_0000_0000_0000;
array[3085] <= 16'b0000_0000_0000_0000;
array[3086] <= 16'b0000_0000_0000_0000;
array[3087] <= 16'b0000_0000_0000_0000;
array[3088] <= 16'b0000_0000_0000_0000;
array[3089] <= 16'b0000_0000_0000_0000;
array[3090] <= 16'b0000_0000_0000_0000;
array[3091] <= 16'b0000_0000_0000_0000;
array[3092] <= 16'b0000_0000_0000_0000;
array[3093] <= 16'b0000_0000_0000_0000;
array[3094] <= 16'b0000_0000_0000_0000;
array[3095] <= 16'b0000_0000_0000_0000;
array[3096] <= 16'b0000_0000_0000_0000;
array[3097] <= 16'b0000_0000_0000_0000;
array[3098] <= 16'b0000_0000_0000_0000;
array[3099] <= 16'b0000_0000_0000_0000;
array[3100] <= 16'b0000_0000_0000_0000;
array[3101] <= 16'b0000_0000_0000_0000;
array[3102] <= 16'b0000_0000_0000_0000;
array[3103] <= 16'b0000_0000_0000_0000;
array[3104] <= 16'b0000_0000_0000_0000;
array[3105] <= 16'b0000_0000_0000_0000;
array[3106] <= 16'b0000_0000_0000_0000;
array[3107] <= 16'b0000_0000_0000_0000;
array[3108] <= 16'b0000_0000_0000_0000;
array[3109] <= 16'b0000_0000_0000_0000;
array[3110] <= 16'b0000_0000_0000_0000;
array[3111] <= 16'b0000_0000_0000_0000;
array[3112] <= 16'b0000_0000_0000_0000;
array[3113] <= 16'b0000_0000_0000_0000;
array[3114] <= 16'b0000_0000_0000_0000;
array[3115] <= 16'b0000_0000_0000_0000;
array[3116] <= 16'b0000_0000_0000_0000;
array[3117] <= 16'b0000_0000_0000_0000;
array[3118] <= 16'b0000_0000_0000_0000;
array[3119] <= 16'b0000_0000_0000_0000;
array[3120] <= 16'b0000_0000_0000_0000;
array[3121] <= 16'b0000_0000_0000_0000;
array[3122] <= 16'b0000_0000_0000_0000;
array[3123] <= 16'b0000_0000_0000_0000;
array[3124] <= 16'b0000_0000_0000_0000;
array[3125] <= 16'b0000_0000_0000_0000;
array[3126] <= 16'b0000_0000_0000_0000;
array[3127] <= 16'b0000_0000_0000_0000;
array[3128] <= 16'b0000_0000_0000_0000;
array[3129] <= 16'b0000_0000_0000_0000;
array[3130] <= 16'b0000_0000_0000_0000;
array[3131] <= 16'b0000_0000_0000_0000;
array[3132] <= 16'b0000_0000_0000_0000;
array[3133] <= 16'b0000_0000_0000_0000;
array[3134] <= 16'b0000_0000_0000_0000;
array[3135] <= 16'b0000_0000_0000_0000;
array[3136] <= 16'b0000_0000_0000_0000;
array[3137] <= 16'b0000_0000_0000_0000;
array[3138] <= 16'b0000_0000_0000_0000;
array[3139] <= 16'b0000_0000_0000_0000;
array[3140] <= 16'b0000_0000_0000_0000;
array[3141] <= 16'b0000_0000_0000_0000;
array[3142] <= 16'b0000_0000_0000_0000;
array[3143] <= 16'b0000_0000_0000_0000;
array[3144] <= 16'b0000_0000_0000_0000;
array[3145] <= 16'b0000_0000_0000_0000;
array[3146] <= 16'b0000_0000_0000_0000;
array[3147] <= 16'b0000_0000_0000_0000;
array[3148] <= 16'b0000_0000_0000_0000;
array[3149] <= 16'b0000_0000_0000_0000;
array[3150] <= 16'b0000_0000_0000_0000;
array[3151] <= 16'b0000_0000_0000_0000;
array[3152] <= 16'b0000_0000_0000_0000;
array[3153] <= 16'b0000_0000_0000_0000;
array[3154] <= 16'b0000_0000_0000_0000;
array[3155] <= 16'b0000_0000_0000_0000;
array[3156] <= 16'b0000_0000_0000_0000;
array[3157] <= 16'b0000_0000_0000_0000;
array[3158] <= 16'b0000_0000_0000_0000;
array[3159] <= 16'b0000_0000_0000_0000;
array[3160] <= 16'b0000_0000_0000_0000;
array[3161] <= 16'b0000_0000_0000_0000;
array[3162] <= 16'b0000_0000_0000_0000;
array[3163] <= 16'b0000_0000_0000_0000;
array[3164] <= 16'b0000_0000_0000_0000;
array[3165] <= 16'b0000_0000_0000_0000;
array[3166] <= 16'b0000_0000_0000_0000;
array[3167] <= 16'b0000_0000_0000_0000;
array[3168] <= 16'b0000_0000_0000_0000;
array[3169] <= 16'b0000_0000_0000_0000;
array[3170] <= 16'b0000_0000_0000_0000;
array[3171] <= 16'b0000_0000_0000_0000;
array[3172] <= 16'b0000_0000_0000_0000;
array[3173] <= 16'b0000_0000_0000_0000;
array[3174] <= 16'b0000_0000_0000_0000;
array[3175] <= 16'b0000_0000_0000_0000;
array[3176] <= 16'b0000_0000_0000_0000;
array[3177] <= 16'b0000_0000_0000_0000;
array[3178] <= 16'b0000_0000_0000_0000;
array[3179] <= 16'b0000_0000_0000_0000;
array[3180] <= 16'b0000_0000_0000_0000;
array[3181] <= 16'b0000_0000_0000_0000;
array[3182] <= 16'b0000_0000_0000_0000;
array[3183] <= 16'b0000_0000_0000_0000;
array[3184] <= 16'b0000_0000_0000_0000;
array[3185] <= 16'b0000_0000_0000_0000;
array[3186] <= 16'b0000_0000_0000_0000;
array[3187] <= 16'b0000_0000_0000_0000;
array[3188] <= 16'b0000_0000_0000_0000;
array[3189] <= 16'b0000_0000_0000_0000;
array[3190] <= 16'b0000_0000_0000_0000;
array[3191] <= 16'b0000_0000_0000_0000;
array[3192] <= 16'b0000_0000_0000_0000;
array[3193] <= 16'b0000_0000_0000_0000;
array[3194] <= 16'b0000_0000_0000_0000;
array[3195] <= 16'b0000_0000_0000_0000;
array[3196] <= 16'b0000_0000_0000_0000;
array[3197] <= 16'b0000_0000_0000_0000;
array[3198] <= 16'b0000_0000_0000_0000;
array[3199] <= 16'b0000_0000_0000_0000;
array[3200] <= 16'b0000_0000_0000_0000;
array[3201] <= 16'b0000_0000_0000_0000;
array[3202] <= 16'b0000_0000_0000_0000;
array[3203] <= 16'b0000_0000_0000_0000;
array[3204] <= 16'b0000_0000_0000_0000;
array[3205] <= 16'b0000_0000_0000_0000;
array[3206] <= 16'b0000_0000_0000_0000;
array[3207] <= 16'b0000_0000_0000_0000;
array[3208] <= 16'b0000_0000_0000_0000;
array[3209] <= 16'b0000_0000_0000_0000;
array[3210] <= 16'b0000_0000_0000_0000;
array[3211] <= 16'b0000_0000_0000_0000;
array[3212] <= 16'b0000_0000_0000_0000;
array[3213] <= 16'b0000_0000_0000_0000;
array[3214] <= 16'b0000_0000_0000_0000;
array[3215] <= 16'b0000_0000_0000_0000;
array[3216] <= 16'b0000_0000_0000_0000;
array[3217] <= 16'b0000_0000_0000_0000;
array[3218] <= 16'b0000_0000_0000_0000;
array[3219] <= 16'b0000_0000_0000_0000;
array[3220] <= 16'b0000_0000_0000_0000;
array[3221] <= 16'b0000_0000_0000_0000;
array[3222] <= 16'b0000_0000_0000_0000;
array[3223] <= 16'b0000_0000_0000_0000;
array[3224] <= 16'b0000_0000_0000_0000;
array[3225] <= 16'b0000_0000_0000_0000;
array[3226] <= 16'b0000_0000_0000_0000;
array[3227] <= 16'b0000_0000_0000_0000;
array[3228] <= 16'b0000_0000_0000_0000;
array[3229] <= 16'b0000_0000_0000_0000;
array[3230] <= 16'b0000_0000_0000_0000;
array[3231] <= 16'b0000_0000_0000_0000;
array[3232] <= 16'b0000_0000_0000_0000;
array[3233] <= 16'b0000_0000_0000_0000;
array[3234] <= 16'b0000_0000_0000_0000;
array[3235] <= 16'b0000_0000_0000_0000;
array[3236] <= 16'b0000_0000_0000_0000;
array[3237] <= 16'b0000_0000_0000_0000;
array[3238] <= 16'b0000_0000_0000_0000;
array[3239] <= 16'b0000_0000_0000_0000;
array[3240] <= 16'b0000_0000_0000_0000;
array[3241] <= 16'b0000_0000_0000_0000;
array[3242] <= 16'b0000_0000_0000_0000;
array[3243] <= 16'b0000_0000_0000_0000;
array[3244] <= 16'b0000_0000_0000_0000;
array[3245] <= 16'b0000_0000_0000_0000;
array[3246] <= 16'b0000_0000_0000_0000;
array[3247] <= 16'b0000_0000_0000_0000;
array[3248] <= 16'b0000_0000_0000_0000;
array[3249] <= 16'b0000_0000_0000_0000;
array[3250] <= 16'b0000_0000_0000_0000;
array[3251] <= 16'b0000_0000_0000_0000;
array[3252] <= 16'b0000_0000_0000_0000;
array[3253] <= 16'b0000_0000_0000_0000;
array[3254] <= 16'b0000_0000_0000_0000;
array[3255] <= 16'b0000_0000_0000_0000;
array[3256] <= 16'b0000_0000_0000_0000;
array[3257] <= 16'b0000_0000_0000_0000;
array[3258] <= 16'b0000_0000_0000_0000;
array[3259] <= 16'b0000_0000_0000_0000;
array[3260] <= 16'b0000_0000_0000_0000;
array[3261] <= 16'b0000_0000_0000_0000;
array[3262] <= 16'b0000_0000_0000_0000;
array[3263] <= 16'b0000_0000_0000_0000;
array[3264] <= 16'b0000_0000_0000_0000;
array[3265] <= 16'b0000_0000_0000_0000;
array[3266] <= 16'b0000_0000_0000_0000;
array[3267] <= 16'b0000_0000_0000_0000;
array[3268] <= 16'b0000_0000_0000_0000;
array[3269] <= 16'b0000_0000_0000_0000;
array[3270] <= 16'b0000_0000_0000_0000;
array[3271] <= 16'b0000_0000_0000_0000;
array[3272] <= 16'b0000_0000_0000_0000;
array[3273] <= 16'b0000_0000_0000_0000;
array[3274] <= 16'b0000_0000_0000_0000;
array[3275] <= 16'b0000_0000_0000_0000;
array[3276] <= 16'b0000_0000_0000_0000;
array[3277] <= 16'b0000_0000_0000_0000;
array[3278] <= 16'b0000_0000_0000_0000;
array[3279] <= 16'b0000_0000_0000_0000;
array[3280] <= 16'b0000_0000_0000_0000;
array[3281] <= 16'b0000_0000_0000_0000;
array[3282] <= 16'b0000_0000_0000_0000;
array[3283] <= 16'b0000_0000_0000_0000;
array[3284] <= 16'b0000_0000_0000_0000;
array[3285] <= 16'b0000_0000_0000_0000;
array[3286] <= 16'b0000_0000_0000_0000;
array[3287] <= 16'b0000_0000_0000_0000;
array[3288] <= 16'b0000_0000_0000_0000;
array[3289] <= 16'b0000_0000_0000_0000;
array[3290] <= 16'b0000_0000_0000_0000;
array[3291] <= 16'b0000_0000_0000_0000;
array[3292] <= 16'b0000_0000_0000_0000;
array[3293] <= 16'b0000_0000_0000_0000;
array[3294] <= 16'b0000_0000_0000_0000;
array[3295] <= 16'b0000_0000_0000_0000;
array[3296] <= 16'b0000_0000_0000_0000;
array[3297] <= 16'b0000_0000_0000_0000;
array[3298] <= 16'b0000_0000_0000_0000;
array[3299] <= 16'b0000_0000_0000_0000;
array[3300] <= 16'b0000_0000_0000_0000;
array[3301] <= 16'b0000_0000_0000_0000;
array[3302] <= 16'b0000_0000_0000_0000;
array[3303] <= 16'b0000_0000_0000_0000;
array[3304] <= 16'b0000_0000_0000_0000;
array[3305] <= 16'b0000_0000_0000_0000;
array[3306] <= 16'b0000_0000_0000_0000;
array[3307] <= 16'b0000_0000_0000_0000;
array[3308] <= 16'b0000_0000_0000_0000;
array[3309] <= 16'b0000_0000_0000_0000;
array[3310] <= 16'b0000_0000_0000_0000;
array[3311] <= 16'b0000_0000_0000_0000;
array[3312] <= 16'b0000_0000_0000_0000;
array[3313] <= 16'b0000_0000_0000_0000;
array[3314] <= 16'b0000_0000_0000_0000;
array[3315] <= 16'b0000_0000_0000_0000;
array[3316] <= 16'b0000_0000_0000_0000;
array[3317] <= 16'b0000_0000_0000_0000;
array[3318] <= 16'b0000_0000_0000_0000;
array[3319] <= 16'b0000_0000_0000_0000;
array[3320] <= 16'b0000_0000_0000_0000;
array[3321] <= 16'b0000_0000_0000_0000;
array[3322] <= 16'b0000_0000_0000_0000;
array[3323] <= 16'b0000_0000_0000_0000;
array[3324] <= 16'b0000_0000_0000_0000;
array[3325] <= 16'b0000_0000_0000_0000;
array[3326] <= 16'b0000_0000_0000_0000;
array[3327] <= 16'b0000_0000_0000_0000;
array[3328] <= 16'b0000_0000_0000_0000;
array[3329] <= 16'b0000_0000_0000_0000;
array[3330] <= 16'b0000_0000_0000_0000;
array[3331] <= 16'b0000_0000_0000_0000;
array[3332] <= 16'b0000_0000_0000_0000;
array[3333] <= 16'b0000_0000_0000_0000;
array[3334] <= 16'b0000_0000_0000_0000;
array[3335] <= 16'b0000_0000_0000_0000;
array[3336] <= 16'b0000_0000_0000_0000;
array[3337] <= 16'b0000_0000_0000_0000;
array[3338] <= 16'b0000_0000_0000_0000;
array[3339] <= 16'b0000_0000_0000_0000;
array[3340] <= 16'b0000_0000_0000_0000;
array[3341] <= 16'b0000_0000_0000_0000;
array[3342] <= 16'b0000_0000_0000_0000;
array[3343] <= 16'b0000_0000_0000_0000;
array[3344] <= 16'b0000_0000_0000_0000;
array[3345] <= 16'b0000_0000_0000_0000;
array[3346] <= 16'b0000_0000_0000_0000;
array[3347] <= 16'b0000_0000_0000_0000;
array[3348] <= 16'b0000_0000_0000_0000;
array[3349] <= 16'b0000_0000_0000_0000;
array[3350] <= 16'b0000_0000_0000_0000;
array[3351] <= 16'b0000_0000_0000_0000;
array[3352] <= 16'b0000_0000_0000_0000;
array[3353] <= 16'b0000_0000_0000_0000;
array[3354] <= 16'b0000_0000_0000_0000;
array[3355] <= 16'b0000_0000_0000_0000;
array[3356] <= 16'b0000_0000_0000_0000;
array[3357] <= 16'b0000_0000_0000_0000;
array[3358] <= 16'b0000_0000_0000_0000;
array[3359] <= 16'b0000_0000_0000_0000;
array[3360] <= 16'b0000_0000_0000_0000;
array[3361] <= 16'b0000_0000_0000_0000;
array[3362] <= 16'b0000_0000_0000_0000;
array[3363] <= 16'b0000_0000_0000_0000;
array[3364] <= 16'b0000_0000_0000_0000;
array[3365] <= 16'b0000_0000_0000_0000;
array[3366] <= 16'b0000_0000_0000_0000;
array[3367] <= 16'b0000_0000_0000_0000;
array[3368] <= 16'b0000_0000_0000_0000;
array[3369] <= 16'b0000_0000_0000_0000;
array[3370] <= 16'b0000_0000_0000_0000;
array[3371] <= 16'b0000_0000_0000_0000;
array[3372] <= 16'b0000_0000_0000_0000;
array[3373] <= 16'b0000_0000_0000_0000;
array[3374] <= 16'b0000_0000_0000_0000;
array[3375] <= 16'b0000_0000_0000_0000;
array[3376] <= 16'b0000_0000_0000_0000;
array[3377] <= 16'b0000_0000_0000_0000;
array[3378] <= 16'b0000_0000_0000_0000;
array[3379] <= 16'b0000_0000_0000_0000;
array[3380] <= 16'b0000_0000_0000_0000;
array[3381] <= 16'b0000_0000_0000_0000;
array[3382] <= 16'b0000_0000_0000_0000;
array[3383] <= 16'b0000_0000_0000_0000;
array[3384] <= 16'b0000_0000_0000_0000;
array[3385] <= 16'b0000_0000_0000_0000;
array[3386] <= 16'b0000_0000_0000_0000;
array[3387] <= 16'b0000_0000_0000_0000;
array[3388] <= 16'b0000_0000_0000_0000;
array[3389] <= 16'b0000_0000_0000_0000;
array[3390] <= 16'b0000_0000_0000_0000;
array[3391] <= 16'b0000_0000_0000_0000;
array[3392] <= 16'b0000_0000_0000_0000;
array[3393] <= 16'b0000_0000_0000_0000;
array[3394] <= 16'b0000_0000_0000_0000;
array[3395] <= 16'b0000_0000_0000_0000;
array[3396] <= 16'b0000_0000_0000_0000;
array[3397] <= 16'b0000_0000_0000_0000;
array[3398] <= 16'b0000_0000_0000_0000;
array[3399] <= 16'b0000_0000_0000_0000;
array[3400] <= 16'b0000_0000_0000_0000;
array[3401] <= 16'b0000_0000_0000_0000;
array[3402] <= 16'b0000_0000_0000_0000;
array[3403] <= 16'b0000_0000_0000_0000;
array[3404] <= 16'b0000_0000_0000_0000;
array[3405] <= 16'b0000_0000_0000_0000;
array[3406] <= 16'b0000_0000_0000_0000;
array[3407] <= 16'b0000_0000_0000_0000;
array[3408] <= 16'b0000_0000_0000_0000;
array[3409] <= 16'b0000_0000_0000_0000;
array[3410] <= 16'b0000_0000_0000_0000;
array[3411] <= 16'b0000_0000_0000_0000;
array[3412] <= 16'b0000_0000_0000_0000;
array[3413] <= 16'b0000_0000_0000_0000;
array[3414] <= 16'b0000_0000_0000_0000;
array[3415] <= 16'b0000_0000_0000_0000;
array[3416] <= 16'b0000_0000_0000_0000;
array[3417] <= 16'b0000_0000_0000_0000;
array[3418] <= 16'b0000_0000_0000_0000;
array[3419] <= 16'b0000_0000_0000_0000;
array[3420] <= 16'b0000_0000_0000_0000;
array[3421] <= 16'b0000_0000_0000_0000;
array[3422] <= 16'b0000_0000_0000_0000;
array[3423] <= 16'b0000_0000_0000_0000;
array[3424] <= 16'b0000_0000_0000_0000;
array[3425] <= 16'b0000_0000_0000_0000;
array[3426] <= 16'b0000_0000_0000_0000;
array[3427] <= 16'b0000_0000_0000_0000;
array[3428] <= 16'b0000_0000_0000_0000;
array[3429] <= 16'b0000_0000_0000_0000;
array[3430] <= 16'b0000_0000_0000_0000;
array[3431] <= 16'b0000_0000_0000_0000;
array[3432] <= 16'b0000_0000_0000_0000;
array[3433] <= 16'b0000_0000_0000_0000;
array[3434] <= 16'b0000_0000_0000_0000;
array[3435] <= 16'b0000_0000_0000_0000;
array[3436] <= 16'b0000_0000_0000_0000;
array[3437] <= 16'b0000_0000_0000_0000;
array[3438] <= 16'b0000_0000_0000_0000;
array[3439] <= 16'b0000_0000_0000_0000;
array[3440] <= 16'b0000_0000_0000_0000;
array[3441] <= 16'b0000_0000_0000_0000;
array[3442] <= 16'b0000_0000_0000_0000;
array[3443] <= 16'b0000_0000_0000_0000;
array[3444] <= 16'b0000_0000_0000_0000;
array[3445] <= 16'b0000_0000_0000_0000;
array[3446] <= 16'b0000_0000_0000_0000;
array[3447] <= 16'b0000_0000_0000_0000;
array[3448] <= 16'b0000_0000_0000_0000;
array[3449] <= 16'b0000_0000_0000_0000;
array[3450] <= 16'b0000_0000_0000_0000;
array[3451] <= 16'b0000_0000_0000_0000;
array[3452] <= 16'b0000_0000_0000_0000;
array[3453] <= 16'b0000_0000_0000_0000;
array[3454] <= 16'b0000_0000_0000_0000;
array[3455] <= 16'b0000_0000_0000_0000;
array[3456] <= 16'b0000_0000_0000_0000;
array[3457] <= 16'b0000_0000_0000_0000;
array[3458] <= 16'b0000_0000_0000_0000;
array[3459] <= 16'b0000_0000_0000_0000;
array[3460] <= 16'b0000_0000_0000_0000;
array[3461] <= 16'b0000_0000_0000_0000;
array[3462] <= 16'b0000_0000_0000_0000;
array[3463] <= 16'b0000_0000_0000_0000;
array[3464] <= 16'b0000_0000_0000_0000;
array[3465] <= 16'b0000_0000_0000_0000;
array[3466] <= 16'b0000_0000_0000_0000;
array[3467] <= 16'b0000_0000_0000_0000;
array[3468] <= 16'b0000_0000_0000_0000;
array[3469] <= 16'b0000_0000_0000_0000;
array[3470] <= 16'b0000_0000_0000_0000;
array[3471] <= 16'b0000_0000_0000_0000;
array[3472] <= 16'b0000_0000_0000_0000;
array[3473] <= 16'b0000_0000_0000_0000;
array[3474] <= 16'b0000_0000_0000_0000;
array[3475] <= 16'b0000_0000_0000_0000;
array[3476] <= 16'b0000_0000_0000_0000;
array[3477] <= 16'b0000_0000_0000_0000;
array[3478] <= 16'b0000_0000_0000_0000;
array[3479] <= 16'b0000_0000_0000_0000;
array[3480] <= 16'b0000_0000_0000_0000;
array[3481] <= 16'b0000_0000_0000_0000;
array[3482] <= 16'b0000_0000_0000_0000;
array[3483] <= 16'b0000_0000_0000_0000;
array[3484] <= 16'b0000_0000_0000_0000;
array[3485] <= 16'b0000_0000_0000_0000;
array[3486] <= 16'b0000_0000_0000_0000;
array[3487] <= 16'b0000_0000_0000_0000;
array[3488] <= 16'b0000_0000_0000_0000;
array[3489] <= 16'b0000_0000_0000_0000;
array[3490] <= 16'b0000_0000_0000_0000;
array[3491] <= 16'b0000_0000_0000_0000;
array[3492] <= 16'b0000_0000_0000_0000;
array[3493] <= 16'b0000_0000_0000_0000;
array[3494] <= 16'b0000_0000_0000_0000;
array[3495] <= 16'b0000_0000_0000_0000;
array[3496] <= 16'b0000_0000_0000_0000;
array[3497] <= 16'b0000_0000_0000_0000;
array[3498] <= 16'b0000_0000_0000_0000;
array[3499] <= 16'b0000_0000_0000_0000;
array[3500] <= 16'b0000_0000_0000_0000;
array[3501] <= 16'b0000_0000_0000_0000;
array[3502] <= 16'b0000_0000_0000_0000;
array[3503] <= 16'b0000_0000_0000_0000;
array[3504] <= 16'b0000_0000_0000_0000;
array[3505] <= 16'b0000_0000_0000_0000;
array[3506] <= 16'b0000_0000_0000_0000;
array[3507] <= 16'b0000_0000_0000_0000;
array[3508] <= 16'b0000_0000_0000_0000;
array[3509] <= 16'b0000_0000_0000_0000;
array[3510] <= 16'b0000_0000_0000_0000;
array[3511] <= 16'b0000_0000_0000_0000;
array[3512] <= 16'b0000_0000_0000_0000;
array[3513] <= 16'b0000_0000_0000_0000;
array[3514] <= 16'b0000_0000_0000_0000;
array[3515] <= 16'b0000_0000_0000_0000;
array[3516] <= 16'b0000_0000_0000_0000;
array[3517] <= 16'b0000_0000_0000_0000;
array[3518] <= 16'b0000_0000_0000_0000;
array[3519] <= 16'b0000_0000_0000_0000;
array[3520] <= 16'b0000_0000_0000_0000;
array[3521] <= 16'b0000_0000_0000_0000;
array[3522] <= 16'b0000_0000_0000_0000;
array[3523] <= 16'b0000_0000_0000_0000;
array[3524] <= 16'b0000_0000_0000_0000;
array[3525] <= 16'b0000_0000_0000_0000;
array[3526] <= 16'b0000_0000_0000_0000;
array[3527] <= 16'b0000_0000_0000_0000;
array[3528] <= 16'b0000_0000_0000_0000;
array[3529] <= 16'b0000_0000_0000_0000;
array[3530] <= 16'b0000_0000_0000_0000;
array[3531] <= 16'b0000_0000_0000_0000;
array[3532] <= 16'b0000_0000_0000_0000;
array[3533] <= 16'b0000_0000_0000_0000;
array[3534] <= 16'b0000_0000_0000_0000;
array[3535] <= 16'b0000_0000_0000_0000;
array[3536] <= 16'b0000_0000_0000_0000;
array[3537] <= 16'b0000_0000_0000_0000;
array[3538] <= 16'b0000_0000_0000_0000;
array[3539] <= 16'b0000_0000_0000_0000;
array[3540] <= 16'b0000_0000_0000_0000;
array[3541] <= 16'b0000_0000_0000_0000;
array[3542] <= 16'b0000_0000_0000_0000;
array[3543] <= 16'b0000_0000_0000_0000;
array[3544] <= 16'b0000_0000_0000_0000;
array[3545] <= 16'b0000_0000_0000_0000;
array[3546] <= 16'b0000_0000_0000_0000;
array[3547] <= 16'b0000_0000_0000_0000;
array[3548] <= 16'b0000_0000_0000_0000;
array[3549] <= 16'b0000_0000_0000_0000;
array[3550] <= 16'b0000_0000_0000_0000;
array[3551] <= 16'b0000_0000_0000_0000;
array[3552] <= 16'b0000_0000_0000_0000;
array[3553] <= 16'b0000_0000_0000_0000;
array[3554] <= 16'b0000_0000_0000_0000;
array[3555] <= 16'b0000_0000_0000_0000;
array[3556] <= 16'b0000_0000_0000_0000;
array[3557] <= 16'b0000_0000_0000_0000;
array[3558] <= 16'b0000_0000_0000_0000;
array[3559] <= 16'b0000_0000_0000_0000;
array[3560] <= 16'b0000_0000_0000_0000;
array[3561] <= 16'b0000_0000_0000_0000;
array[3562] <= 16'b0000_0000_0000_0000;
array[3563] <= 16'b0000_0000_0000_0000;
array[3564] <= 16'b0000_0000_0000_0000;
array[3565] <= 16'b0000_0000_0000_0000;
array[3566] <= 16'b0000_0000_0000_0000;
array[3567] <= 16'b0000_0000_0000_0000;
array[3568] <= 16'b0000_0000_0000_0000;
array[3569] <= 16'b0000_0000_0000_0000;
array[3570] <= 16'b0000_0000_0000_0000;
array[3571] <= 16'b0000_0000_0000_0000;
array[3572] <= 16'b0000_0000_0000_0000;
array[3573] <= 16'b0000_0000_0000_0000;
array[3574] <= 16'b0000_0000_0000_0000;
array[3575] <= 16'b0000_0000_0000_0000;
array[3576] <= 16'b0000_0000_0000_0000;
array[3577] <= 16'b0000_0000_0000_0000;
array[3578] <= 16'b0000_0000_0000_0000;
array[3579] <= 16'b0000_0000_0000_0000;
array[3580] <= 16'b0000_0000_0000_0000;
array[3581] <= 16'b0000_0000_0000_0000;
array[3582] <= 16'b0000_0000_0000_0000;
array[3583] <= 16'b0000_0000_0000_0000;
array[3584] <= 16'b0000_0000_0000_0000;
array[3585] <= 16'b0000_0000_0000_0000;
array[3586] <= 16'b0000_0000_0000_0000;
array[3587] <= 16'b0000_0000_0000_0000;
array[3588] <= 16'b0000_0000_0000_0000;
array[3589] <= 16'b0000_0000_0000_0000;
array[3590] <= 16'b0000_0000_0000_0000;
array[3591] <= 16'b0000_0000_0000_0000;
array[3592] <= 16'b0000_0000_0000_0000;
array[3593] <= 16'b0000_0000_0000_0000;
array[3594] <= 16'b0000_0000_0000_0000;
array[3595] <= 16'b0000_0000_0000_0000;
array[3596] <= 16'b0000_0000_0000_0000;
array[3597] <= 16'b0000_0000_0000_0000;
array[3598] <= 16'b0000_0000_0000_0000;
array[3599] <= 16'b0000_0000_0000_0000;
array[3600] <= 16'b0000_0000_0000_0000;
array[3601] <= 16'b0000_0000_0000_0000;
array[3602] <= 16'b0000_0000_0000_0000;
array[3603] <= 16'b0000_0000_0000_0000;
array[3604] <= 16'b0000_0000_0000_0000;
array[3605] <= 16'b0000_0000_0000_0000;
array[3606] <= 16'b0000_0000_0000_0000;
array[3607] <= 16'b0000_0000_0000_0000;
array[3608] <= 16'b0000_0000_0000_0000;
array[3609] <= 16'b0000_0000_0000_0000;
array[3610] <= 16'b0000_0000_0000_0000;
array[3611] <= 16'b0000_0000_0000_0000;
array[3612] <= 16'b0000_0000_0000_0000;
array[3613] <= 16'b0000_0000_0000_0000;
array[3614] <= 16'b0000_0000_0000_0000;
array[3615] <= 16'b0000_0000_0000_0000;
array[3616] <= 16'b0000_0000_0000_0000;
array[3617] <= 16'b0000_0000_0000_0000;
array[3618] <= 16'b0000_0000_0000_0000;
array[3619] <= 16'b0000_0000_0000_0000;
array[3620] <= 16'b0000_0000_0000_0000;
array[3621] <= 16'b0000_0000_0000_0000;
array[3622] <= 16'b0000_0000_0000_0000;
array[3623] <= 16'b0000_0000_0000_0000;
array[3624] <= 16'b0000_0000_0000_0000;
array[3625] <= 16'b0000_0000_0000_0000;
array[3626] <= 16'b0000_0000_0000_0000;
array[3627] <= 16'b0000_0000_0000_0000;
array[3628] <= 16'b0000_0000_0000_0000;
array[3629] <= 16'b0000_0000_0000_0000;
array[3630] <= 16'b0000_0000_0000_0000;
array[3631] <= 16'b0000_0000_0000_0000;
array[3632] <= 16'b0000_0000_0000_0000;
array[3633] <= 16'b0000_0000_0000_0000;
array[3634] <= 16'b0000_0000_0000_0000;
array[3635] <= 16'b0000_0000_0000_0000;
array[3636] <= 16'b0000_0000_0000_0000;
array[3637] <= 16'b0000_0000_0000_0000;
array[3638] <= 16'b0000_0000_0000_0000;
array[3639] <= 16'b0000_0000_0000_0000;
array[3640] <= 16'b0000_0000_0000_0000;
array[3641] <= 16'b0000_0000_0000_0000;
array[3642] <= 16'b0000_0000_0000_0000;
array[3643] <= 16'b0000_0000_0000_0000;
array[3644] <= 16'b0000_0000_0000_0000;
array[3645] <= 16'b0000_0000_0000_0000;
array[3646] <= 16'b0000_0000_0000_0000;
array[3647] <= 16'b0000_0000_0000_0000;
array[3648] <= 16'b0000_0000_0000_0000;
array[3649] <= 16'b0000_0000_0000_0000;
array[3650] <= 16'b0000_0000_0000_0000;
array[3651] <= 16'b0000_0000_0000_0000;
array[3652] <= 16'b0000_0000_0000_0000;
array[3653] <= 16'b0000_0000_0000_0000;
array[3654] <= 16'b0000_0000_0000_0000;
array[3655] <= 16'b0000_0000_0000_0000;
array[3656] <= 16'b0000_0000_0000_0000;
array[3657] <= 16'b0000_0000_0000_0000;
array[3658] <= 16'b0000_0000_0000_0000;
array[3659] <= 16'b0000_0000_0000_0000;
array[3660] <= 16'b0000_0000_0000_0000;
array[3661] <= 16'b0000_0000_0000_0000;
array[3662] <= 16'b0000_0000_0000_0000;
array[3663] <= 16'b0000_0000_0000_0000;
array[3664] <= 16'b0000_0000_0000_0000;
array[3665] <= 16'b0000_0000_0000_0000;
array[3666] <= 16'b0000_0000_0000_0000;
array[3667] <= 16'b0000_0000_0000_0000;
array[3668] <= 16'b0000_0000_0000_0000;
array[3669] <= 16'b0000_0000_0000_0000;
array[3670] <= 16'b0000_0000_0000_0000;
array[3671] <= 16'b0000_0000_0000_0000;
array[3672] <= 16'b0000_0000_0000_0000;
array[3673] <= 16'b0000_0000_0000_0000;
array[3674] <= 16'b0000_0000_0000_0000;
array[3675] <= 16'b0000_0000_0000_0000;
array[3676] <= 16'b0000_0000_0000_0000;
array[3677] <= 16'b0000_0000_0000_0000;
array[3678] <= 16'b0000_0000_0000_0000;
array[3679] <= 16'b0000_0000_0000_0000;
array[3680] <= 16'b0000_0000_0000_0000;
array[3681] <= 16'b0000_0000_0000_0000;
array[3682] <= 16'b0000_0000_0000_0000;
array[3683] <= 16'b0000_0000_0000_0000;
array[3684] <= 16'b0000_0000_0000_0000;
array[3685] <= 16'b0000_0000_0000_0000;
array[3686] <= 16'b0000_0000_0000_0000;
array[3687] <= 16'b0000_0000_0000_0000;
array[3688] <= 16'b0000_0000_0000_0000;
array[3689] <= 16'b0000_0000_0000_0000;
array[3690] <= 16'b0000_0000_0000_0000;
array[3691] <= 16'b0000_0000_0000_0000;
array[3692] <= 16'b0000_0000_0000_0000;
array[3693] <= 16'b0000_0000_0000_0000;
array[3694] <= 16'b0000_0000_0000_0000;
array[3695] <= 16'b0000_0000_0000_0000;
array[3696] <= 16'b0000_0000_0000_0000;
array[3697] <= 16'b0000_0000_0000_0000;
array[3698] <= 16'b0000_0000_0000_0000;
array[3699] <= 16'b0000_0000_0000_0000;
array[3700] <= 16'b0000_0000_0000_0000;
array[3701] <= 16'b0000_0000_0000_0000;
array[3702] <= 16'b0000_0000_0000_0000;
array[3703] <= 16'b0000_0000_0000_0000;
array[3704] <= 16'b0000_0000_0000_0000;
array[3705] <= 16'b0000_0000_0000_0000;
array[3706] <= 16'b0000_0000_0000_0000;
array[3707] <= 16'b0000_0000_0000_0000;
array[3708] <= 16'b0000_0000_0000_0000;
array[3709] <= 16'b0000_0000_0000_0000;
array[3710] <= 16'b0000_0000_0000_0000;
array[3711] <= 16'b0000_0000_0000_0000;
array[3712] <= 16'b0000_0000_0000_0000;
array[3713] <= 16'b0000_0000_0000_0000;
array[3714] <= 16'b0000_0000_0000_0000;
array[3715] <= 16'b0000_0000_0000_0000;
array[3716] <= 16'b0000_0000_0000_0000;
array[3717] <= 16'b0000_0000_0000_0000;
array[3718] <= 16'b0000_0000_0000_0000;
array[3719] <= 16'b0000_0000_0000_0000;
array[3720] <= 16'b0000_0000_0000_0000;
array[3721] <= 16'b0000_0000_0000_0000;
array[3722] <= 16'b0000_0000_0000_0000;
array[3723] <= 16'b0000_0000_0000_0000;
array[3724] <= 16'b0000_0000_0000_0000;
array[3725] <= 16'b0000_0000_0000_0000;
array[3726] <= 16'b0000_0000_0000_0000;
array[3727] <= 16'b0000_0000_0000_0000;
array[3728] <= 16'b0000_0000_0000_0000;
array[3729] <= 16'b0000_0000_0000_0000;
array[3730] <= 16'b0000_0000_0000_0000;
array[3731] <= 16'b0000_0000_0000_0000;
array[3732] <= 16'b0000_0000_0000_0000;
array[3733] <= 16'b0000_0000_0000_0000;
array[3734] <= 16'b0000_0000_0000_0000;
array[3735] <= 16'b0000_0000_0000_0000;
array[3736] <= 16'b0000_0000_0000_0000;
array[3737] <= 16'b0000_0000_0000_0000;
array[3738] <= 16'b0000_0000_0000_0000;
array[3739] <= 16'b0000_0000_0000_0000;
array[3740] <= 16'b0000_0000_0000_0000;
array[3741] <= 16'b0000_0000_0000_0000;
array[3742] <= 16'b0000_0000_0000_0000;
array[3743] <= 16'b0000_0000_0000_0000;
array[3744] <= 16'b0000_0000_0000_0000;
array[3745] <= 16'b0000_0000_0000_0000;
array[3746] <= 16'b0000_0000_0000_0000;
array[3747] <= 16'b0000_0000_0000_0000;
array[3748] <= 16'b0000_0000_0000_0000;
array[3749] <= 16'b0000_0000_0000_0000;
array[3750] <= 16'b0000_0000_0000_0000;
array[3751] <= 16'b0000_0000_0000_0000;
array[3752] <= 16'b0000_0000_0000_0000;
array[3753] <= 16'b0000_0000_0000_0000;
array[3754] <= 16'b0000_0000_0000_0000;
array[3755] <= 16'b0000_0000_0000_0000;
array[3756] <= 16'b0000_0000_0000_0000;
array[3757] <= 16'b0000_0000_0000_0000;
array[3758] <= 16'b0000_0000_0000_0000;
array[3759] <= 16'b0000_0000_0000_0000;
array[3760] <= 16'b0000_0000_0000_0000;
array[3761] <= 16'b0000_0000_0000_0000;
array[3762] <= 16'b0000_0000_0000_0000;
array[3763] <= 16'b0000_0000_0000_0000;
array[3764] <= 16'b0000_0000_0000_0000;
array[3765] <= 16'b0000_0000_0000_0000;
array[3766] <= 16'b0000_0000_0000_0000;
array[3767] <= 16'b0000_0000_0000_0000;
array[3768] <= 16'b0000_0000_0000_0000;
array[3769] <= 16'b0000_0000_0000_0000;
array[3770] <= 16'b0000_0000_0000_0000;
array[3771] <= 16'b0000_0000_0000_0000;
array[3772] <= 16'b0000_0000_0000_0000;
array[3773] <= 16'b0000_0000_0000_0000;
array[3774] <= 16'b0000_0000_0000_0000;
array[3775] <= 16'b0000_0000_0000_0000;
array[3776] <= 16'b0000_0000_0000_0000;
array[3777] <= 16'b0000_0000_0000_0000;
array[3778] <= 16'b0000_0000_0000_0000;
array[3779] <= 16'b0000_0000_0000_0000;
array[3780] <= 16'b0000_0000_0000_0000;
array[3781] <= 16'b0000_0000_0000_0000;
array[3782] <= 16'b0000_0000_0000_0000;
array[3783] <= 16'b0000_0000_0000_0000;
array[3784] <= 16'b0000_0000_0000_0000;
array[3785] <= 16'b0000_0000_0000_0000;
array[3786] <= 16'b0000_0000_0000_0000;
array[3787] <= 16'b0000_0000_0000_0000;
array[3788] <= 16'b0000_0000_0000_0000;
array[3789] <= 16'b0000_0000_0000_0000;
array[3790] <= 16'b0000_0000_0000_0000;
array[3791] <= 16'b0000_0000_0000_0000;
array[3792] <= 16'b0000_0000_0000_0000;
array[3793] <= 16'b0000_0000_0000_0000;
array[3794] <= 16'b0000_0000_0000_0000;
array[3795] <= 16'b0000_0000_0000_0000;
array[3796] <= 16'b0000_0000_0000_0000;
array[3797] <= 16'b0000_0000_0000_0000;
array[3798] <= 16'b0000_0000_0000_0000;
array[3799] <= 16'b0000_0000_0000_0000;
array[3800] <= 16'b0000_0000_0000_0000;
array[3801] <= 16'b0000_0000_0000_0000;
array[3802] <= 16'b0000_0000_0000_0000;
array[3803] <= 16'b0000_0000_0000_0000;
array[3804] <= 16'b0000_0000_0000_0000;
array[3805] <= 16'b0000_0000_0000_0000;
array[3806] <= 16'b0000_0000_0000_0000;
array[3807] <= 16'b0000_0000_0000_0000;
array[3808] <= 16'b0000_0000_0000_0000;
array[3809] <= 16'b0000_0000_0000_0000;
array[3810] <= 16'b0000_0000_0000_0000;
array[3811] <= 16'b0000_0000_0000_0000;
array[3812] <= 16'b0000_0000_0000_0000;
array[3813] <= 16'b0000_0000_0000_0000;
array[3814] <= 16'b0000_0000_0000_0000;
array[3815] <= 16'b0000_0000_0000_0000;
array[3816] <= 16'b0000_0000_0000_0000;
array[3817] <= 16'b0000_0000_0000_0000;
array[3818] <= 16'b0000_0000_0000_0000;
array[3819] <= 16'b0000_0000_0000_0000;
array[3820] <= 16'b0000_0000_0000_0000;
array[3821] <= 16'b0000_0000_0000_0000;
array[3822] <= 16'b0000_0000_0000_0000;
array[3823] <= 16'b0000_0000_0000_0000;
array[3824] <= 16'b0000_0000_0000_0000;
array[3825] <= 16'b0000_0000_0000_0000;
array[3826] <= 16'b0000_0000_0000_0000;
array[3827] <= 16'b0000_0000_0000_0000;
array[3828] <= 16'b0000_0000_0000_0000;
array[3829] <= 16'b0000_0000_0000_0000;
array[3830] <= 16'b0000_0000_0000_0000;
array[3831] <= 16'b0000_0000_0000_0000;
array[3832] <= 16'b0000_0000_0000_0000;
array[3833] <= 16'b0000_0000_0000_0000;
array[3834] <= 16'b0000_0000_0000_0000;
array[3835] <= 16'b0000_0000_0000_0000;
array[3836] <= 16'b0000_0000_0000_0000;
array[3837] <= 16'b0000_0000_0000_0000;
array[3838] <= 16'b0000_0000_0000_0000;
array[3839] <= 16'b0000_0000_0000_0000;
array[3840] <= 16'b0000_0000_0000_0000;
array[3841] <= 16'b0000_0000_0000_0000;
array[3842] <= 16'b0000_0000_0000_0000;
array[3843] <= 16'b0000_0000_0000_0000;
array[3844] <= 16'b0000_0000_0000_0000;
array[3845] <= 16'b0000_0000_0000_0000;
array[3846] <= 16'b0000_0000_0000_0000;
array[3847] <= 16'b0000_0000_0000_0000;
array[3848] <= 16'b0000_0000_0000_0000;
array[3849] <= 16'b0000_0000_0000_0000;
array[3850] <= 16'b0000_0000_0000_0000;
array[3851] <= 16'b0000_0000_0000_0000;
array[3852] <= 16'b0000_0000_0000_0000;
array[3853] <= 16'b0000_0000_0000_0000;
array[3854] <= 16'b0000_0000_0000_0000;
array[3855] <= 16'b0000_0000_0000_0000;
array[3856] <= 16'b0000_0000_0000_0000;
array[3857] <= 16'b0000_0000_0000_0000;
array[3858] <= 16'b0000_0000_0000_0000;
array[3859] <= 16'b0000_0000_0000_0000;
array[3860] <= 16'b0000_0000_0000_0000;
array[3861] <= 16'b0000_0000_0000_0000;
array[3862] <= 16'b0000_0000_0000_0000;
array[3863] <= 16'b0000_0000_0000_0000;
array[3864] <= 16'b0000_0000_0000_0000;
array[3865] <= 16'b0000_0000_0000_0000;
array[3866] <= 16'b0000_0000_0000_0000;
array[3867] <= 16'b0000_0000_0000_0000;
array[3868] <= 16'b0000_0000_0000_0000;
array[3869] <= 16'b0000_0000_0000_0000;
array[3870] <= 16'b0000_0000_0000_0000;
array[3871] <= 16'b0000_0000_0000_0000;
array[3872] <= 16'b0000_0000_0000_0000;
array[3873] <= 16'b0000_0000_0000_0000;
array[3874] <= 16'b0000_0000_0000_0000;
array[3875] <= 16'b0000_0000_0000_0000;
array[3876] <= 16'b0000_0000_0000_0000;
array[3877] <= 16'b0000_0000_0000_0000;
array[3878] <= 16'b0000_0000_0000_0000;
array[3879] <= 16'b0000_0000_0000_0000;
array[3880] <= 16'b0000_0000_0000_0000;
array[3881] <= 16'b0000_0000_0000_0000;
array[3882] <= 16'b0000_0000_0000_0000;
array[3883] <= 16'b0000_0000_0000_0000;
array[3884] <= 16'b0000_0000_0000_0000;
array[3885] <= 16'b0000_0000_0000_0000;
array[3886] <= 16'b0000_0000_0000_0000;
array[3887] <= 16'b0000_0000_0000_0000;
array[3888] <= 16'b0000_0000_0000_0000;
array[3889] <= 16'b0000_0000_0000_0000;
array[3890] <= 16'b0000_0000_0000_0000;
array[3891] <= 16'b0000_0000_0000_0000;
array[3892] <= 16'b0000_0000_0000_0000;
array[3893] <= 16'b0000_0000_0000_0000;
array[3894] <= 16'b0000_0000_0000_0000;
array[3895] <= 16'b0000_0000_0000_0000;
array[3896] <= 16'b0000_0000_0000_0000;
array[3897] <= 16'b0000_0000_0000_0000;
array[3898] <= 16'b0000_0000_0000_0000;
array[3899] <= 16'b0000_0000_0000_0000;
array[3900] <= 16'b0000_0000_0000_0000;
array[3901] <= 16'b0000_0000_0000_0000;
array[3902] <= 16'b0000_0000_0000_0000;
array[3903] <= 16'b0000_0000_0000_0000;
array[3904] <= 16'b0000_0000_0000_0000;
array[3905] <= 16'b0000_0000_0000_0000;
array[3906] <= 16'b0000_0000_0000_0000;
array[3907] <= 16'b0000_0000_0000_0000;
array[3908] <= 16'b0000_0000_0000_0000;
array[3909] <= 16'b0000_0000_0000_0000;
array[3910] <= 16'b0000_0000_0000_0000;
array[3911] <= 16'b0000_0000_0000_0000;
array[3912] <= 16'b0000_0000_0000_0000;
array[3913] <= 16'b0000_0000_0000_0000;
array[3914] <= 16'b0000_0000_0000_0000;
array[3915] <= 16'b0000_0000_0000_0000;
array[3916] <= 16'b0000_0000_0000_0000;
array[3917] <= 16'b0000_0000_0000_0000;
array[3918] <= 16'b0000_0000_0000_0000;
array[3919] <= 16'b0000_0000_0000_0000;
array[3920] <= 16'b0000_0000_0000_0000;
array[3921] <= 16'b0000_0000_0000_0000;
array[3922] <= 16'b0000_0000_0000_0000;
array[3923] <= 16'b0000_0000_0000_0000;
array[3924] <= 16'b0000_0000_0000_0000;
array[3925] <= 16'b0000_0000_0000_0000;
array[3926] <= 16'b0000_0000_0000_0000;
array[3927] <= 16'b0000_0000_0000_0000;
array[3928] <= 16'b0000_0000_0000_0000;
array[3929] <= 16'b0000_0000_0000_0000;
array[3930] <= 16'b0000_0000_0000_0000;
array[3931] <= 16'b0000_0000_0000_0000;
array[3932] <= 16'b0000_0000_0000_0000;
array[3933] <= 16'b0000_0000_0000_0000;
array[3934] <= 16'b0000_0000_0000_0000;
array[3935] <= 16'b0000_0000_0000_0000;
array[3936] <= 16'b0000_0000_0000_0000;
array[3937] <= 16'b0000_0000_0000_0000;
array[3938] <= 16'b0000_0000_0000_0000;
array[3939] <= 16'b0000_0000_0000_0000;
array[3940] <= 16'b0000_0000_0000_0000;
array[3941] <= 16'b0000_0000_0000_0000;
array[3942] <= 16'b0000_0000_0000_0000;
array[3943] <= 16'b0000_0000_0000_0000;
array[3944] <= 16'b0000_0000_0000_0000;
array[3945] <= 16'b0000_0000_0000_0000;
array[3946] <= 16'b0000_0000_0000_0000;
array[3947] <= 16'b0000_0000_0000_0000;
array[3948] <= 16'b0000_0000_0000_0000;
array[3949] <= 16'b0000_0000_0000_0000;
array[3950] <= 16'b0000_0000_0000_0000;
array[3951] <= 16'b0000_0000_0000_0000;
array[3952] <= 16'b0000_0000_0000_0000;
array[3953] <= 16'b0000_0000_0000_0000;
array[3954] <= 16'b0000_0000_0000_0000;
array[3955] <= 16'b0000_0000_0000_0000;
array[3956] <= 16'b0000_0000_0000_0000;
array[3957] <= 16'b0000_0000_0000_0000;
array[3958] <= 16'b0000_0000_0000_0000;
array[3959] <= 16'b0000_0000_0000_0000;
array[3960] <= 16'b0000_0000_0000_0000;
array[3961] <= 16'b0000_0000_0000_0000;
array[3962] <= 16'b0000_0000_0000_0000;
array[3963] <= 16'b0000_0000_0000_0000;
array[3964] <= 16'b0000_0000_0000_0000;
array[3965] <= 16'b0000_0000_0000_0000;
array[3966] <= 16'b0000_0000_0000_0000;
array[3967] <= 16'b0000_0000_0000_0000;
array[3968] <= 16'b0000_0000_0000_0000;
array[3969] <= 16'b0000_0000_0000_0000;
array[3970] <= 16'b0000_0000_0000_0000;
array[3971] <= 16'b0000_0000_0000_0000;
array[3972] <= 16'b0000_0000_0000_0000;
array[3973] <= 16'b0000_0000_0000_0000;
array[3974] <= 16'b0000_0000_0000_0000;
array[3975] <= 16'b0000_0000_0000_0000;
array[3976] <= 16'b0000_0000_0000_0000;
array[3977] <= 16'b0000_0000_0000_0000;
array[3978] <= 16'b0000_0000_0000_0000;
array[3979] <= 16'b0000_0000_0000_0000;
array[3980] <= 16'b0000_0000_0000_0000;
array[3981] <= 16'b0000_0000_0000_0000;
array[3982] <= 16'b0000_0000_0000_0000;
array[3983] <= 16'b0000_0000_0000_0000;
array[3984] <= 16'b0000_0000_0000_0000;
array[3985] <= 16'b0000_0000_0000_0000;
array[3986] <= 16'b0000_0000_0000_0000;
array[3987] <= 16'b0000_0000_0000_0000;
array[3988] <= 16'b0000_0000_0000_0000;
array[3989] <= 16'b0000_0000_0000_0000;
array[3990] <= 16'b0000_0000_0000_0000;
array[3991] <= 16'b0000_0000_0000_0000;
array[3992] <= 16'b0000_0000_0000_0000;
array[3993] <= 16'b0000_0000_0000_0000;
array[3994] <= 16'b0000_0000_0000_0000;
array[3995] <= 16'b0000_0000_0000_0000;
array[3996] <= 16'b0000_0000_0000_0000;
array[3997] <= 16'b0000_0000_0000_0000;
array[3998] <= 16'b0000_0000_0000_0000;
array[3999] <= 16'b0000_0000_0000_0000;
array[4000] <= 16'b0000_0000_0000_0000;
array[4001] <= 16'b0000_0000_0000_0000;
array[4002] <= 16'b0000_0000_0000_0000;
array[4003] <= 16'b0000_0000_0000_0000;
array[4004] <= 16'b0000_0000_0000_0000;
array[4005] <= 16'b0000_0000_0000_0000;
array[4006] <= 16'b0000_0000_0000_0000;
array[4007] <= 16'b0000_0000_0000_0000;
array[4008] <= 16'b0000_0000_0000_0000;
array[4009] <= 16'b0000_0000_0000_0000;
array[4010] <= 16'b0000_0000_0000_0000;
array[4011] <= 16'b0000_0000_0000_0000;
array[4012] <= 16'b0000_0000_0000_0000;
array[4013] <= 16'b0000_0000_0000_0000;
array[4014] <= 16'b0000_0000_0000_0000;
array[4015] <= 16'b0000_0000_0000_0000;
array[4016] <= 16'b0000_0000_0000_0000;
array[4017] <= 16'b0000_0000_0000_0000;
array[4018] <= 16'b0000_0000_0000_0000;
array[4019] <= 16'b0000_0000_0000_0000;
array[4020] <= 16'b0000_0000_0000_0000;
array[4021] <= 16'b0000_0000_0000_0000;
array[4022] <= 16'b0000_0000_0000_0000;
array[4023] <= 16'b0000_0000_0000_0000;
array[4024] <= 16'b0000_0000_0000_0000;
array[4025] <= 16'b0000_0000_0000_0000;
array[4026] <= 16'b0000_0000_0000_0000;
array[4027] <= 16'b0000_0000_0000_0000;
array[4028] <= 16'b0000_0000_0000_0000;
array[4029] <= 16'b0000_0000_0000_0000;
array[4030] <= 16'b0000_0000_0000_0000;
array[4031] <= 16'b0000_0000_0000_0000;
array[4032] <= 16'b0000_0000_0000_0000;
array[4033] <= 16'b0000_0000_0000_0000;
array[4034] <= 16'b0000_0000_0000_0000;
array[4035] <= 16'b0000_0000_0000_0000;
array[4036] <= 16'b0000_0000_0000_0000;
array[4037] <= 16'b0000_0000_0000_0000;
array[4038] <= 16'b0000_0000_0000_0000;
array[4039] <= 16'b0000_0000_0000_0000;
array[4040] <= 16'b0000_0000_0000_0000;
array[4041] <= 16'b0000_0000_0000_0000;
array[4042] <= 16'b0000_0000_0000_0000;
array[4043] <= 16'b0000_0000_0000_0000;
array[4044] <= 16'b0000_0000_0000_0000;
array[4045] <= 16'b0000_0000_0000_0000;
array[4046] <= 16'b0000_0000_0000_0000;
array[4047] <= 16'b0000_0000_0000_0000;
array[4048] <= 16'b0000_0000_0000_0000;
array[4049] <= 16'b0000_0000_0000_0000;
array[4050] <= 16'b0000_0000_0000_0000;
array[4051] <= 16'b0000_0000_0000_0000;
array[4052] <= 16'b0000_0000_0000_0000;
array[4053] <= 16'b0000_0000_0000_0000;
array[4054] <= 16'b0000_0000_0000_0000;
array[4055] <= 16'b0000_0000_0000_0000;
array[4056] <= 16'b0000_0000_0000_0000;
array[4057] <= 16'b0000_0000_0000_0000;
array[4058] <= 16'b0000_0000_0000_0000;
array[4059] <= 16'b0000_0000_0000_0000;
array[4060] <= 16'b0000_0000_0000_0000;
array[4061] <= 16'b0000_0000_0000_0000;
array[4062] <= 16'b0000_0000_0000_0000;
array[4063] <= 16'b0000_0000_0000_0000;
array[4064] <= 16'b0000_0000_0000_0000;
array[4065] <= 16'b0000_0000_0000_0000;
array[4066] <= 16'b0000_0000_0000_0000;
array[4067] <= 16'b0000_0000_0000_0000;
array[4068] <= 16'b0000_0000_0000_0000;
array[4069] <= 16'b0000_0000_0000_0000;
array[4070] <= 16'b0000_0000_0000_0000;
array[4071] <= 16'b0000_0000_0000_0000;
array[4072] <= 16'b0000_0000_0000_0000;
array[4073] <= 16'b0000_0000_0000_0000;
array[4074] <= 16'b0000_0000_0000_0000;
array[4075] <= 16'b0000_0000_0000_0000;
array[4076] <= 16'b0000_0000_0000_0000;
array[4077] <= 16'b0000_0000_0000_0000;
array[4078] <= 16'b0000_0000_0000_0000;
array[4079] <= 16'b0000_0000_0000_0000;
array[4080] <= 16'b0000_0000_0000_0000;
array[4081] <= 16'b0000_0000_0000_0000;
array[4082] <= 16'b0000_0000_0000_0000;
array[4083] <= 16'b0000_0000_0000_0000;
array[4084] <= 16'b0000_0000_0000_0000;
array[4085] <= 16'b0000_0000_0000_0000;
array[4086] <= 16'b0000_0000_0000_0000;
array[4087] <= 16'b0000_0000_0000_0000;
array[4088] <= 16'b0000_0000_0000_0000;
array[4089] <= 16'b0000_0000_0000_0000;
array[4090] <= 16'b0000_0000_0000_0000;
array[4091] <= 16'b0000_0000_0000_0000;
array[4092] <= 16'b0000_0000_0000_0000;
array[4093] <= 16'b0000_0000_0000_0000;
array[4094] <= 16'b0000_0000_0000_0000;
array[4095] <= 16'b0000_0000_0000_0000;
array[4096] <= 16'b0000_0000_0000_0000;
array[4097] <= 16'b0000_0000_0000_0000;
array[4098] <= 16'b0000_0000_0000_0000;
array[4099] <= 16'b0000_0000_0000_0000;
array[4100] <= 16'b0000_0000_0000_0000;
array[4101] <= 16'b0000_0000_0000_0000;
array[4102] <= 16'b0000_0000_0000_0000;
array[4103] <= 16'b0000_0000_0000_0000;
array[4104] <= 16'b0000_0000_0000_0000;
array[4105] <= 16'b0000_0000_0000_0000;
array[4106] <= 16'b0000_0000_0000_0000;
array[4107] <= 16'b0000_0000_0000_0000;
array[4108] <= 16'b0000_0000_0000_0000;
array[4109] <= 16'b0000_0000_0000_0000;
array[4110] <= 16'b0000_0000_0000_0000;
array[4111] <= 16'b0000_0000_0000_0000;
array[4112] <= 16'b0000_0000_0000_0000;
array[4113] <= 16'b0000_0000_0000_0000;
array[4114] <= 16'b0000_0000_0000_0000;
array[4115] <= 16'b0000_0000_0000_0000;
array[4116] <= 16'b0000_0000_0000_0000;
array[4117] <= 16'b0000_0000_0000_0000;
array[4118] <= 16'b0000_0000_0000_0000;
array[4119] <= 16'b0000_0000_0000_0000;
array[4120] <= 16'b0000_0000_0000_0000;
array[4121] <= 16'b0000_0000_0000_0000;
array[4122] <= 16'b0000_0000_0000_0000;
array[4123] <= 16'b0000_0000_0000_0000;
array[4124] <= 16'b0000_0000_0000_0000;
array[4125] <= 16'b0000_0000_0000_0000;
array[4126] <= 16'b0000_0000_0000_0000;
array[4127] <= 16'b0000_0000_0000_0000;
array[4128] <= 16'b0000_0000_0000_0000;
array[4129] <= 16'b0000_0000_0000_0000;
array[4130] <= 16'b0000_0000_0000_0000;
array[4131] <= 16'b0000_0000_0000_0000;
array[4132] <= 16'b0000_0000_0000_0000;
array[4133] <= 16'b0000_0000_0000_0000;
array[4134] <= 16'b0000_0000_0000_0000;
array[4135] <= 16'b0000_0000_0000_0000;
array[4136] <= 16'b0000_0000_0000_0000;
array[4137] <= 16'b0000_0000_0000_0000;
array[4138] <= 16'b0000_0000_0000_0000;
array[4139] <= 16'b0000_0000_0000_0000;
array[4140] <= 16'b0000_0000_0000_0000;
array[4141] <= 16'b0000_0000_0000_0000;
array[4142] <= 16'b0000_0000_0000_0000;
array[4143] <= 16'b0000_0000_0000_0000;
array[4144] <= 16'b0000_0000_0000_0000;
array[4145] <= 16'b0000_0000_0000_0000;
array[4146] <= 16'b0000_0000_0000_0000;
array[4147] <= 16'b0000_0000_0000_0000;
array[4148] <= 16'b0000_0000_0000_0000;
array[4149] <= 16'b0000_0000_0000_0000;
array[4150] <= 16'b0000_0000_0000_0000;
array[4151] <= 16'b0000_0000_0000_0000;
array[4152] <= 16'b0000_0000_0000_0000;
array[4153] <= 16'b0000_0000_0000_0000;
array[4154] <= 16'b0000_0000_0000_0000;
array[4155] <= 16'b0000_0000_0000_0000;
array[4156] <= 16'b0000_0000_0000_0000;
array[4157] <= 16'b0000_0000_0000_0000;
array[4158] <= 16'b0000_0000_0000_0000;
array[4159] <= 16'b0000_0000_0000_0000;
array[4160] <= 16'b0000_0000_0000_0000;
array[4161] <= 16'b0000_0000_0000_0000;
array[4162] <= 16'b0000_0000_0000_0000;
array[4163] <= 16'b0000_0000_0000_0000;
array[4164] <= 16'b0000_0000_0000_0000;
array[4165] <= 16'b0000_0000_0000_0000;
array[4166] <= 16'b0000_0000_0000_0000;
array[4167] <= 16'b0000_0000_0000_0000;
array[4168] <= 16'b0000_0000_0000_0000;
array[4169] <= 16'b0000_0000_0000_0000;
array[4170] <= 16'b0000_0000_0000_0000;
array[4171] <= 16'b0000_0000_0000_0000;
array[4172] <= 16'b0000_0000_0000_0000;
array[4173] <= 16'b0000_0000_0000_0000;
array[4174] <= 16'b0000_0000_0000_0000;
array[4175] <= 16'b0000_0000_0000_0000;
array[4176] <= 16'b0000_0000_0000_0000;
array[4177] <= 16'b0000_0000_0000_0000;
array[4178] <= 16'b0000_0000_0000_0000;
array[4179] <= 16'b0000_0000_0000_0000;
array[4180] <= 16'b0000_0000_0000_0000;
array[4181] <= 16'b0000_0000_0000_0000;
array[4182] <= 16'b0000_0000_0000_0000;
array[4183] <= 16'b0000_0000_0000_0000;
array[4184] <= 16'b0000_0000_0000_0000;
array[4185] <= 16'b0000_0000_0000_0000;
array[4186] <= 16'b0000_0000_0000_0000;
array[4187] <= 16'b0000_0000_0000_0000;
array[4188] <= 16'b0000_0000_0000_0000;
array[4189] <= 16'b0000_0000_0000_0000;
array[4190] <= 16'b0000_0000_0000_0000;
array[4191] <= 16'b0000_0000_0000_0000;
array[4192] <= 16'b0000_0000_0000_0000;
array[4193] <= 16'b0000_0000_0000_0000;
array[4194] <= 16'b0000_0000_0000_0000;
array[4195] <= 16'b0000_0000_0000_0000;
array[4196] <= 16'b0000_0000_0000_0000;
array[4197] <= 16'b0000_0000_0000_0000;
array[4198] <= 16'b0000_0000_0000_0000;
array[4199] <= 16'b0000_0000_0000_0000;
array[4200] <= 16'b0000_0000_0000_0000;
array[4201] <= 16'b0000_0000_0000_0000;
array[4202] <= 16'b0000_0000_0000_0000;
array[4203] <= 16'b0000_0000_0000_0000;
array[4204] <= 16'b0000_0000_0000_0000;
array[4205] <= 16'b0000_0000_0000_0000;
array[4206] <= 16'b0000_0000_0000_0000;
array[4207] <= 16'b0000_0000_0000_0000;
array[4208] <= 16'b0000_0000_0000_0000;
array[4209] <= 16'b0000_0000_0000_0000;
array[4210] <= 16'b0000_0000_0000_0000;
array[4211] <= 16'b0000_0000_0000_0000;
array[4212] <= 16'b0000_0000_0000_0000;
array[4213] <= 16'b0000_0000_0000_0000;
array[4214] <= 16'b0000_0000_0000_0000;
array[4215] <= 16'b0000_0000_0000_0000;
array[4216] <= 16'b0000_0000_0000_0000;
array[4217] <= 16'b0000_0000_0000_0000;
array[4218] <= 16'b0000_0000_0000_0000;
array[4219] <= 16'b0000_0000_0000_0000;
array[4220] <= 16'b0000_0000_0000_0000;
array[4221] <= 16'b0000_0000_0000_0000;
array[4222] <= 16'b0000_0000_0000_0000;
array[4223] <= 16'b0000_0000_0000_0000;
array[4224] <= 16'b0000_0000_0000_0000;
array[4225] <= 16'b0000_0000_0000_0000;
array[4226] <= 16'b0000_0000_0000_0000;
array[4227] <= 16'b0000_0000_0000_0000;
array[4228] <= 16'b0000_0000_0000_0000;
array[4229] <= 16'b0000_0000_0000_0000;
array[4230] <= 16'b0000_0000_0000_0000;
array[4231] <= 16'b0000_0000_0000_0000;
array[4232] <= 16'b0000_0000_0000_0000;
array[4233] <= 16'b0000_0000_0000_0000;
array[4234] <= 16'b0000_0000_0000_0000;
array[4235] <= 16'b0000_0000_0000_0000;
array[4236] <= 16'b0000_0000_0000_0000;
array[4237] <= 16'b0000_0000_0000_0000;
array[4238] <= 16'b0000_0000_0000_0000;
array[4239] <= 16'b0000_0000_0000_0000;
array[4240] <= 16'b0000_0000_0000_0000;
array[4241] <= 16'b0000_0000_0000_0000;
array[4242] <= 16'b0000_0000_0000_0000;
array[4243] <= 16'b0000_0000_0000_0000;
array[4244] <= 16'b0000_0000_0000_0000;
array[4245] <= 16'b0000_0000_0000_0000;
array[4246] <= 16'b0000_0000_0000_0000;
array[4247] <= 16'b0000_0000_0000_0000;
array[4248] <= 16'b0000_0000_0000_0000;
array[4249] <= 16'b0000_0000_0000_0000;
array[4250] <= 16'b0000_0000_0000_0000;
array[4251] <= 16'b0000_0000_0000_0000;
array[4252] <= 16'b0000_0000_0000_0000;
array[4253] <= 16'b0000_0000_0000_0000;
array[4254] <= 16'b0000_0000_0000_0000;
array[4255] <= 16'b0000_0000_0000_0000;
array[4256] <= 16'b0000_0000_0000_0000;
array[4257] <= 16'b0000_0000_0000_0000;
array[4258] <= 16'b0000_0000_0000_0000;
array[4259] <= 16'b0000_0000_0000_0000;
array[4260] <= 16'b0000_0000_0000_0000;
array[4261] <= 16'b0000_0000_0000_0000;
array[4262] <= 16'b0000_0000_0000_0000;
array[4263] <= 16'b0000_0000_0000_0000;
array[4264] <= 16'b0000_0000_0000_0000;
array[4265] <= 16'b0000_0000_0000_0000;
array[4266] <= 16'b0000_0000_0000_0000;
array[4267] <= 16'b0000_0000_0000_0000;
array[4268] <= 16'b0000_0000_0000_0000;
array[4269] <= 16'b0000_0000_0000_0000;
array[4270] <= 16'b0000_0000_0000_0000;
array[4271] <= 16'b0000_0000_0000_0000;
array[4272] <= 16'b0000_0000_0000_0000;
array[4273] <= 16'b0000_0000_0000_0000;
array[4274] <= 16'b0000_0000_0000_0000;
array[4275] <= 16'b0000_0000_0000_0000;
array[4276] <= 16'b0000_0000_0000_0000;
array[4277] <= 16'b0000_0000_0000_0000;
array[4278] <= 16'b0000_0000_0000_0000;
array[4279] <= 16'b0000_0000_0000_0000;
array[4280] <= 16'b0000_0000_0000_0000;
array[4281] <= 16'b0000_0000_0000_0000;
array[4282] <= 16'b0000_0000_0000_0000;
array[4283] <= 16'b0000_0000_0000_0000;
array[4284] <= 16'b0000_0000_0000_0000;
array[4285] <= 16'b0000_0000_0000_0000;
array[4286] <= 16'b0000_0000_0000_0000;
array[4287] <= 16'b0000_0000_0000_0000;
array[4288] <= 16'b0000_0000_0000_0000;
array[4289] <= 16'b0000_0000_0000_0000;
array[4290] <= 16'b0000_0000_0000_0000;
array[4291] <= 16'b0000_0000_0000_0000;
array[4292] <= 16'b0000_0000_0000_0000;
array[4293] <= 16'b0000_0000_0000_0000;
array[4294] <= 16'b0000_0000_0000_0000;
array[4295] <= 16'b0000_0000_0000_0000;
array[4296] <= 16'b0000_0000_0000_0000;
array[4297] <= 16'b0000_0000_0000_0000;
array[4298] <= 16'b0000_0000_0000_0000;
array[4299] <= 16'b0000_0000_0000_0000;
array[4300] <= 16'b0000_0000_0000_0000;
array[4301] <= 16'b0000_0000_0000_0000;
array[4302] <= 16'b0000_0000_0000_0000;
array[4303] <= 16'b0000_0000_0000_0000;
array[4304] <= 16'b0000_0000_0000_0000;
array[4305] <= 16'b0000_0000_0000_0000;
array[4306] <= 16'b0000_0000_0000_0000;
array[4307] <= 16'b0000_0000_0000_0000;
array[4308] <= 16'b0000_0000_0000_0000;
array[4309] <= 16'b0000_0000_0000_0000;
array[4310] <= 16'b0000_0000_0000_0000;
array[4311] <= 16'b0000_0000_0000_0000;
array[4312] <= 16'b0000_0000_0000_0000;
array[4313] <= 16'b0000_0000_0000_0000;
array[4314] <= 16'b0000_0000_0000_0000;
array[4315] <= 16'b0000_0000_0000_0000;
array[4316] <= 16'b0000_0000_0000_0000;
array[4317] <= 16'b0000_0000_0000_0000;
array[4318] <= 16'b0000_0000_0000_0000;
array[4319] <= 16'b0000_0000_0000_0000;
array[4320] <= 16'b0000_0000_0000_0000;
array[4321] <= 16'b0000_0000_0000_0000;
array[4322] <= 16'b0000_0000_0000_0000;
array[4323] <= 16'b0000_0000_0000_0000;
array[4324] <= 16'b0000_0000_0000_0000;
array[4325] <= 16'b0000_0000_0000_0000;
array[4326] <= 16'b0000_0000_0000_0000;
array[4327] <= 16'b0000_0000_0000_0000;
array[4328] <= 16'b0000_0000_0000_0000;
array[4329] <= 16'b0000_0000_0000_0000;
array[4330] <= 16'b0000_0000_0000_0000;
array[4331] <= 16'b0000_0000_0000_0000;
array[4332] <= 16'b0000_0000_0000_0000;
array[4333] <= 16'b0000_0000_0000_0000;
array[4334] <= 16'b0000_0000_0000_0000;
array[4335] <= 16'b0000_0000_0000_0000;
array[4336] <= 16'b0000_0000_0000_0000;
array[4337] <= 16'b0000_0000_0000_0000;
array[4338] <= 16'b0000_0000_0000_0000;
array[4339] <= 16'b0000_0000_0000_0000;
array[4340] <= 16'b0000_0000_0000_0000;
array[4341] <= 16'b0000_0000_0000_0000;
array[4342] <= 16'b0000_0000_0000_0000;
array[4343] <= 16'b0000_0000_0000_0000;
array[4344] <= 16'b0000_0000_0000_0000;
array[4345] <= 16'b0000_0000_0000_0000;
array[4346] <= 16'b0000_0000_0000_0000;
array[4347] <= 16'b0000_0000_0000_0000;
array[4348] <= 16'b0000_0000_0000_0000;
array[4349] <= 16'b0000_0000_0000_0000;
array[4350] <= 16'b0000_0000_0000_0000;
array[4351] <= 16'b0000_0000_0000_0000;
array[4352] <= 16'b0000_0000_0000_0000;
array[4353] <= 16'b0000_0000_0000_0000;
array[4354] <= 16'b0000_0000_0000_0000;
array[4355] <= 16'b0000_0000_0000_0000;
array[4356] <= 16'b0000_0000_0000_0000;
array[4357] <= 16'b0000_0000_0000_0000;
array[4358] <= 16'b0000_0000_0000_0000;
array[4359] <= 16'b0000_0000_0000_0000;
array[4360] <= 16'b0000_0000_0000_0000;
array[4361] <= 16'b0000_0000_0000_0000;
array[4362] <= 16'b0000_0000_0000_0000;
array[4363] <= 16'b0000_0000_0000_0000;
array[4364] <= 16'b0000_0000_0000_0000;
array[4365] <= 16'b0000_0000_0000_0000;
array[4366] <= 16'b0000_0000_0000_0000;
array[4367] <= 16'b0000_0000_0000_0000;
array[4368] <= 16'b0000_0000_0000_0000;
array[4369] <= 16'b0000_0000_0000_0000;
array[4370] <= 16'b0000_0000_0000_0000;
array[4371] <= 16'b0000_0000_0000_0000;
array[4372] <= 16'b0000_0000_0000_0000;
array[4373] <= 16'b0000_0000_0000_0000;
array[4374] <= 16'b0000_0000_0000_0000;
array[4375] <= 16'b0000_0000_0000_0000;
array[4376] <= 16'b0000_0000_0000_0000;
array[4377] <= 16'b0000_0000_0000_0000;
array[4378] <= 16'b0000_0000_0000_0000;
array[4379] <= 16'b0000_0000_0000_0000;
array[4380] <= 16'b0000_0000_0000_0000;
array[4381] <= 16'b0000_0000_0000_0000;
array[4382] <= 16'b0000_0000_0000_0000;
array[4383] <= 16'b0000_0000_0000_0000;
array[4384] <= 16'b0000_0000_0000_0000;
array[4385] <= 16'b0000_0000_0000_0000;
array[4386] <= 16'b0000_0000_0000_0000;
array[4387] <= 16'b0000_0000_0000_0000;
array[4388] <= 16'b0000_0000_0000_0000;
array[4389] <= 16'b0000_0000_0000_0000;
array[4390] <= 16'b0000_0000_0000_0000;
array[4391] <= 16'b0000_0000_0000_0000;
array[4392] <= 16'b0000_0000_0000_0000;
array[4393] <= 16'b0000_0000_0000_0000;
array[4394] <= 16'b0000_0000_0000_0000;
array[4395] <= 16'b0000_0000_0000_0000;
array[4396] <= 16'b0000_0000_0000_0000;
array[4397] <= 16'b0000_0000_0000_0000;
array[4398] <= 16'b0000_0000_0000_0000;
array[4399] <= 16'b0000_0000_0000_0000;
array[4400] <= 16'b0000_0000_0000_0000;
array[4401] <= 16'b0000_0000_0000_0000;
array[4402] <= 16'b0000_0000_0000_0000;
array[4403] <= 16'b0000_0000_0000_0000;
array[4404] <= 16'b0000_0000_0000_0000;
array[4405] <= 16'b0000_0000_0000_0000;
array[4406] <= 16'b0000_0000_0000_0000;
array[4407] <= 16'b0000_0000_0000_0000;
array[4408] <= 16'b0000_0000_0000_0000;
array[4409] <= 16'b0000_0000_0000_0000;
array[4410] <= 16'b0000_0000_0000_0000;
array[4411] <= 16'b0000_0000_0000_0000;
array[4412] <= 16'b0000_0000_0000_0000;
array[4413] <= 16'b0000_0000_0000_0000;
array[4414] <= 16'b0000_0000_0000_0000;
array[4415] <= 16'b0000_0000_0000_0000;
array[4416] <= 16'b0000_0000_0000_0000;
array[4417] <= 16'b0000_0000_0000_0000;
array[4418] <= 16'b0000_0000_0000_0000;
array[4419] <= 16'b0000_0000_0000_0000;
array[4420] <= 16'b0000_0000_0000_0000;
array[4421] <= 16'b0000_0000_0000_0000;
array[4422] <= 16'b0000_0000_0000_0000;
array[4423] <= 16'b0000_0000_0000_0000;
array[4424] <= 16'b0000_0000_0000_0000;
array[4425] <= 16'b0000_0000_0000_0000;
array[4426] <= 16'b0000_0000_0000_0000;
array[4427] <= 16'b0000_0000_0000_0000;
array[4428] <= 16'b0000_0000_0000_0000;
array[4429] <= 16'b0000_0000_0000_0000;
array[4430] <= 16'b0000_0000_0000_0000;
array[4431] <= 16'b0000_0000_0000_0000;
array[4432] <= 16'b0000_0000_0000_0000;
array[4433] <= 16'b0000_0000_0000_0000;
array[4434] <= 16'b0000_0000_0000_0000;
array[4435] <= 16'b0000_0000_0000_0000;
array[4436] <= 16'b0000_0000_0000_0000;
array[4437] <= 16'b0000_0000_0000_0000;
array[4438] <= 16'b0000_0000_0000_0000;
array[4439] <= 16'b0000_0000_0000_0000;
array[4440] <= 16'b0000_0000_0000_0000;
array[4441] <= 16'b0000_0000_0000_0000;
array[4442] <= 16'b0000_0000_0000_0000;
array[4443] <= 16'b0000_0000_0000_0000;
array[4444] <= 16'b0000_0000_0000_0000;
array[4445] <= 16'b0000_0000_0000_0000;
array[4446] <= 16'b0000_0000_0000_0000;
array[4447] <= 16'b0000_0000_0000_0000;
array[4448] <= 16'b0000_0000_0000_0000;
array[4449] <= 16'b0000_0000_0000_0000;
array[4450] <= 16'b0000_0000_0000_0000;
array[4451] <= 16'b0000_0000_0000_0000;
array[4452] <= 16'b0000_0000_0000_0000;
array[4453] <= 16'b0000_0000_0000_0000;
array[4454] <= 16'b0000_0000_0000_0000;
array[4455] <= 16'b0000_0000_0000_0000;
array[4456] <= 16'b0000_0000_0000_0000;
array[4457] <= 16'b0000_0000_0000_0000;
array[4458] <= 16'b0000_0000_0000_0000;
array[4459] <= 16'b0000_0000_0000_0000;
array[4460] <= 16'b0000_0000_0000_0000;
array[4461] <= 16'b0000_0000_0000_0000;
array[4462] <= 16'b0000_0000_0000_0000;
array[4463] <= 16'b0000_0000_0000_0000;
array[4464] <= 16'b0000_0000_0000_0000;
array[4465] <= 16'b0000_0000_0000_0000;
array[4466] <= 16'b0000_0000_0000_0000;
array[4467] <= 16'b0000_0000_0000_0000;
array[4468] <= 16'b0000_0000_0000_0000;
array[4469] <= 16'b0000_0000_0000_0000;
array[4470] <= 16'b0000_0000_0000_0000;
array[4471] <= 16'b0000_0000_0000_0000;
array[4472] <= 16'b0000_0000_0000_0000;
array[4473] <= 16'b0000_0000_0000_0000;
array[4474] <= 16'b0000_0000_0000_0000;
array[4475] <= 16'b0000_0000_0000_0000;
array[4476] <= 16'b0000_0000_0000_0000;
array[4477] <= 16'b0000_0000_0000_0000;
array[4478] <= 16'b0000_0000_0000_0000;
array[4479] <= 16'b0000_0000_0000_0000;
array[4480] <= 16'b0000_0000_0000_0000;
array[4481] <= 16'b0000_0000_0000_0000;
array[4482] <= 16'b0000_0000_0000_0000;
array[4483] <= 16'b0000_0000_0000_0000;
array[4484] <= 16'b0000_0000_0000_0000;
array[4485] <= 16'b0000_0000_0000_0000;
array[4486] <= 16'b0000_0000_0000_0000;
array[4487] <= 16'b0000_0000_0000_0000;
array[4488] <= 16'b0000_0000_0000_0000;
array[4489] <= 16'b0000_0000_0000_0000;
array[4490] <= 16'b0000_0000_0000_0000;
array[4491] <= 16'b0000_0000_0000_0000;
array[4492] <= 16'b0000_0000_0000_0000;
array[4493] <= 16'b0000_0000_0000_0000;
array[4494] <= 16'b0000_0000_0000_0000;
array[4495] <= 16'b0000_0000_0000_0000;
array[4496] <= 16'b0000_0000_0000_0000;
array[4497] <= 16'b0000_0000_0000_0000;
array[4498] <= 16'b0000_0000_0000_0000;
array[4499] <= 16'b0000_0000_0000_0000;
array[4500] <= 16'b0000_0000_0000_0000;
array[4501] <= 16'b0000_0000_0000_0000;
array[4502] <= 16'b0000_0000_0000_0000;
array[4503] <= 16'b0000_0000_0000_0000;
array[4504] <= 16'b0000_0000_0000_0000;
array[4505] <= 16'b0000_0000_0000_0000;
array[4506] <= 16'b0000_0000_0000_0000;
array[4507] <= 16'b0000_0000_0000_0000;
array[4508] <= 16'b0000_0000_0000_0000;
array[4509] <= 16'b0000_0000_0000_0000;
array[4510] <= 16'b0000_0000_0000_0000;
array[4511] <= 16'b0000_0000_0000_0000;
array[4512] <= 16'b0000_0000_0000_0000;
array[4513] <= 16'b0000_0000_0000_0000;
array[4514] <= 16'b0000_0000_0000_0000;
array[4515] <= 16'b0000_0000_0000_0000;
array[4516] <= 16'b0000_0000_0000_0000;
array[4517] <= 16'b0000_0000_0000_0000;
array[4518] <= 16'b0000_0000_0000_0000;
array[4519] <= 16'b0000_0000_0000_0000;
array[4520] <= 16'b0000_0000_0000_0000;
array[4521] <= 16'b0000_0000_0000_0000;
array[4522] <= 16'b0000_0000_0000_0000;
array[4523] <= 16'b0000_0000_0000_0000;
array[4524] <= 16'b0000_0000_0000_0000;
array[4525] <= 16'b0000_0000_0000_0000;
array[4526] <= 16'b0000_0000_0000_0000;
array[4527] <= 16'b0000_0000_0000_0000;
array[4528] <= 16'b0000_0000_0000_0000;
array[4529] <= 16'b0000_0000_0000_0000;
array[4530] <= 16'b0000_0000_0000_0000;
array[4531] <= 16'b0000_0000_0000_0000;
array[4532] <= 16'b0000_0000_0000_0000;
array[4533] <= 16'b0000_0000_0000_0000;
array[4534] <= 16'b0000_0000_0000_0000;
array[4535] <= 16'b0000_0000_0000_0000;
array[4536] <= 16'b0000_0000_0000_0000;
array[4537] <= 16'b0000_0000_0000_0000;
array[4538] <= 16'b0000_0000_0000_0000;
array[4539] <= 16'b0000_0000_0000_0000;
array[4540] <= 16'b0000_0000_0000_0000;
array[4541] <= 16'b0000_0000_0000_0000;
array[4542] <= 16'b0000_0000_0000_0000;
array[4543] <= 16'b0000_0000_0000_0000;
array[4544] <= 16'b0000_0000_0000_0000;
array[4545] <= 16'b0000_0000_0000_0000;
array[4546] <= 16'b0000_0000_0000_0000;
array[4547] <= 16'b0000_0000_0000_0000;
array[4548] <= 16'b0000_0000_0000_0000;
array[4549] <= 16'b0000_0000_0000_0000;
array[4550] <= 16'b0000_0000_0000_0000;
array[4551] <= 16'b0000_0000_0000_0000;
array[4552] <= 16'b0000_0000_0000_0000;
array[4553] <= 16'b0000_0000_0000_0000;
array[4554] <= 16'b0000_0000_0000_0000;
array[4555] <= 16'b0000_0000_0000_0000;
array[4556] <= 16'b0000_0000_0000_0000;
array[4557] <= 16'b0000_0000_0000_0000;
array[4558] <= 16'b0000_0000_0000_0000;
array[4559] <= 16'b0000_0000_0000_0000;
array[4560] <= 16'b0000_0000_0000_0000;
array[4561] <= 16'b0000_0000_0000_0000;
array[4562] <= 16'b0000_0000_0000_0000;
array[4563] <= 16'b0000_0000_0000_0000;
array[4564] <= 16'b0000_0000_0000_0000;
array[4565] <= 16'b0000_0000_0000_0000;
array[4566] <= 16'b0000_0000_0000_0000;
array[4567] <= 16'b0000_0000_0000_0000;
array[4568] <= 16'b0000_0000_0000_0000;
array[4569] <= 16'b0000_0000_0000_0000;
array[4570] <= 16'b0000_0000_0000_0000;
array[4571] <= 16'b0000_0000_0000_0000;
array[4572] <= 16'b0000_0000_0000_0000;
array[4573] <= 16'b0000_0000_0000_0000;
array[4574] <= 16'b0000_0000_0000_0000;
array[4575] <= 16'b0000_0000_0000_0000;
array[4576] <= 16'b0000_0000_0000_0000;
array[4577] <= 16'b0000_0000_0000_0000;
array[4578] <= 16'b0000_0000_0000_0000;
array[4579] <= 16'b0000_0000_0000_0000;
array[4580] <= 16'b0000_0000_0000_0000;
array[4581] <= 16'b0000_0000_0000_0000;
array[4582] <= 16'b0000_0000_0000_0000;
array[4583] <= 16'b0000_0000_0000_0000;
array[4584] <= 16'b0000_0000_0000_0000;
array[4585] <= 16'b0000_0000_0000_0000;
array[4586] <= 16'b0000_0000_0000_0000;
array[4587] <= 16'b0000_0000_0000_0000;
array[4588] <= 16'b0000_0000_0000_0000;
array[4589] <= 16'b0000_0000_0000_0000;
array[4590] <= 16'b0000_0000_0000_0000;
array[4591] <= 16'b0000_0000_0000_0000;
array[4592] <= 16'b0000_0000_0000_0000;
array[4593] <= 16'b0000_0000_0000_0000;
array[4594] <= 16'b0000_0000_0000_0000;
array[4595] <= 16'b0000_0000_0000_0000;
array[4596] <= 16'b0000_0000_0000_0000;
array[4597] <= 16'b0000_0000_0000_0000;
array[4598] <= 16'b0000_0000_0000_0000;
array[4599] <= 16'b0000_0000_0000_0000;
array[4600] <= 16'b0000_0000_0000_0000;
array[4601] <= 16'b0000_0000_0000_0000;
array[4602] <= 16'b0000_0000_0000_0000;
array[4603] <= 16'b0000_0000_0000_0000;
array[4604] <= 16'b0000_0000_0000_0000;
array[4605] <= 16'b0000_0000_0000_0000;
array[4606] <= 16'b0000_0000_0000_0000;
array[4607] <= 16'b0000_0000_0000_0000;
array[4608] <= 16'b0000_0000_0000_0000;
array[4609] <= 16'b0000_0000_0000_0000;
array[4610] <= 16'b0000_0000_0000_0000;
array[4611] <= 16'b0000_0000_0000_0000;
array[4612] <= 16'b0000_0000_0000_0000;
array[4613] <= 16'b0000_0000_0000_0000;
array[4614] <= 16'b0000_0000_0000_0000;
array[4615] <= 16'b0000_0000_0000_0000;
array[4616] <= 16'b0000_0000_0000_0000;
array[4617] <= 16'b0000_0000_0000_0000;
array[4618] <= 16'b0000_0000_0000_0000;
array[4619] <= 16'b0000_0000_0000_0000;
array[4620] <= 16'b0000_0000_0000_0000;
array[4621] <= 16'b0000_0000_0000_0000;
array[4622] <= 16'b0000_0000_0000_0000;
array[4623] <= 16'b0000_0000_0000_0000;
array[4624] <= 16'b0000_0000_0000_0000;
array[4625] <= 16'b0000_0000_0000_0000;
array[4626] <= 16'b0000_0000_0000_0000;
array[4627] <= 16'b0000_0000_0000_0000;
array[4628] <= 16'b0000_0000_0000_0000;
array[4629] <= 16'b0000_0000_0000_0000;
array[4630] <= 16'b0000_0000_0000_0000;
array[4631] <= 16'b0000_0000_0000_0000;
array[4632] <= 16'b0000_0000_0000_0000;
array[4633] <= 16'b0000_0000_0000_0000;
array[4634] <= 16'b0000_0000_0000_0000;
array[4635] <= 16'b0000_0000_0000_0000;
array[4636] <= 16'b0000_0000_0000_0000;
array[4637] <= 16'b0000_0000_0000_0000;
array[4638] <= 16'b0000_0000_0000_0000;
array[4639] <= 16'b0000_0000_0000_0000;
array[4640] <= 16'b0000_0000_0000_0000;
array[4641] <= 16'b0000_0000_0000_0000;
array[4642] <= 16'b0000_0000_0000_0000;
array[4643] <= 16'b0000_0000_0000_0000;
array[4644] <= 16'b0000_0000_0000_0000;
array[4645] <= 16'b0000_0000_0000_0000;
array[4646] <= 16'b0000_0000_0000_0000;
array[4647] <= 16'b0000_0000_0000_0000;
array[4648] <= 16'b0000_0000_0000_0000;
array[4649] <= 16'b0000_0000_0000_0000;
array[4650] <= 16'b0000_0000_0000_0000;
array[4651] <= 16'b0000_0000_0000_0000;
array[4652] <= 16'b0000_0000_0000_0000;
array[4653] <= 16'b0000_0000_0000_0000;
array[4654] <= 16'b0000_0000_0000_0000;
array[4655] <= 16'b0000_0000_0000_0000;
array[4656] <= 16'b0000_0000_0000_0000;
array[4657] <= 16'b0000_0000_0000_0000;
array[4658] <= 16'b0000_0000_0000_0000;
array[4659] <= 16'b0000_0000_0000_0000;
array[4660] <= 16'b0000_0000_0000_0000;
array[4661] <= 16'b0000_0000_0000_0000;
array[4662] <= 16'b0000_0000_0000_0000;
array[4663] <= 16'b0000_0000_0000_0000;
array[4664] <= 16'b0000_0000_0000_0000;
array[4665] <= 16'b0000_0000_0000_0000;
array[4666] <= 16'b0000_0000_0000_0000;
array[4667] <= 16'b0000_0000_0000_0000;
array[4668] <= 16'b0000_0000_0000_0000;
array[4669] <= 16'b0000_0000_0000_0000;
array[4670] <= 16'b0000_0000_0000_0000;
array[4671] <= 16'b0000_0000_0000_0000;
array[4672] <= 16'b0000_0000_0000_0000;
array[4673] <= 16'b0000_0000_0000_0000;
array[4674] <= 16'b0000_0000_0000_0000;
array[4675] <= 16'b0000_0000_0000_0000;
array[4676] <= 16'b0000_0000_0000_0000;
array[4677] <= 16'b0000_0000_0000_0000;
array[4678] <= 16'b0000_0000_0000_0000;
array[4679] <= 16'b0000_0000_0000_0000;
array[4680] <= 16'b0000_0000_0000_0000;
array[4681] <= 16'b0000_0000_0000_0000;
array[4682] <= 16'b0000_0000_0000_0000;
array[4683] <= 16'b0000_0000_0000_0000;
array[4684] <= 16'b0000_0000_0000_0000;
array[4685] <= 16'b0000_0000_0000_0000;
array[4686] <= 16'b0000_0000_0000_0000;
array[4687] <= 16'b0000_0000_0000_0000;
array[4688] <= 16'b0000_0000_0000_0000;
array[4689] <= 16'b0000_0000_0000_0000;
array[4690] <= 16'b0000_0000_0000_0000;
array[4691] <= 16'b0000_0000_0000_0000;
array[4692] <= 16'b0000_0000_0000_0000;
array[4693] <= 16'b0000_0000_0000_0000;
array[4694] <= 16'b0000_0000_0000_0000;
array[4695] <= 16'b0000_0000_0000_0000;
array[4696] <= 16'b0000_0000_0000_0000;
array[4697] <= 16'b0000_0000_0000_0000;
array[4698] <= 16'b0000_0000_0000_0000;
array[4699] <= 16'b0000_0000_0000_0000;
array[4700] <= 16'b0000_0000_0000_0000;
array[4701] <= 16'b0000_0000_0000_0000;
array[4702] <= 16'b0000_0000_0000_0000;
array[4703] <= 16'b0000_0000_0000_0000;
array[4704] <= 16'b0000_0000_0000_0000;
array[4705] <= 16'b0000_0000_0000_0000;
array[4706] <= 16'b0000_0000_0000_0000;
array[4707] <= 16'b0000_0000_0000_0000;
array[4708] <= 16'b0000_0000_0000_0000;
array[4709] <= 16'b0000_0000_0000_0000;
array[4710] <= 16'b0000_0000_0000_0000;
array[4711] <= 16'b0000_0000_0000_0000;
array[4712] <= 16'b0000_0000_0000_0000;
array[4713] <= 16'b0000_0000_0000_0000;
array[4714] <= 16'b0000_0000_0000_0000;
array[4715] <= 16'b0000_0000_0000_0000;
array[4716] <= 16'b0000_0000_0000_0000;
array[4717] <= 16'b0000_0000_0000_0000;
array[4718] <= 16'b0000_0000_0000_0000;
array[4719] <= 16'b0000_0000_0000_0000;
array[4720] <= 16'b0000_0000_0000_0000;
array[4721] <= 16'b0000_0000_0000_0000;
array[4722] <= 16'b0000_0000_0000_0000;
array[4723] <= 16'b0000_0000_0000_0000;
array[4724] <= 16'b0000_0000_0000_0000;
array[4725] <= 16'b0000_0000_0000_0000;
array[4726] <= 16'b0000_0000_0000_0000;
array[4727] <= 16'b0000_0000_0000_0000;
array[4728] <= 16'b0000_0000_0000_0000;
array[4729] <= 16'b0000_0000_0000_0000;
array[4730] <= 16'b0000_0000_0000_0000;
array[4731] <= 16'b0000_0000_0000_0000;
array[4732] <= 16'b0000_0000_0000_0000;
array[4733] <= 16'b0000_0000_0000_0000;
array[4734] <= 16'b0000_0000_0000_0000;
array[4735] <= 16'b0000_0000_0000_0000;
array[4736] <= 16'b0000_0000_0000_0000;
array[4737] <= 16'b0000_0000_0000_0000;
array[4738] <= 16'b0000_0000_0000_0000;
array[4739] <= 16'b0000_0000_0000_0000;
array[4740] <= 16'b0000_0000_0000_0000;
array[4741] <= 16'b0000_0000_0000_0000;
array[4742] <= 16'b0000_0000_0000_0000;
array[4743] <= 16'b0000_0000_0000_0000;
array[4744] <= 16'b0000_0000_0000_0000;
array[4745] <= 16'b0000_0000_0000_0000;
array[4746] <= 16'b0000_0000_0000_0000;
array[4747] <= 16'b0000_0000_0000_0000;
array[4748] <= 16'b0000_0000_0000_0000;
array[4749] <= 16'b0000_0000_0000_0000;
array[4750] <= 16'b0000_0000_0000_0000;
array[4751] <= 16'b0000_0000_0000_0000;
array[4752] <= 16'b0000_0000_0000_0000;
array[4753] <= 16'b0000_0000_0000_0000;
array[4754] <= 16'b0000_0000_0000_0000;
array[4755] <= 16'b0000_0000_0000_0000;
array[4756] <= 16'b0000_0000_0000_0000;
array[4757] <= 16'b0000_0000_0000_0000;
array[4758] <= 16'b0000_0000_0000_0000;
array[4759] <= 16'b0000_0000_0000_0000;
array[4760] <= 16'b0000_0000_0000_0000;
array[4761] <= 16'b0000_0000_0000_0000;
array[4762] <= 16'b0000_0000_0000_0000;
array[4763] <= 16'b0000_0000_0000_0000;
array[4764] <= 16'b0000_0000_0000_0000;
array[4765] <= 16'b0000_0000_0000_0000;
array[4766] <= 16'b0000_0000_0000_0000;
array[4767] <= 16'b0000_0000_0000_0000;
array[4768] <= 16'b0000_0000_0000_0000;
array[4769] <= 16'b0000_0000_0000_0000;
array[4770] <= 16'b0000_0000_0000_0000;
array[4771] <= 16'b0000_0000_0000_0000;
array[4772] <= 16'b0000_0000_0000_0000;
array[4773] <= 16'b0000_0000_0000_0000;
array[4774] <= 16'b0000_0000_0000_0000;
array[4775] <= 16'b0000_0000_0000_0000;
array[4776] <= 16'b0000_0000_0000_0000;
array[4777] <= 16'b0000_0000_0000_0000;
array[4778] <= 16'b0000_0000_0000_0000;
array[4779] <= 16'b0000_0000_0000_0000;
array[4780] <= 16'b0000_0000_0000_0000;
array[4781] <= 16'b0000_0000_0000_0000;
array[4782] <= 16'b0000_0000_0000_0000;
array[4783] <= 16'b0000_0000_0000_0000;
array[4784] <= 16'b0000_0000_0000_0000;
array[4785] <= 16'b0000_0000_0000_0000;
array[4786] <= 16'b0000_0000_0000_0000;
array[4787] <= 16'b0000_0000_0000_0000;
array[4788] <= 16'b0000_0000_0000_0000;
array[4789] <= 16'b0000_0000_0000_0000;
array[4790] <= 16'b0000_0000_0000_0000;
array[4791] <= 16'b0000_0000_0000_0000;
array[4792] <= 16'b0000_0000_0000_0000;
array[4793] <= 16'b0000_0000_0000_0000;
array[4794] <= 16'b0000_0000_0000_0000;
array[4795] <= 16'b0000_0000_0000_0000;
array[4796] <= 16'b0000_0000_0000_0000;
array[4797] <= 16'b0000_0000_0000_0000;
array[4798] <= 16'b0000_0000_0000_0000;
array[4799] <= 16'b0000_0000_0000_0000;
array[4800] <= 16'b0000_0000_0000_0000;
array[4801] <= 16'b0000_0000_0000_0000;
array[4802] <= 16'b0000_0000_0000_0000;
array[4803] <= 16'b0000_0000_0000_0000;
array[4804] <= 16'b0000_0000_0000_0000;
array[4805] <= 16'b0000_0000_0000_0000;
array[4806] <= 16'b0000_0000_0000_0000;
array[4807] <= 16'b0000_0000_0000_0000;
array[4808] <= 16'b0000_0000_0000_0000;
array[4809] <= 16'b0000_0000_0000_0000;
array[4810] <= 16'b0000_0000_0000_0000;
array[4811] <= 16'b0000_0000_0000_0000;
array[4812] <= 16'b0000_0000_0000_0000;
array[4813] <= 16'b0000_0000_0000_0000;
array[4814] <= 16'b0000_0000_0000_0000;
array[4815] <= 16'b0000_0000_0000_0000;
array[4816] <= 16'b0000_0000_0000_0000;
array[4817] <= 16'b0000_0000_0000_0000;
array[4818] <= 16'b0000_0000_0000_0000;
array[4819] <= 16'b0000_0000_0000_0000;
array[4820] <= 16'b0000_0000_0000_0000;
array[4821] <= 16'b0000_0000_0000_0000;
array[4822] <= 16'b0000_0000_0000_0000;
array[4823] <= 16'b0000_0000_0000_0000;
array[4824] <= 16'b0000_0000_0000_0000;
array[4825] <= 16'b0000_0000_0000_0000;
array[4826] <= 16'b0000_0000_0000_0000;
array[4827] <= 16'b0000_0000_0000_0000;
array[4828] <= 16'b0000_0000_0000_0000;
array[4829] <= 16'b0000_0000_0000_0000;
array[4830] <= 16'b0000_0000_0000_0000;
array[4831] <= 16'b0000_0000_0000_0000;
array[4832] <= 16'b0000_0000_0000_0000;
array[4833] <= 16'b0000_0000_0000_0000;
array[4834] <= 16'b0000_0000_0000_0000;
array[4835] <= 16'b0000_0000_0000_0000;
array[4836] <= 16'b0000_0000_0000_0000;
array[4837] <= 16'b0000_0000_0000_0000;
array[4838] <= 16'b0000_0000_0000_0000;
array[4839] <= 16'b0000_0000_0000_0000;
array[4840] <= 16'b0000_0000_0000_0000;
array[4841] <= 16'b0000_0000_0000_0000;
array[4842] <= 16'b0000_0000_0000_0000;
array[4843] <= 16'b0000_0000_0000_0000;
array[4844] <= 16'b0000_0000_0000_0000;
array[4845] <= 16'b0000_0000_0000_0000;
array[4846] <= 16'b0000_0000_0000_0000;
array[4847] <= 16'b0000_0000_0000_0000;
array[4848] <= 16'b0000_0000_0000_0000;
array[4849] <= 16'b0000_0000_0000_0000;
array[4850] <= 16'b0000_0000_0000_0000;
array[4851] <= 16'b0000_0000_0000_0000;
array[4852] <= 16'b0000_0000_0000_0000;
array[4853] <= 16'b0000_0000_0000_0000;
array[4854] <= 16'b0000_0000_0000_0000;
array[4855] <= 16'b0000_0000_0000_0000;
array[4856] <= 16'b0000_0000_0000_0000;
array[4857] <= 16'b0000_0000_0000_0000;
array[4858] <= 16'b0000_0000_0000_0000;
array[4859] <= 16'b0000_0000_0000_0000;
array[4860] <= 16'b0000_0000_0000_0000;
array[4861] <= 16'b0000_0000_0000_0000;
array[4862] <= 16'b0000_0000_0000_0000;
array[4863] <= 16'b0000_0000_0000_0000;
array[4864] <= 16'b0000_0000_0000_0000;
array[4865] <= 16'b0000_0000_0000_0000;
array[4866] <= 16'b0000_0000_0000_0000;
array[4867] <= 16'b0000_0000_0000_0000;
array[4868] <= 16'b0000_0000_0000_0000;
array[4869] <= 16'b0000_0000_0000_0000;
array[4870] <= 16'b0000_0000_0000_0000;
array[4871] <= 16'b0000_0000_0000_0000;
array[4872] <= 16'b0000_0000_0000_0000;
array[4873] <= 16'b0000_0000_0000_0000;
array[4874] <= 16'b0000_0000_0000_0000;
array[4875] <= 16'b0000_0000_0000_0000;
array[4876] <= 16'b0000_0000_0000_0000;
array[4877] <= 16'b0000_0000_0000_0000;
array[4878] <= 16'b0000_0000_0000_0000;
array[4879] <= 16'b0000_0000_0000_0000;
array[4880] <= 16'b0000_0000_0000_0000;
array[4881] <= 16'b0000_0000_0000_0000;
array[4882] <= 16'b0000_0000_0000_0000;
array[4883] <= 16'b0000_0000_0000_0000;
array[4884] <= 16'b0000_0000_0000_0000;
array[4885] <= 16'b0000_0000_0000_0000;
array[4886] <= 16'b0000_0000_0000_0000;
array[4887] <= 16'b0000_0000_0000_0000;
array[4888] <= 16'b0000_0000_0000_0000;
array[4889] <= 16'b0000_0000_0000_0000;
array[4890] <= 16'b0000_0000_0000_0000;
array[4891] <= 16'b0000_0000_0000_0000;
array[4892] <= 16'b0000_0000_0000_0000;
array[4893] <= 16'b0000_0000_0000_0000;
array[4894] <= 16'b0000_0000_0000_0000;
array[4895] <= 16'b0000_0000_0000_0000;
array[4896] <= 16'b0000_0000_0000_0000;
array[4897] <= 16'b0000_0000_0000_0000;
array[4898] <= 16'b0000_0000_0000_0000;
array[4899] <= 16'b0000_0000_0000_0000;
array[4900] <= 16'b0000_0000_0000_0000;
array[4901] <= 16'b0000_0000_0000_0000;
array[4902] <= 16'b0000_0000_0000_0000;
array[4903] <= 16'b0000_0000_0000_0000;
array[4904] <= 16'b0000_0000_0000_0000;
array[4905] <= 16'b0000_0000_0000_0000;
array[4906] <= 16'b0000_0000_0000_0000;
array[4907] <= 16'b0000_0000_0000_0000;
array[4908] <= 16'b0000_0000_0000_0000;
array[4909] <= 16'b0000_0000_0000_0000;
array[4910] <= 16'b0000_0000_0000_0000;
array[4911] <= 16'b0000_0000_0000_0000;
array[4912] <= 16'b0000_0000_0000_0000;
array[4913] <= 16'b0000_0000_0000_0000;
array[4914] <= 16'b0000_0000_0000_0000;
array[4915] <= 16'b0000_0000_0000_0000;
array[4916] <= 16'b0000_0000_0000_0000;
array[4917] <= 16'b0000_0000_0000_0000;
array[4918] <= 16'b0000_0000_0000_0000;
array[4919] <= 16'b0000_0000_0000_0000;
array[4920] <= 16'b0000_0000_0000_0000;
array[4921] <= 16'b0000_0000_0000_0000;
array[4922] <= 16'b0000_0000_0000_0000;
array[4923] <= 16'b0000_0000_0000_0000;
array[4924] <= 16'b0000_0000_0000_0000;
array[4925] <= 16'b0000_0000_0000_0000;
array[4926] <= 16'b0000_0000_0000_0000;
array[4927] <= 16'b0000_0000_0000_0000;
array[4928] <= 16'b0000_0000_0000_0000;
array[4929] <= 16'b0000_0000_0000_0000;
array[4930] <= 16'b0000_0000_0000_0000;
array[4931] <= 16'b0000_0000_0000_0000;
array[4932] <= 16'b0000_0000_0000_0000;
array[4933] <= 16'b0000_0000_0000_0000;
array[4934] <= 16'b0000_0000_0000_0000;
array[4935] <= 16'b0000_0000_0000_0000;
array[4936] <= 16'b0000_0000_0000_0000;
array[4937] <= 16'b0000_0000_0000_0000;
array[4938] <= 16'b0000_0000_0000_0000;
array[4939] <= 16'b0000_0000_0000_0000;
array[4940] <= 16'b0000_0000_0000_0000;
array[4941] <= 16'b0000_0000_0000_0000;
array[4942] <= 16'b0000_0000_0000_0000;
array[4943] <= 16'b0000_0000_0000_0000;
array[4944] <= 16'b0000_0000_0000_0000;
array[4945] <= 16'b0000_0000_0000_0000;
array[4946] <= 16'b0000_0000_0000_0000;
array[4947] <= 16'b0000_0000_0000_0000;
array[4948] <= 16'b0000_0000_0000_0000;
array[4949] <= 16'b0000_0000_0000_0000;
array[4950] <= 16'b0000_0000_0000_0000;
array[4951] <= 16'b0000_0000_0000_0000;
array[4952] <= 16'b0000_0000_0000_0000;
array[4953] <= 16'b0000_0000_0000_0000;
array[4954] <= 16'b0000_0000_0000_0000;
array[4955] <= 16'b0000_0000_0000_0000;
array[4956] <= 16'b0000_0000_0000_0000;
array[4957] <= 16'b0000_0000_0000_0000;
array[4958] <= 16'b0000_0000_0000_0000;
array[4959] <= 16'b0000_0000_0000_0000;
array[4960] <= 16'b0000_0000_0000_0000;
array[4961] <= 16'b0000_0000_0000_0000;
array[4962] <= 16'b0000_0000_0000_0000;
array[4963] <= 16'b0000_0000_0000_0000;
array[4964] <= 16'b0000_0000_0000_0000;
array[4965] <= 16'b0000_0000_0000_0000;
array[4966] <= 16'b0000_0000_0000_0000;
array[4967] <= 16'b0000_0000_0000_0000;
array[4968] <= 16'b0000_0000_0000_0000;
array[4969] <= 16'b0000_0000_0000_0000;
array[4970] <= 16'b0000_0000_0000_0000;
array[4971] <= 16'b0000_0000_0000_0000;
array[4972] <= 16'b0000_0000_0000_0000;
array[4973] <= 16'b0000_0000_0000_0000;
array[4974] <= 16'b0000_0000_0000_0000;
array[4975] <= 16'b0000_0000_0000_0000;
array[4976] <= 16'b0000_0000_0000_0000;
array[4977] <= 16'b0000_0000_0000_0000;
array[4978] <= 16'b0000_0000_0000_0000;
array[4979] <= 16'b0000_0000_0000_0000;
array[4980] <= 16'b0000_0000_0000_0000;
array[4981] <= 16'b0000_0000_0000_0000;
array[4982] <= 16'b0000_0000_0000_0000;
array[4983] <= 16'b0000_0000_0000_0000;
array[4984] <= 16'b0000_0000_0000_0000;
array[4985] <= 16'b0000_0000_0000_0000;
array[4986] <= 16'b0000_0000_0000_0000;
array[4987] <= 16'b0000_0000_0000_0000;
array[4988] <= 16'b0000_0000_0000_0000;
array[4989] <= 16'b0000_0000_0000_0000;
array[4990] <= 16'b0000_0000_0000_0000;
array[4991] <= 16'b0000_0000_0000_0000;
array[4992] <= 16'b0000_0000_0000_0000;
array[4993] <= 16'b0000_0000_0000_0000;
array[4994] <= 16'b0000_0000_0000_0000;
array[4995] <= 16'b0000_0000_0000_0000;
array[4996] <= 16'b0000_0000_0000_0000;
array[4997] <= 16'b0000_0000_0000_0000;
array[4998] <= 16'b0000_0000_0000_0000;
array[4999] <= 16'b0000_0000_0000_0000;
array[5000] <= 16'b0000_0000_0000_0000;
array[5001] <= 16'b0000_0000_0000_0000;
array[5002] <= 16'b0000_0000_0000_0000;
array[5003] <= 16'b0000_0000_0000_0000;
array[5004] <= 16'b0000_0000_0000_0000;
array[5005] <= 16'b0000_0000_0000_0000;
array[5006] <= 16'b0000_0000_0000_0000;
array[5007] <= 16'b0000_0000_0000_0000;
array[5008] <= 16'b0000_0000_0000_0000;
array[5009] <= 16'b0000_0000_0000_0000;
array[5010] <= 16'b0000_0000_0000_0000;
array[5011] <= 16'b0000_0000_0000_0000;
array[5012] <= 16'b0000_0000_0000_0000;
array[5013] <= 16'b0000_0000_0000_0000;
array[5014] <= 16'b0000_0000_0000_0000;
array[5015] <= 16'b0000_0000_0000_0000;
array[5016] <= 16'b0000_0000_0000_0000;
array[5017] <= 16'b0000_0000_0000_0000;
array[5018] <= 16'b0000_0000_0000_0000;
array[5019] <= 16'b0000_0000_0000_0000;
array[5020] <= 16'b0000_0000_0000_0000;
array[5021] <= 16'b0000_0000_0000_0000;
array[5022] <= 16'b0000_0000_0000_0000;
array[5023] <= 16'b0000_0000_0000_0000;
array[5024] <= 16'b0000_0000_0000_0000;
array[5025] <= 16'b0000_0000_0000_0000;
array[5026] <= 16'b0000_0000_0000_0000;
array[5027] <= 16'b0000_0000_0000_0000;
array[5028] <= 16'b0000_0000_0000_0000;
array[5029] <= 16'b0000_0000_0000_0000;
array[5030] <= 16'b0000_0000_0000_0000;
array[5031] <= 16'b0000_0000_0000_0000;
array[5032] <= 16'b0000_0000_0000_0000;
array[5033] <= 16'b0000_0000_0000_0000;
array[5034] <= 16'b0000_0000_0000_0000;
array[5035] <= 16'b0000_0000_0000_0000;
array[5036] <= 16'b0000_0000_0000_0000;
array[5037] <= 16'b0000_0000_0000_0000;
array[5038] <= 16'b0000_0000_0000_0000;
array[5039] <= 16'b0000_0000_0000_0000;
array[5040] <= 16'b0000_0000_0000_0000;
array[5041] <= 16'b0000_0000_0000_0000;
array[5042] <= 16'b0000_0000_0000_0000;
array[5043] <= 16'b0000_0000_0000_0000;
array[5044] <= 16'b0000_0000_0000_0000;
array[5045] <= 16'b0000_0000_0000_0000;
array[5046] <= 16'b0000_0000_0000_0000;
array[5047] <= 16'b0000_0000_0000_0000;
array[5048] <= 16'b0000_0000_0000_0000;
array[5049] <= 16'b0000_0000_0000_0000;
array[5050] <= 16'b0000_0000_0000_0000;
array[5051] <= 16'b0000_0000_0000_0000;
array[5052] <= 16'b0000_0000_0000_0000;
array[5053] <= 16'b0000_0000_0000_0000;
array[5054] <= 16'b0000_0000_0000_0000;
array[5055] <= 16'b0000_0000_0000_0000;
array[5056] <= 16'b0000_0000_0000_0000;
array[5057] <= 16'b0000_0000_0000_0000;
array[5058] <= 16'b0000_0000_0000_0000;
array[5059] <= 16'b0000_0000_0000_0000;
array[5060] <= 16'b0000_0000_0000_0000;
array[5061] <= 16'b0000_0000_0000_0000;
array[5062] <= 16'b0000_0000_0000_0000;
array[5063] <= 16'b0000_0000_0000_0000;
array[5064] <= 16'b0000_0000_0000_0000;
array[5065] <= 16'b0000_0000_0000_0000;
array[5066] <= 16'b0000_0000_0000_0000;
array[5067] <= 16'b0000_0000_0000_0000;
array[5068] <= 16'b0000_0000_0000_0000;
array[5069] <= 16'b0000_0000_0000_0000;
array[5070] <= 16'b0000_0000_0000_0000;
array[5071] <= 16'b0000_0000_0000_0000;
array[5072] <= 16'b0000_0000_0000_0000;
array[5073] <= 16'b0000_0000_0000_0000;
array[5074] <= 16'b0000_0000_0000_0000;
array[5075] <= 16'b0000_0000_0000_0000;
array[5076] <= 16'b0000_0000_0000_0000;
array[5077] <= 16'b0000_0000_0000_0000;
array[5078] <= 16'b0000_0000_0000_0000;
array[5079] <= 16'b0000_0000_0000_0000;
array[5080] <= 16'b0000_0000_0000_0000;
array[5081] <= 16'b0000_0000_0000_0000;
array[5082] <= 16'b0000_0000_0000_0000;
array[5083] <= 16'b0000_0000_0000_0000;
array[5084] <= 16'b0000_0000_0000_0000;
array[5085] <= 16'b0000_0000_0000_0000;
array[5086] <= 16'b0000_0000_0000_0000;
array[5087] <= 16'b0000_0000_0000_0000;
array[5088] <= 16'b0000_0000_0000_0000;
array[5089] <= 16'b0000_0000_0000_0000;
array[5090] <= 16'b0000_0000_0000_0000;
array[5091] <= 16'b0000_0000_0000_0000;
array[5092] <= 16'b0000_0000_0000_0000;
array[5093] <= 16'b0000_0000_0000_0000;
array[5094] <= 16'b0000_0000_0000_0000;
array[5095] <= 16'b0000_0000_0000_0000;
array[5096] <= 16'b0000_0000_0000_0000;
array[5097] <= 16'b0000_0000_0000_0000;
array[5098] <= 16'b0000_0000_0000_0000;
array[5099] <= 16'b0000_0000_0000_0000;
array[5100] <= 16'b0000_0000_0000_0000;
array[5101] <= 16'b0000_0000_0000_0000;
array[5102] <= 16'b0000_0000_0000_0000;
array[5103] <= 16'b0000_0000_0000_0000;
array[5104] <= 16'b0000_0000_0000_0000;
array[5105] <= 16'b0000_0000_0000_0000;
array[5106] <= 16'b0000_0000_0000_0000;
array[5107] <= 16'b0000_0000_0000_0000;
array[5108] <= 16'b0000_0000_0000_0000;
array[5109] <= 16'b0000_0000_0000_0000;
array[5110] <= 16'b0000_0000_0000_0000;
array[5111] <= 16'b0000_0000_0000_0000;
array[5112] <= 16'b0000_0000_0000_0000;
array[5113] <= 16'b0000_0000_0000_0000;
array[5114] <= 16'b0000_0000_0000_0000;
array[5115] <= 16'b0000_0000_0000_0000;
array[5116] <= 16'b0000_0000_0000_0000;
array[5117] <= 16'b0000_0000_0000_0000;
array[5118] <= 16'b0000_0000_0000_0000;
array[5119] <= 16'b0000_0000_0000_0000;
array[5120] <= 16'b0000_0000_0000_0000;
array[5121] <= 16'b0000_0000_0000_0000;
array[5122] <= 16'b0000_0000_0000_0000;
array[5123] <= 16'b0000_0000_0000_0000;
array[5124] <= 16'b0000_0000_0000_0000;
array[5125] <= 16'b0000_0000_0000_0000;
array[5126] <= 16'b0000_0000_0000_0000;
array[5127] <= 16'b0000_0000_0000_0000;
array[5128] <= 16'b0000_0000_0000_0000;
array[5129] <= 16'b0000_0000_0000_0000;
array[5130] <= 16'b0000_0000_0000_0000;
array[5131] <= 16'b0000_0000_0000_0000;
array[5132] <= 16'b0000_0000_0000_0000;
array[5133] <= 16'b0000_0000_0000_0000;
array[5134] <= 16'b0000_0000_0000_0000;
array[5135] <= 16'b0000_0000_0000_0000;
array[5136] <= 16'b0000_0000_0000_0000;
array[5137] <= 16'b0000_0000_0000_0000;
array[5138] <= 16'b0000_0000_0000_0000;
array[5139] <= 16'b0000_0000_0000_0000;
array[5140] <= 16'b0000_0000_0000_0000;
array[5141] <= 16'b0000_0000_0000_0000;
array[5142] <= 16'b0000_0000_0000_0000;
array[5143] <= 16'b0000_0000_0000_0000;
array[5144] <= 16'b0000_0000_0000_0000;
array[5145] <= 16'b0000_0000_0000_0000;
array[5146] <= 16'b0000_0000_0000_0000;
array[5147] <= 16'b0000_0000_0000_0000;
array[5148] <= 16'b0000_0000_0000_0000;
array[5149] <= 16'b0000_0000_0000_0000;
array[5150] <= 16'b0000_0000_0000_0000;
array[5151] <= 16'b0000_0000_0000_0000;
array[5152] <= 16'b0000_0000_0000_0000;
array[5153] <= 16'b0000_0000_0000_0000;
array[5154] <= 16'b0000_0000_0000_0000;
array[5155] <= 16'b0000_0000_0000_0000;
array[5156] <= 16'b0000_0000_0000_0000;
array[5157] <= 16'b0000_0000_0000_0000;
array[5158] <= 16'b0000_0000_0000_0000;
array[5159] <= 16'b0000_0000_0000_0000;
array[5160] <= 16'b0000_0000_0000_0000;
array[5161] <= 16'b0000_0000_0000_0000;
array[5162] <= 16'b0000_0000_0000_0000;
array[5163] <= 16'b0000_0000_0000_0000;
array[5164] <= 16'b0000_0000_0000_0000;
array[5165] <= 16'b0000_0000_0000_0000;
array[5166] <= 16'b0000_0000_0000_0000;
array[5167] <= 16'b0000_0000_0000_0000;
array[5168] <= 16'b0000_0000_0000_0000;
array[5169] <= 16'b0000_0000_0000_0000;
array[5170] <= 16'b0000_0000_0000_0000;
array[5171] <= 16'b0000_0000_0000_0000;
array[5172] <= 16'b0000_0000_0000_0000;
array[5173] <= 16'b0000_0000_0000_0000;
array[5174] <= 16'b0000_0000_0000_0000;
array[5175] <= 16'b0000_0000_0000_0000;
array[5176] <= 16'b0000_0000_0000_0000;
array[5177] <= 16'b0000_0000_0000_0000;
array[5178] <= 16'b0000_0000_0000_0000;
array[5179] <= 16'b0000_0000_0000_0000;
array[5180] <= 16'b0000_0000_0000_0000;
array[5181] <= 16'b0000_0000_0000_0000;
array[5182] <= 16'b0000_0000_0000_0000;
array[5183] <= 16'b0000_0000_0000_0000;
array[5184] <= 16'b0000_0000_0000_0000;
array[5185] <= 16'b0000_0000_0000_0000;
array[5186] <= 16'b0000_0000_0000_0000;
array[5187] <= 16'b0000_0000_0000_0000;
array[5188] <= 16'b0000_0000_0000_0000;
array[5189] <= 16'b0000_0000_0000_0000;
array[5190] <= 16'b0000_0000_0000_0000;
array[5191] <= 16'b0000_0000_0000_0000;
array[5192] <= 16'b0000_0000_0000_0000;
array[5193] <= 16'b0000_0000_0000_0000;
array[5194] <= 16'b0000_0000_0000_0000;
array[5195] <= 16'b0000_0000_0000_0000;
array[5196] <= 16'b0000_0000_0000_0000;
array[5197] <= 16'b0000_0000_0000_0000;
array[5198] <= 16'b0000_0000_0000_0000;
array[5199] <= 16'b0000_0000_0000_0000;
array[5200] <= 16'b0000_0000_0000_0000;
array[5201] <= 16'b0000_0000_0000_0000;
array[5202] <= 16'b0000_0000_0000_0000;
array[5203] <= 16'b0000_0000_0000_0000;
array[5204] <= 16'b0000_0000_0000_0000;
array[5205] <= 16'b0000_0000_0000_0000;
array[5206] <= 16'b0000_0000_0000_0000;
array[5207] <= 16'b0000_0000_0000_0000;
array[5208] <= 16'b0000_0000_0000_0000;
array[5209] <= 16'b0000_0000_0000_0000;
array[5210] <= 16'b0000_0000_0000_0000;
array[5211] <= 16'b0000_0000_0000_0000;
array[5212] <= 16'b0000_0000_0000_0000;
array[5213] <= 16'b0000_0000_0000_0000;
array[5214] <= 16'b0000_0000_0000_0000;
array[5215] <= 16'b0000_0000_0000_0000;
array[5216] <= 16'b0000_0000_0000_0000;
array[5217] <= 16'b0000_0000_0000_0000;
array[5218] <= 16'b0000_0000_0000_0000;
array[5219] <= 16'b0000_0000_0000_0000;
array[5220] <= 16'b0000_0000_0000_0000;
array[5221] <= 16'b0000_0000_0000_0000;
array[5222] <= 16'b0000_0000_0000_0000;
array[5223] <= 16'b0000_0000_0000_0000;
array[5224] <= 16'b0000_0000_0000_0000;
array[5225] <= 16'b0000_0000_0000_0000;
array[5226] <= 16'b0000_0000_0000_0000;
array[5227] <= 16'b0000_0000_0000_0000;
array[5228] <= 16'b0000_0000_0000_0000;
array[5229] <= 16'b0000_0000_0000_0000;
array[5230] <= 16'b0000_0000_0000_0000;
array[5231] <= 16'b0000_0000_0000_0000;
array[5232] <= 16'b0000_0000_0000_0000;
array[5233] <= 16'b0000_0000_0000_0000;
array[5234] <= 16'b0000_0000_0000_0000;
array[5235] <= 16'b0000_0000_0000_0000;
array[5236] <= 16'b0000_0000_0000_0000;
array[5237] <= 16'b0000_0000_0000_0000;
array[5238] <= 16'b0000_0000_0000_0000;
array[5239] <= 16'b0000_0000_0000_0000;
array[5240] <= 16'b0000_0000_0000_0000;
array[5241] <= 16'b0000_0000_0000_0000;
array[5242] <= 16'b0000_0000_0000_0000;
array[5243] <= 16'b0000_0000_0000_0000;
array[5244] <= 16'b0000_0000_0000_0000;
array[5245] <= 16'b0000_0000_0000_0000;
array[5246] <= 16'b0000_0000_0000_0000;
array[5247] <= 16'b0000_0000_0000_0000;
array[5248] <= 16'b0000_0000_0000_0000;
array[5249] <= 16'b0000_0000_0000_0000;
array[5250] <= 16'b0000_0000_0000_0000;
array[5251] <= 16'b0000_0000_0000_0000;
array[5252] <= 16'b0000_0000_0000_0000;
array[5253] <= 16'b0000_0000_0000_0000;
array[5254] <= 16'b0000_0000_0000_0000;
array[5255] <= 16'b0000_0000_0000_0000;
array[5256] <= 16'b0000_0000_0000_0000;
array[5257] <= 16'b0000_0000_0000_0000;
array[5258] <= 16'b0000_0000_0000_0000;
array[5259] <= 16'b0000_0000_0000_0000;
array[5260] <= 16'b0000_0000_0000_0000;
array[5261] <= 16'b0000_0000_0000_0000;
array[5262] <= 16'b0000_0000_0000_0000;
array[5263] <= 16'b0000_0000_0000_0000;
array[5264] <= 16'b0000_0000_0000_0000;
array[5265] <= 16'b0000_0000_0000_0000;
array[5266] <= 16'b0000_0000_0000_0000;
array[5267] <= 16'b0000_0000_0000_0000;
array[5268] <= 16'b0000_0000_0000_0000;
array[5269] <= 16'b0000_0000_0000_0000;
array[5270] <= 16'b0000_0000_0000_0000;
array[5271] <= 16'b0000_0000_0000_0000;
array[5272] <= 16'b0000_0000_0000_0000;
array[5273] <= 16'b0000_0000_0000_0000;
array[5274] <= 16'b0000_0000_0000_0000;
array[5275] <= 16'b0000_0000_0000_0000;
array[5276] <= 16'b0000_0000_0000_0000;
array[5277] <= 16'b0000_0000_0000_0000;
array[5278] <= 16'b0000_0000_0000_0000;
array[5279] <= 16'b0000_0000_0000_0000;
array[5280] <= 16'b0000_0000_0000_0000;
array[5281] <= 16'b0000_0000_0000_0000;
array[5282] <= 16'b0000_0000_0000_0000;
array[5283] <= 16'b0000_0000_0000_0000;
array[5284] <= 16'b0000_0000_0000_0000;
array[5285] <= 16'b0000_0000_0000_0000;
array[5286] <= 16'b0000_0000_0000_0000;
array[5287] <= 16'b0000_0000_0000_0000;
array[5288] <= 16'b0000_0000_0000_0000;
array[5289] <= 16'b0000_0000_0000_0000;
array[5290] <= 16'b0000_0000_0000_0000;
array[5291] <= 16'b0000_0000_0000_0000;
array[5292] <= 16'b0000_0000_0000_0000;
array[5293] <= 16'b0000_0000_0000_0000;
array[5294] <= 16'b0000_0000_0000_0000;
array[5295] <= 16'b0000_0000_0000_0000;
array[5296] <= 16'b0000_0000_0000_0000;
array[5297] <= 16'b0000_0000_0000_0000;
array[5298] <= 16'b0000_0000_0000_0000;
array[5299] <= 16'b0000_0000_0000_0000;
array[5300] <= 16'b0000_0000_0000_0000;
array[5301] <= 16'b0000_0000_0000_0000;
array[5302] <= 16'b0000_0000_0000_0000;
array[5303] <= 16'b0000_0000_0000_0000;
array[5304] <= 16'b0000_0000_0000_0000;
array[5305] <= 16'b0000_0000_0000_0000;
array[5306] <= 16'b0000_0000_0000_0000;
array[5307] <= 16'b0000_0000_0000_0000;
array[5308] <= 16'b0000_0000_0000_0000;
array[5309] <= 16'b0000_0000_0000_0000;
array[5310] <= 16'b0000_0000_0000_0000;
array[5311] <= 16'b0000_0000_0000_0000;
array[5312] <= 16'b0000_0000_0000_0000;
array[5313] <= 16'b0000_0000_0000_0000;
array[5314] <= 16'b0000_0000_0000_0000;
array[5315] <= 16'b0000_0000_0000_0000;
array[5316] <= 16'b0000_0000_0000_0000;
array[5317] <= 16'b0000_0000_0000_0000;
array[5318] <= 16'b0000_0000_0000_0000;
array[5319] <= 16'b0000_0000_0000_0000;
array[5320] <= 16'b0000_0000_0000_0000;
array[5321] <= 16'b0000_0000_0000_0000;
array[5322] <= 16'b0000_0000_0000_0000;
array[5323] <= 16'b0000_0000_0000_0000;
array[5324] <= 16'b0000_0000_0000_0000;
array[5325] <= 16'b0000_0000_0000_0000;
array[5326] <= 16'b0000_0000_0000_0000;
array[5327] <= 16'b0000_0000_0000_0000;
array[5328] <= 16'b0000_0000_0000_0000;
array[5329] <= 16'b0000_0000_0000_0000;
array[5330] <= 16'b0000_0000_0000_0000;
array[5331] <= 16'b0000_0000_0000_0000;
array[5332] <= 16'b0000_0000_0000_0000;
array[5333] <= 16'b0000_0000_0000_0000;
array[5334] <= 16'b0000_0000_0000_0000;
array[5335] <= 16'b0000_0000_0000_0000;
array[5336] <= 16'b0000_0000_0000_0000;
array[5337] <= 16'b0000_0000_0000_0000;
array[5338] <= 16'b0000_0000_0000_0000;
array[5339] <= 16'b0000_0000_0000_0000;
array[5340] <= 16'b0000_0000_0000_0000;
array[5341] <= 16'b0000_0000_0000_0000;
array[5342] <= 16'b0000_0000_0000_0000;
array[5343] <= 16'b0000_0000_0000_0000;
array[5344] <= 16'b0000_0000_0000_0000;
array[5345] <= 16'b0000_0000_0000_0000;
array[5346] <= 16'b0000_0000_0000_0000;
array[5347] <= 16'b0000_0000_0000_0000;
array[5348] <= 16'b0000_0000_0000_0000;
array[5349] <= 16'b0000_0000_0000_0000;
array[5350] <= 16'b0000_0000_0000_0000;
array[5351] <= 16'b0000_0000_0000_0000;
array[5352] <= 16'b0000_0000_0000_0000;
array[5353] <= 16'b0000_0000_0000_0000;
array[5354] <= 16'b0000_0000_0000_0000;
array[5355] <= 16'b0000_0000_0000_0000;
array[5356] <= 16'b0000_0000_0000_0000;
array[5357] <= 16'b0000_0000_0000_0000;
array[5358] <= 16'b0000_0000_0000_0000;
array[5359] <= 16'b0000_0000_0000_0000;
array[5360] <= 16'b0000_0000_0000_0000;
array[5361] <= 16'b0000_0000_0000_0000;
array[5362] <= 16'b0000_0000_0000_0000;
array[5363] <= 16'b0000_0000_0000_0000;
array[5364] <= 16'b0000_0000_0000_0000;
array[5365] <= 16'b0000_0000_0000_0000;
array[5366] <= 16'b0000_0000_0000_0000;
array[5367] <= 16'b0000_0000_0000_0000;
array[5368] <= 16'b0000_0000_0000_0000;
array[5369] <= 16'b0000_0000_0000_0000;
array[5370] <= 16'b0000_0000_0000_0000;
array[5371] <= 16'b0000_0000_0000_0000;
array[5372] <= 16'b0000_0000_0000_0000;
array[5373] <= 16'b0000_0000_0000_0000;
array[5374] <= 16'b0000_0000_0000_0000;
array[5375] <= 16'b0000_0000_0000_0000;
array[5376] <= 16'b0000_0000_0000_0000;
array[5377] <= 16'b0000_0000_0000_0000;
array[5378] <= 16'b0000_0000_0000_0000;
array[5379] <= 16'b0000_0000_0000_0000;
array[5380] <= 16'b0000_0000_0000_0000;
array[5381] <= 16'b0000_0000_0000_0000;
array[5382] <= 16'b0000_0000_0000_0000;
array[5383] <= 16'b0000_0000_0000_0000;
array[5384] <= 16'b0000_0000_0000_0000;
array[5385] <= 16'b0000_0000_0000_0000;
array[5386] <= 16'b0000_0000_0000_0000;
array[5387] <= 16'b0000_0000_0000_0000;
array[5388] <= 16'b0000_0000_0000_0000;
array[5389] <= 16'b0000_0000_0000_0000;
array[5390] <= 16'b0000_0000_0000_0000;
array[5391] <= 16'b0000_0000_0000_0000;
array[5392] <= 16'b0000_0000_0000_0000;
array[5393] <= 16'b0000_0000_0000_0000;
array[5394] <= 16'b0000_0000_0000_0000;
array[5395] <= 16'b0000_0000_0000_0000;
array[5396] <= 16'b0000_0000_0000_0000;
array[5397] <= 16'b0000_0000_0000_0000;
array[5398] <= 16'b0000_0000_0000_0000;
array[5399] <= 16'b0000_0000_0000_0000;
array[5400] <= 16'b0000_0000_0000_0000;
array[5401] <= 16'b0000_0000_0000_0000;
array[5402] <= 16'b0000_0000_0000_0000;
array[5403] <= 16'b0000_0000_0000_0000;
array[5404] <= 16'b0000_0000_0000_0000;
array[5405] <= 16'b0000_0000_0000_0000;
array[5406] <= 16'b0000_0000_0000_0000;
array[5407] <= 16'b0000_0000_0000_0000;
array[5408] <= 16'b0000_0000_0000_0000;
array[5409] <= 16'b0000_0000_0000_0000;
array[5410] <= 16'b0000_0000_0000_0000;
array[5411] <= 16'b0000_0000_0000_0000;
array[5412] <= 16'b0000_0000_0000_0000;
array[5413] <= 16'b0000_0000_0000_0000;
array[5414] <= 16'b0000_0000_0000_0000;
array[5415] <= 16'b0000_0000_0000_0000;
array[5416] <= 16'b0000_0000_0000_0000;
array[5417] <= 16'b0000_0000_0000_0000;
array[5418] <= 16'b0000_0000_0000_0000;
array[5419] <= 16'b0000_0000_0000_0000;
array[5420] <= 16'b0000_0000_0000_0000;
array[5421] <= 16'b0000_0000_0000_0000;
array[5422] <= 16'b0000_0000_0000_0000;
array[5423] <= 16'b0000_0000_0000_0000;
array[5424] <= 16'b0000_0000_0000_0000;
array[5425] <= 16'b0000_0000_0000_0000;
array[5426] <= 16'b0000_0000_0000_0000;
array[5427] <= 16'b0000_0000_0000_0000;
array[5428] <= 16'b0000_0000_0000_0000;
array[5429] <= 16'b0000_0000_0000_0000;
array[5430] <= 16'b0000_0000_0000_0000;
array[5431] <= 16'b0000_0000_0000_0000;
array[5432] <= 16'b0000_0000_0000_0000;
array[5433] <= 16'b0000_0000_0000_0000;
array[5434] <= 16'b0000_0000_0000_0000;
array[5435] <= 16'b0000_0000_0000_0000;
array[5436] <= 16'b0000_0000_0000_0000;
array[5437] <= 16'b0000_0000_0000_0000;
array[5438] <= 16'b0000_0000_0000_0000;
array[5439] <= 16'b0000_0000_0000_0000;
array[5440] <= 16'b0000_0000_0000_0000;
array[5441] <= 16'b0000_0000_0000_0000;
array[5442] <= 16'b0000_0000_0000_0000;
array[5443] <= 16'b0000_0000_0000_0000;
array[5444] <= 16'b0000_0000_0000_0000;
array[5445] <= 16'b0000_0000_0000_0000;
array[5446] <= 16'b0000_0000_0000_0000;
array[5447] <= 16'b0000_0000_0000_0000;
array[5448] <= 16'b0000_0000_0000_0000;
array[5449] <= 16'b0000_0000_0000_0000;
array[5450] <= 16'b0000_0000_0000_0000;
array[5451] <= 16'b0000_0000_0000_0000;
array[5452] <= 16'b0000_0000_0000_0000;
array[5453] <= 16'b0000_0000_0000_0000;
array[5454] <= 16'b0000_0000_0000_0000;
array[5455] <= 16'b0000_0000_0000_0000;
array[5456] <= 16'b0000_0000_0000_0000;
array[5457] <= 16'b0000_0000_0000_0000;
array[5458] <= 16'b0000_0000_0000_0000;
array[5459] <= 16'b0000_0000_0000_0000;
array[5460] <= 16'b0000_0000_0000_0000;
array[5461] <= 16'b0000_0000_0000_0000;
array[5462] <= 16'b0000_0000_0000_0000;
array[5463] <= 16'b0000_0000_0000_0000;
array[5464] <= 16'b0000_0000_0000_0000;
array[5465] <= 16'b0000_0000_0000_0000;
array[5466] <= 16'b0000_0000_0000_0000;
array[5467] <= 16'b0000_0000_0000_0000;
array[5468] <= 16'b0000_0000_0000_0000;
array[5469] <= 16'b0000_0000_0000_0000;
array[5470] <= 16'b0000_0000_0000_0000;
array[5471] <= 16'b0000_0000_0000_0000;
array[5472] <= 16'b0000_0000_0000_0000;
array[5473] <= 16'b0000_0000_0000_0000;
array[5474] <= 16'b0000_0000_0000_0000;
array[5475] <= 16'b0000_0000_0000_0000;
array[5476] <= 16'b0000_0000_0000_0000;
array[5477] <= 16'b0000_0000_0000_0000;
array[5478] <= 16'b0000_0000_0000_0000;
array[5479] <= 16'b0000_0000_0000_0000;
array[5480] <= 16'b0000_0000_0000_0000;
array[5481] <= 16'b0000_0000_0000_0000;
array[5482] <= 16'b0000_0000_0000_0000;
array[5483] <= 16'b0000_0000_0000_0000;
array[5484] <= 16'b0000_0000_0000_0000;
array[5485] <= 16'b0000_0000_0000_0000;
array[5486] <= 16'b0000_0000_0000_0000;
array[5487] <= 16'b0000_0000_0000_0000;
array[5488] <= 16'b0000_0000_0000_0000;
array[5489] <= 16'b0000_0000_0000_0000;
array[5490] <= 16'b0000_0000_0000_0000;
array[5491] <= 16'b0000_0000_0000_0000;
array[5492] <= 16'b0000_0000_0000_0000;
array[5493] <= 16'b0000_0000_0000_0000;
array[5494] <= 16'b0000_0000_0000_0000;
array[5495] <= 16'b0000_0000_0000_0000;
array[5496] <= 16'b0000_0000_0000_0000;
array[5497] <= 16'b0000_0000_0000_0000;
array[5498] <= 16'b0000_0000_0000_0000;
array[5499] <= 16'b0000_0000_0000_0000;
array[5500] <= 16'b0000_0000_0000_0000;
array[5501] <= 16'b0000_0000_0000_0000;
array[5502] <= 16'b0000_0000_0000_0000;
array[5503] <= 16'b0000_0000_0000_0000;
array[5504] <= 16'b0000_0000_0000_0000;
array[5505] <= 16'b0000_0000_0000_0000;
array[5506] <= 16'b0000_0000_0000_0000;
array[5507] <= 16'b0000_0000_0000_0000;
array[5508] <= 16'b0000_0000_0000_0000;
array[5509] <= 16'b0000_0000_0000_0000;
array[5510] <= 16'b0000_0000_0000_0000;
array[5511] <= 16'b0000_0000_0000_0000;
array[5512] <= 16'b0000_0000_0000_0000;
array[5513] <= 16'b0000_0000_0000_0000;
array[5514] <= 16'b0000_0000_0000_0000;
array[5515] <= 16'b0000_0000_0000_0000;
array[5516] <= 16'b0000_0000_0000_0000;
array[5517] <= 16'b0000_0000_0000_0000;
array[5518] <= 16'b0000_0000_0000_0000;
array[5519] <= 16'b0000_0000_0000_0000;
array[5520] <= 16'b0000_0000_0000_0000;
array[5521] <= 16'b0000_0000_0000_0000;
array[5522] <= 16'b0000_0000_0000_0000;
array[5523] <= 16'b0000_0000_0000_0000;
array[5524] <= 16'b0000_0000_0000_0000;
array[5525] <= 16'b0000_0000_0000_0000;
array[5526] <= 16'b0000_0000_0000_0000;
array[5527] <= 16'b0000_0000_0000_0000;
array[5528] <= 16'b0000_0000_0000_0000;
array[5529] <= 16'b0000_0000_0000_0000;
array[5530] <= 16'b0000_0000_0000_0000;
array[5531] <= 16'b0000_0000_0000_0000;
array[5532] <= 16'b0000_0000_0000_0000;
array[5533] <= 16'b0000_0000_0000_0000;
array[5534] <= 16'b0000_0000_0000_0000;
array[5535] <= 16'b0000_0000_0000_0000;
array[5536] <= 16'b0000_0000_0000_0000;
array[5537] <= 16'b0000_0000_0000_0000;
array[5538] <= 16'b0000_0000_0000_0000;
array[5539] <= 16'b0000_0000_0000_0000;
array[5540] <= 16'b0000_0000_0000_0000;
array[5541] <= 16'b0000_0000_0000_0000;
array[5542] <= 16'b0000_0000_0000_0000;
array[5543] <= 16'b0000_0000_0000_0000;
array[5544] <= 16'b0000_0000_0000_0000;
array[5545] <= 16'b0000_0000_0000_0000;
array[5546] <= 16'b0000_0000_0000_0000;
array[5547] <= 16'b0000_0000_0000_0000;
array[5548] <= 16'b0000_0000_0000_0000;
array[5549] <= 16'b0000_0000_0000_0000;
array[5550] <= 16'b0000_0000_0000_0000;
array[5551] <= 16'b0000_0000_0000_0000;
array[5552] <= 16'b0000_0000_0000_0000;
array[5553] <= 16'b0000_0000_0000_0000;
array[5554] <= 16'b0000_0000_0000_0000;
array[5555] <= 16'b0000_0000_0000_0000;
array[5556] <= 16'b0000_0000_0000_0000;
array[5557] <= 16'b0000_0000_0000_0000;
array[5558] <= 16'b0000_0000_0000_0000;
array[5559] <= 16'b0000_0000_0000_0000;
array[5560] <= 16'b0000_0000_0000_0000;
array[5561] <= 16'b0000_0000_0000_0000;
array[5562] <= 16'b0000_0000_0000_0000;
array[5563] <= 16'b0000_0000_0000_0000;
array[5564] <= 16'b0000_0000_0000_0000;
array[5565] <= 16'b0000_0000_0000_0000;
array[5566] <= 16'b0000_0000_0000_0000;
array[5567] <= 16'b0000_0000_0000_0000;
array[5568] <= 16'b0000_0000_0000_0000;
array[5569] <= 16'b0000_0000_0000_0000;
array[5570] <= 16'b0000_0000_0000_0000;
array[5571] <= 16'b0000_0000_0000_0000;
array[5572] <= 16'b0000_0000_0000_0000;
array[5573] <= 16'b0000_0000_0000_0000;
array[5574] <= 16'b0000_0000_0000_0000;
array[5575] <= 16'b0000_0000_0000_0000;
array[5576] <= 16'b0000_0000_0000_0000;
array[5577] <= 16'b0000_0000_0000_0000;
array[5578] <= 16'b0000_0000_0000_0000;
array[5579] <= 16'b0000_0000_0000_0000;
array[5580] <= 16'b0000_0000_0000_0000;
array[5581] <= 16'b0000_0000_0000_0000;
array[5582] <= 16'b0000_0000_0000_0000;
array[5583] <= 16'b0000_0000_0000_0000;
array[5584] <= 16'b0000_0000_0000_0000;
array[5585] <= 16'b0000_0000_0000_0000;
array[5586] <= 16'b0000_0000_0000_0000;
array[5587] <= 16'b0000_0000_0000_0000;
array[5588] <= 16'b0000_0000_0000_0000;
array[5589] <= 16'b0000_0000_0000_0000;
array[5590] <= 16'b0000_0000_0000_0000;
array[5591] <= 16'b0000_0000_0000_0000;
array[5592] <= 16'b0000_0000_0000_0000;
array[5593] <= 16'b0000_0000_0000_0000;
array[5594] <= 16'b0000_0000_0000_0000;
array[5595] <= 16'b0000_0000_0000_0000;
array[5596] <= 16'b0000_0000_0000_0000;
array[5597] <= 16'b0000_0000_0000_0000;
array[5598] <= 16'b0000_0000_0000_0000;
array[5599] <= 16'b0000_0000_0000_0000;
array[5600] <= 16'b0000_0000_0000_0000;
array[5601] <= 16'b0000_0000_0000_0000;
array[5602] <= 16'b0000_0000_0000_0000;
array[5603] <= 16'b0000_0000_0000_0000;
array[5604] <= 16'b0000_0000_0000_0000;
array[5605] <= 16'b0000_0000_0000_0000;
array[5606] <= 16'b0000_0000_0000_0000;
array[5607] <= 16'b0000_0000_0000_0000;
array[5608] <= 16'b0000_0000_0000_0000;
array[5609] <= 16'b0000_0000_0000_0000;
array[5610] <= 16'b0000_0000_0000_0000;
array[5611] <= 16'b0000_0000_0000_0000;
array[5612] <= 16'b0000_0000_0000_0000;
array[5613] <= 16'b0000_0000_0000_0000;
array[5614] <= 16'b0000_0000_0000_0000;
array[5615] <= 16'b0000_0000_0000_0000;
array[5616] <= 16'b0000_0000_0000_0000;
array[5617] <= 16'b0000_0000_0000_0000;
array[5618] <= 16'b0000_0000_0000_0000;
array[5619] <= 16'b0000_0000_0000_0000;
array[5620] <= 16'b0000_0000_0000_0000;
array[5621] <= 16'b0000_0000_0000_0000;
array[5622] <= 16'b0000_0000_0000_0000;
array[5623] <= 16'b0000_0000_0000_0000;
array[5624] <= 16'b0000_0000_0000_0000;
array[5625] <= 16'b0000_0000_0000_0000;
array[5626] <= 16'b0000_0000_0000_0000;
array[5627] <= 16'b0000_0000_0000_0000;
array[5628] <= 16'b0000_0000_0000_0000;
array[5629] <= 16'b0000_0000_0000_0000;
array[5630] <= 16'b0000_0000_0000_0000;
array[5631] <= 16'b0000_0000_0000_0000;
array[5632] <= 16'b0000_0000_0000_0000;
array[5633] <= 16'b0000_0000_0000_0000;
array[5634] <= 16'b0000_0000_0000_0000;
array[5635] <= 16'b0000_0000_0000_0000;
array[5636] <= 16'b0000_0000_0000_0000;
array[5637] <= 16'b0000_0000_0000_0000;
array[5638] <= 16'b0000_0000_0000_0000;
array[5639] <= 16'b0000_0000_0000_0000;
array[5640] <= 16'b0000_0000_0000_0000;
array[5641] <= 16'b0000_0000_0000_0000;
array[5642] <= 16'b0000_0000_0000_0000;
array[5643] <= 16'b0000_0000_0000_0000;
array[5644] <= 16'b0000_0000_0000_0000;
array[5645] <= 16'b0000_0000_0000_0000;
array[5646] <= 16'b0000_0000_0000_0000;
array[5647] <= 16'b0000_0000_0000_0000;
array[5648] <= 16'b0000_0000_0000_0000;
array[5649] <= 16'b0000_0000_0000_0000;
array[5650] <= 16'b0000_0000_0000_0000;
array[5651] <= 16'b0000_0000_0000_0000;
array[5652] <= 16'b0000_0000_0000_0000;
array[5653] <= 16'b0000_0000_0000_0000;
array[5654] <= 16'b0000_0000_0000_0000;
array[5655] <= 16'b0000_0000_0000_0000;
array[5656] <= 16'b0000_0000_0000_0000;
array[5657] <= 16'b0000_0000_0000_0000;
array[5658] <= 16'b0000_0000_0000_0000;
array[5659] <= 16'b0000_0000_0000_0000;
array[5660] <= 16'b0000_0000_0000_0000;
array[5661] <= 16'b0000_0000_0000_0000;
array[5662] <= 16'b0000_0000_0000_0000;
array[5663] <= 16'b0000_0000_0000_0000;
array[5664] <= 16'b0000_0000_0000_0000;
array[5665] <= 16'b0000_0000_0000_0000;
array[5666] <= 16'b0000_0000_0000_0000;
array[5667] <= 16'b0000_0000_0000_0000;
array[5668] <= 16'b0000_0000_0000_0000;
array[5669] <= 16'b0000_0000_0000_0000;
array[5670] <= 16'b0000_0000_0000_0000;
array[5671] <= 16'b0000_0000_0000_0000;
array[5672] <= 16'b0000_0000_0000_0000;
array[5673] <= 16'b0000_0000_0000_0000;
array[5674] <= 16'b0000_0000_0000_0000;
array[5675] <= 16'b0000_0000_0000_0000;
array[5676] <= 16'b0000_0000_0000_0000;
array[5677] <= 16'b0000_0000_0000_0000;
array[5678] <= 16'b0000_0000_0000_0000;
array[5679] <= 16'b0000_0000_0000_0000;
array[5680] <= 16'b0000_0000_0000_0000;
array[5681] <= 16'b0000_0000_0000_0000;
array[5682] <= 16'b0000_0000_0000_0000;
array[5683] <= 16'b0000_0000_0000_0000;
array[5684] <= 16'b0000_0000_0000_0000;
array[5685] <= 16'b0000_0000_0000_0000;
array[5686] <= 16'b0000_0000_0000_0000;
array[5687] <= 16'b0000_0000_0000_0000;
array[5688] <= 16'b0000_0000_0000_0000;
array[5689] <= 16'b0000_0000_0000_0000;
array[5690] <= 16'b0000_0000_0000_0000;
array[5691] <= 16'b0000_0000_0000_0000;
array[5692] <= 16'b0000_0000_0000_0000;
array[5693] <= 16'b0000_0000_0000_0000;
array[5694] <= 16'b0000_0000_0000_0000;
array[5695] <= 16'b0000_0000_0000_0000;
array[5696] <= 16'b0000_0000_0000_0000;
array[5697] <= 16'b0000_0000_0000_0000;
array[5698] <= 16'b0000_0000_0000_0000;
array[5699] <= 16'b0000_0000_0000_0000;
array[5700] <= 16'b0000_0000_0000_0000;
array[5701] <= 16'b0000_0000_0000_0000;
array[5702] <= 16'b0000_0000_0000_0000;
array[5703] <= 16'b0000_0000_0000_0000;
array[5704] <= 16'b0000_0000_0000_0000;
array[5705] <= 16'b0000_0000_0000_0000;
array[5706] <= 16'b0000_0000_0000_0000;
array[5707] <= 16'b0000_0000_0000_0000;
array[5708] <= 16'b0000_0000_0000_0000;
array[5709] <= 16'b0000_0000_0000_0000;
array[5710] <= 16'b0000_0000_0000_0000;
array[5711] <= 16'b0000_0000_0000_0000;
array[5712] <= 16'b0000_0000_0000_0000;
array[5713] <= 16'b0000_0000_0000_0000;
array[5714] <= 16'b0000_0000_0000_0000;
array[5715] <= 16'b0000_0000_0000_0000;
array[5716] <= 16'b0000_0000_0000_0000;
array[5717] <= 16'b0000_0000_0000_0000;
array[5718] <= 16'b0000_0000_0000_0000;
array[5719] <= 16'b0000_0000_0000_0000;
array[5720] <= 16'b0000_0000_0000_0000;
array[5721] <= 16'b0000_0000_0000_0000;
array[5722] <= 16'b0000_0000_0000_0000;
array[5723] <= 16'b0000_0000_0000_0000;
array[5724] <= 16'b0000_0000_0000_0000;
array[5725] <= 16'b0000_0000_0000_0000;
array[5726] <= 16'b0000_0000_0000_0000;
array[5727] <= 16'b0000_0000_0000_0000;
array[5728] <= 16'b0000_0000_0000_0000;
array[5729] <= 16'b0000_0000_0000_0000;
array[5730] <= 16'b0000_0000_0000_0000;
array[5731] <= 16'b0000_0000_0000_0000;
array[5732] <= 16'b0000_0000_0000_0000;
array[5733] <= 16'b0000_0000_0000_0000;
array[5734] <= 16'b0000_0000_0000_0000;
array[5735] <= 16'b0000_0000_0000_0000;
array[5736] <= 16'b0000_0000_0000_0000;
array[5737] <= 16'b0000_0000_0000_0000;
array[5738] <= 16'b0000_0000_0000_0000;
array[5739] <= 16'b0000_0000_0000_0000;
array[5740] <= 16'b0000_0000_0000_0000;
array[5741] <= 16'b0000_0000_0000_0000;
array[5742] <= 16'b0000_0000_0000_0000;
array[5743] <= 16'b0000_0000_0000_0000;
array[5744] <= 16'b0000_0000_0000_0000;
array[5745] <= 16'b0000_0000_0000_0000;
array[5746] <= 16'b0000_0000_0000_0000;
array[5747] <= 16'b0000_0000_0000_0000;
array[5748] <= 16'b0000_0000_0000_0000;
array[5749] <= 16'b0000_0000_0000_0000;
array[5750] <= 16'b0000_0000_0000_0000;
array[5751] <= 16'b0000_0000_0000_0000;
array[5752] <= 16'b0000_0000_0000_0000;
array[5753] <= 16'b0000_0000_0000_0000;
array[5754] <= 16'b0000_0000_0000_0000;
array[5755] <= 16'b0000_0000_0000_0000;
array[5756] <= 16'b0000_0000_0000_0000;
array[5757] <= 16'b0000_0000_0000_0000;
array[5758] <= 16'b0000_0000_0000_0000;
array[5759] <= 16'b0000_0000_0000_0000;
array[5760] <= 16'b0000_0000_0000_0000;
array[5761] <= 16'b0000_0000_0000_0000;
array[5762] <= 16'b0000_0000_0000_0000;
array[5763] <= 16'b0000_0000_0000_0000;
array[5764] <= 16'b0000_0000_0000_0000;
array[5765] <= 16'b0000_0000_0000_0000;
array[5766] <= 16'b0000_0000_0000_0000;
array[5767] <= 16'b0000_0000_0000_0000;
array[5768] <= 16'b0000_0000_0000_0000;
array[5769] <= 16'b0000_0000_0000_0000;
array[5770] <= 16'b0000_0000_0000_0000;
array[5771] <= 16'b0000_0000_0000_0000;
array[5772] <= 16'b0000_0000_0000_0000;
array[5773] <= 16'b0000_0000_0000_0000;
array[5774] <= 16'b0000_0000_0000_0000;
array[5775] <= 16'b0000_0000_0000_0000;
array[5776] <= 16'b0000_0000_0000_0000;
array[5777] <= 16'b0000_0000_0000_0000;
array[5778] <= 16'b0000_0000_0000_0000;
array[5779] <= 16'b0000_0000_0000_0000;
array[5780] <= 16'b0000_0000_0000_0000;
array[5781] <= 16'b0000_0000_0000_0000;
array[5782] <= 16'b0000_0000_0000_0000;
array[5783] <= 16'b0000_0000_0000_0000;
array[5784] <= 16'b0000_0000_0000_0000;
array[5785] <= 16'b0000_0000_0000_0000;
array[5786] <= 16'b0000_0000_0000_0000;
array[5787] <= 16'b0000_0000_0000_0000;
array[5788] <= 16'b0000_0000_0000_0000;
array[5789] <= 16'b0000_0000_0000_0000;
array[5790] <= 16'b0000_0000_0000_0000;
array[5791] <= 16'b0000_0000_0000_0000;
array[5792] <= 16'b0000_0000_0000_0000;
array[5793] <= 16'b0000_0000_0000_0000;
array[5794] <= 16'b0000_0000_0000_0000;
array[5795] <= 16'b0000_0000_0000_0000;
array[5796] <= 16'b0000_0000_0000_0000;
array[5797] <= 16'b0000_0000_0000_0000;
array[5798] <= 16'b0000_0000_0000_0000;
array[5799] <= 16'b0000_0000_0000_0000;
array[5800] <= 16'b0000_0000_0000_0000;
array[5801] <= 16'b0000_0000_0000_0000;
array[5802] <= 16'b0000_0000_0000_0000;
array[5803] <= 16'b0000_0000_0000_0000;
array[5804] <= 16'b0000_0000_0000_0000;
array[5805] <= 16'b0000_0000_0000_0000;
array[5806] <= 16'b0000_0000_0000_0000;
array[5807] <= 16'b0000_0000_0000_0000;
array[5808] <= 16'b0000_0000_0000_0000;
array[5809] <= 16'b0000_0000_0000_0000;
array[5810] <= 16'b0000_0000_0000_0000;
array[5811] <= 16'b0000_0000_0000_0000;
array[5812] <= 16'b0000_0000_0000_0000;
array[5813] <= 16'b0000_0000_0000_0000;
array[5814] <= 16'b0000_0000_0000_0000;
array[5815] <= 16'b0000_0000_0000_0000;
array[5816] <= 16'b0000_0000_0000_0000;
array[5817] <= 16'b0000_0000_0000_0000;
array[5818] <= 16'b0000_0000_0000_0000;
array[5819] <= 16'b0000_0000_0000_0000;
array[5820] <= 16'b0000_0000_0000_0000;
array[5821] <= 16'b0000_0000_0000_0000;
array[5822] <= 16'b0000_0000_0000_0000;
array[5823] <= 16'b0000_0000_0000_0000;
array[5824] <= 16'b0000_0000_0000_0000;
array[5825] <= 16'b0000_0000_0000_0000;
array[5826] <= 16'b0000_0000_0000_0000;
array[5827] <= 16'b0000_0000_0000_0000;
array[5828] <= 16'b0000_0000_0000_0000;
array[5829] <= 16'b0000_0000_0000_0000;
array[5830] <= 16'b0000_0000_0000_0000;
array[5831] <= 16'b0000_0000_0000_0000;
array[5832] <= 16'b0000_0000_0000_0000;
array[5833] <= 16'b0000_0000_0000_0000;
array[5834] <= 16'b0000_0000_0000_0000;
array[5835] <= 16'b0000_0000_0000_0000;
array[5836] <= 16'b0000_0000_0000_0000;
array[5837] <= 16'b0000_0000_0000_0000;
array[5838] <= 16'b0000_0000_0000_0000;
array[5839] <= 16'b0000_0000_0000_0000;
array[5840] <= 16'b0000_0000_0000_0000;
array[5841] <= 16'b0000_0000_0000_0000;
array[5842] <= 16'b0000_0000_0000_0000;
array[5843] <= 16'b0000_0000_0000_0000;
array[5844] <= 16'b0000_0000_0000_0000;
array[5845] <= 16'b0000_0000_0000_0000;
array[5846] <= 16'b0000_0000_0000_0000;
array[5847] <= 16'b0000_0000_0000_0000;
array[5848] <= 16'b0000_0000_0000_0000;
array[5849] <= 16'b0000_0000_0000_0000;
array[5850] <= 16'b0000_0000_0000_0000;
array[5851] <= 16'b0000_0000_0000_0000;
array[5852] <= 16'b0000_0000_0000_0000;
array[5853] <= 16'b0000_0000_0000_0000;
array[5854] <= 16'b0000_0000_0000_0000;
array[5855] <= 16'b0000_0000_0000_0000;
array[5856] <= 16'b0000_0000_0000_0000;
array[5857] <= 16'b0000_0000_0000_0000;
array[5858] <= 16'b0000_0000_0000_0000;
array[5859] <= 16'b0000_0000_0000_0000;
array[5860] <= 16'b0000_0000_0000_0000;
array[5861] <= 16'b0000_0000_0000_0000;
array[5862] <= 16'b0000_0000_0000_0000;
array[5863] <= 16'b0000_0000_0000_0000;
array[5864] <= 16'b0000_0000_0000_0000;
array[5865] <= 16'b0000_0000_0000_0000;
array[5866] <= 16'b0000_0000_0000_0000;
array[5867] <= 16'b0000_0000_0000_0000;
array[5868] <= 16'b0000_0000_0000_0000;
array[5869] <= 16'b0000_0000_0000_0000;
array[5870] <= 16'b0000_0000_0000_0000;
array[5871] <= 16'b0000_0000_0000_0000;
array[5872] <= 16'b0000_0000_0000_0000;
array[5873] <= 16'b0000_0000_0000_0000;
array[5874] <= 16'b0000_0000_0000_0000;
array[5875] <= 16'b0000_0000_0000_0000;
array[5876] <= 16'b0000_0000_0000_0000;
array[5877] <= 16'b0000_0000_0000_0000;
array[5878] <= 16'b0000_0000_0000_0000;
array[5879] <= 16'b0000_0000_0000_0000;
array[5880] <= 16'b0000_0000_0000_0000;
array[5881] <= 16'b0000_0000_0000_0000;
array[5882] <= 16'b0000_0000_0000_0000;
array[5883] <= 16'b0000_0000_0000_0000;
array[5884] <= 16'b0000_0000_0000_0000;
array[5885] <= 16'b0000_0000_0000_0000;
array[5886] <= 16'b0000_0000_0000_0000;
array[5887] <= 16'b0000_0000_0000_0000;
array[5888] <= 16'b0000_0000_0000_0000;
array[5889] <= 16'b0000_0000_0000_0000;
array[5890] <= 16'b0000_0000_0000_0000;
array[5891] <= 16'b0000_0000_0000_0000;
array[5892] <= 16'b0000_0000_0000_0000;
array[5893] <= 16'b0000_0000_0000_0000;
array[5894] <= 16'b0000_0000_0000_0000;
array[5895] <= 16'b0000_0000_0000_0000;
array[5896] <= 16'b0000_0000_0000_0000;
array[5897] <= 16'b0000_0000_0000_0000;
array[5898] <= 16'b0000_0000_0000_0000;
array[5899] <= 16'b0000_0000_0000_0000;
array[5900] <= 16'b0000_0000_0000_0000;
array[5901] <= 16'b0000_0000_0000_0000;
array[5902] <= 16'b0000_0000_0000_0000;
array[5903] <= 16'b0000_0000_0000_0000;
array[5904] <= 16'b0000_0000_0000_0000;
array[5905] <= 16'b0000_0000_0000_0000;
array[5906] <= 16'b0000_0000_0000_0000;
array[5907] <= 16'b0000_0000_0000_0000;
array[5908] <= 16'b0000_0000_0000_0000;
array[5909] <= 16'b0000_0000_0000_0000;
array[5910] <= 16'b0000_0000_0000_0000;
array[5911] <= 16'b0000_0000_0000_0000;
array[5912] <= 16'b0000_0000_0000_0000;
array[5913] <= 16'b0000_0000_0000_0000;
array[5914] <= 16'b0000_0000_0000_0000;
array[5915] <= 16'b0000_0000_0000_0000;
array[5916] <= 16'b0000_0000_0000_0000;
array[5917] <= 16'b0000_0000_0000_0000;
array[5918] <= 16'b0000_0000_0000_0000;
array[5919] <= 16'b0000_0000_0000_0000;
array[5920] <= 16'b0000_0000_0000_0000;
array[5921] <= 16'b0000_0000_0000_0000;
array[5922] <= 16'b0000_0000_0000_0000;
array[5923] <= 16'b0000_0000_0000_0000;
array[5924] <= 16'b0000_0000_0000_0000;
array[5925] <= 16'b0000_0000_0000_0000;
array[5926] <= 16'b0000_0000_0000_0000;
array[5927] <= 16'b0000_0000_0000_0000;
array[5928] <= 16'b0000_0000_0000_0000;
array[5929] <= 16'b0000_0000_0000_0000;
array[5930] <= 16'b0000_0000_0000_0000;
array[5931] <= 16'b0000_0000_0000_0000;
array[5932] <= 16'b0000_0000_0000_0000;
array[5933] <= 16'b0000_0000_0000_0000;
array[5934] <= 16'b0000_0000_0000_0000;
array[5935] <= 16'b0000_0000_0000_0000;
array[5936] <= 16'b0000_0000_0000_0000;
array[5937] <= 16'b0000_0000_0000_0000;
array[5938] <= 16'b0000_0000_0000_0000;
array[5939] <= 16'b0000_0000_0000_0000;
array[5940] <= 16'b0000_0000_0000_0000;
array[5941] <= 16'b0000_0000_0000_0000;
array[5942] <= 16'b0000_0000_0000_0000;
array[5943] <= 16'b0000_0000_0000_0000;
array[5944] <= 16'b0000_0000_0000_0000;
array[5945] <= 16'b0000_0000_0000_0000;
array[5946] <= 16'b0000_0000_0000_0000;
array[5947] <= 16'b0000_0000_0000_0000;
array[5948] <= 16'b0000_0000_0000_0000;
array[5949] <= 16'b0000_0000_0000_0000;
array[5950] <= 16'b0000_0000_0000_0000;
array[5951] <= 16'b0000_0000_0000_0000;
array[5952] <= 16'b0000_0000_0000_0000;
array[5953] <= 16'b0000_0000_0000_0000;
array[5954] <= 16'b0000_0000_0000_0000;
array[5955] <= 16'b0000_0000_0000_0000;
array[5956] <= 16'b0000_0000_0000_0000;
array[5957] <= 16'b0000_0000_0000_0000;
array[5958] <= 16'b0000_0000_0000_0000;
array[5959] <= 16'b0000_0000_0000_0000;
array[5960] <= 16'b0000_0000_0000_0000;
array[5961] <= 16'b0000_0000_0000_0000;
array[5962] <= 16'b0000_0000_0000_0000;
array[5963] <= 16'b0000_0000_0000_0000;
array[5964] <= 16'b0000_0000_0000_0000;
array[5965] <= 16'b0000_0000_0000_0000;
array[5966] <= 16'b0000_0000_0000_0000;
array[5967] <= 16'b0000_0000_0000_0000;
array[5968] <= 16'b0000_0000_0000_0000;
array[5969] <= 16'b0000_0000_0000_0000;
array[5970] <= 16'b0000_0000_0000_0000;
array[5971] <= 16'b0000_0000_0000_0000;
array[5972] <= 16'b0000_0000_0000_0000;
array[5973] <= 16'b0000_0000_0000_0000;
array[5974] <= 16'b0000_0000_0000_0000;
array[5975] <= 16'b0000_0000_0000_0000;
array[5976] <= 16'b0000_0000_0000_0000;
array[5977] <= 16'b0000_0000_0000_0000;
array[5978] <= 16'b0000_0000_0000_0000;
array[5979] <= 16'b0000_0000_0000_0000;
array[5980] <= 16'b0000_0000_0000_0000;
array[5981] <= 16'b0000_0000_0000_0000;
array[5982] <= 16'b0000_0000_0000_0000;
array[5983] <= 16'b0000_0000_0000_0000;
array[5984] <= 16'b0000_0000_0000_0000;
array[5985] <= 16'b0000_0000_0000_0000;
array[5986] <= 16'b0000_0000_0000_0000;
array[5987] <= 16'b0000_0000_0000_0000;
array[5988] <= 16'b0000_0000_0000_0000;
array[5989] <= 16'b0000_0000_0000_0000;
array[5990] <= 16'b0000_0000_0000_0000;
array[5991] <= 16'b0000_0000_0000_0000;
array[5992] <= 16'b0000_0000_0000_0000;
array[5993] <= 16'b0000_0000_0000_0000;
array[5994] <= 16'b0000_0000_0000_0000;
array[5995] <= 16'b0000_0000_0000_0000;
array[5996] <= 16'b0000_0000_0000_0000;
array[5997] <= 16'b0000_0000_0000_0000;
array[5998] <= 16'b0000_0000_0000_0000;
array[5999] <= 16'b0000_0000_0000_0000;
array[6000] <= 16'b0000_0000_0000_0000;
array[6001] <= 16'b0000_0000_0000_0000;
array[6002] <= 16'b0000_0000_0000_0000;
array[6003] <= 16'b0000_0000_0000_0000;
array[6004] <= 16'b0000_0000_0000_0000;
array[6005] <= 16'b0000_0000_0000_0000;
array[6006] <= 16'b0000_0000_0000_0000;
array[6007] <= 16'b0000_0000_0000_0000;
array[6008] <= 16'b0000_0000_0000_0000;
array[6009] <= 16'b0000_0000_0000_0000;
array[6010] <= 16'b0000_0000_0000_0000;
array[6011] <= 16'b0000_0000_0000_0000;
array[6012] <= 16'b0000_0000_0000_0000;
array[6013] <= 16'b0000_0000_0000_0000;
array[6014] <= 16'b0000_0000_0000_0000;
array[6015] <= 16'b0000_0000_0000_0000;
array[6016] <= 16'b0000_0000_0000_0000;
array[6017] <= 16'b0000_0000_0000_0000;
array[6018] <= 16'b0000_0000_0000_0000;
array[6019] <= 16'b0000_0000_0000_0000;
array[6020] <= 16'b0000_0000_0000_0000;
array[6021] <= 16'b0000_0000_0000_0000;
array[6022] <= 16'b0000_0000_0000_0000;
array[6023] <= 16'b0000_0000_0000_0000;
array[6024] <= 16'b0000_0000_0000_0000;
array[6025] <= 16'b0000_0000_0000_0000;
array[6026] <= 16'b0000_0000_0000_0000;
array[6027] <= 16'b0000_0000_0000_0000;
array[6028] <= 16'b0000_0000_0000_0000;
array[6029] <= 16'b0000_0000_0000_0000;
array[6030] <= 16'b0000_0000_0000_0000;
array[6031] <= 16'b0000_0000_0000_0000;
array[6032] <= 16'b0000_0000_0000_0000;
array[6033] <= 16'b0000_0000_0000_0000;
array[6034] <= 16'b0000_0000_0000_0000;
array[6035] <= 16'b0000_0000_0000_0000;
array[6036] <= 16'b0000_0000_0000_0000;
array[6037] <= 16'b0000_0000_0000_0000;
array[6038] <= 16'b0000_0000_0000_0000;
array[6039] <= 16'b0000_0000_0000_0000;
array[6040] <= 16'b0000_0000_0000_0000;
array[6041] <= 16'b0000_0000_0000_0000;
array[6042] <= 16'b0000_0000_0000_0000;
array[6043] <= 16'b0000_0000_0000_0000;
array[6044] <= 16'b0000_0000_0000_0000;
array[6045] <= 16'b0000_0000_0000_0000;
array[6046] <= 16'b0000_0000_0000_0000;
array[6047] <= 16'b0000_0000_0000_0000;
array[6048] <= 16'b0000_0000_0000_0000;
array[6049] <= 16'b0000_0000_0000_0000;
array[6050] <= 16'b0000_0000_0000_0000;
array[6051] <= 16'b0000_0000_0000_0000;
array[6052] <= 16'b0000_0000_0000_0000;
array[6053] <= 16'b0000_0000_0000_0000;
array[6054] <= 16'b0000_0000_0000_0000;
array[6055] <= 16'b0000_0000_0000_0000;
array[6056] <= 16'b0000_0000_0000_0000;
array[6057] <= 16'b0000_0000_0000_0000;
array[6058] <= 16'b0000_0000_0000_0000;
array[6059] <= 16'b0000_0000_0000_0000;
array[6060] <= 16'b0000_0000_0000_0000;
array[6061] <= 16'b0000_0000_0000_0000;
array[6062] <= 16'b0000_0000_0000_0000;
array[6063] <= 16'b0000_0000_0000_0000;
array[6064] <= 16'b0000_0000_0000_0000;
array[6065] <= 16'b0000_0000_0000_0000;
array[6066] <= 16'b0000_0000_0000_0000;
array[6067] <= 16'b0000_0000_0000_0000;
array[6068] <= 16'b0000_0000_0000_0000;
array[6069] <= 16'b0000_0000_0000_0000;
array[6070] <= 16'b0000_0000_0000_0000;
array[6071] <= 16'b0000_0000_0000_0000;
array[6072] <= 16'b0000_0000_0000_0000;
array[6073] <= 16'b0000_0000_0000_0000;
array[6074] <= 16'b0000_0000_0000_0000;
array[6075] <= 16'b0000_0000_0000_0000;
array[6076] <= 16'b0000_0000_0000_0000;
array[6077] <= 16'b0000_0000_0000_0000;
array[6078] <= 16'b0000_0000_0000_0000;
array[6079] <= 16'b0000_0000_0000_0000;
array[6080] <= 16'b0000_0000_0000_0000;
array[6081] <= 16'b0000_0000_0000_0000;
array[6082] <= 16'b0000_0000_0000_0000;
array[6083] <= 16'b0000_0000_0000_0000;
array[6084] <= 16'b0000_0000_0000_0000;
array[6085] <= 16'b0000_0000_0000_0000;
array[6086] <= 16'b0000_0000_0000_0000;
array[6087] <= 16'b0000_0000_0000_0000;
array[6088] <= 16'b0000_0000_0000_0000;
array[6089] <= 16'b0000_0000_0000_0000;
array[6090] <= 16'b0000_0000_0000_0000;
array[6091] <= 16'b0000_0000_0000_0000;
array[6092] <= 16'b0000_0000_0000_0000;
array[6093] <= 16'b0000_0000_0000_0000;
array[6094] <= 16'b0000_0000_0000_0000;
array[6095] <= 16'b0000_0000_0000_0000;
array[6096] <= 16'b0000_0000_0000_0000;
array[6097] <= 16'b0000_0000_0000_0000;
array[6098] <= 16'b0000_0000_0000_0000;
array[6099] <= 16'b0000_0000_0000_0000;
array[6100] <= 16'b0000_0000_0000_0000;
array[6101] <= 16'b0000_0000_0000_0000;
array[6102] <= 16'b0000_0000_0000_0000;
array[6103] <= 16'b0000_0000_0000_0000;
array[6104] <= 16'b0000_0000_0000_0000;
array[6105] <= 16'b0000_0000_0000_0000;
array[6106] <= 16'b0000_0000_0000_0000;
array[6107] <= 16'b0000_0000_0000_0000;
array[6108] <= 16'b0000_0000_0000_0000;
array[6109] <= 16'b0000_0000_0000_0000;
array[6110] <= 16'b0000_0000_0000_0000;
array[6111] <= 16'b0000_0000_0000_0000;
array[6112] <= 16'b0000_0000_0000_0000;
array[6113] <= 16'b0000_0000_0000_0000;
array[6114] <= 16'b0000_0000_0000_0000;
array[6115] <= 16'b0000_0000_0000_0000;
array[6116] <= 16'b0000_0000_0000_0000;
array[6117] <= 16'b0000_0000_0000_0000;
array[6118] <= 16'b0000_0000_0000_0000;
array[6119] <= 16'b0000_0000_0000_0000;
array[6120] <= 16'b0000_0000_0000_0000;
array[6121] <= 16'b0000_0000_0000_0000;
array[6122] <= 16'b0000_0000_0000_0000;
array[6123] <= 16'b0000_0000_0000_0000;
array[6124] <= 16'b0000_0000_0000_0000;
array[6125] <= 16'b0000_0000_0000_0000;
array[6126] <= 16'b0000_0000_0000_0000;
array[6127] <= 16'b0000_0000_0000_0000;
array[6128] <= 16'b0000_0000_0000_0000;
array[6129] <= 16'b0000_0000_0000_0000;
array[6130] <= 16'b0000_0000_0000_0000;
array[6131] <= 16'b0000_0000_0000_0000;
array[6132] <= 16'b0000_0000_0000_0000;
array[6133] <= 16'b0000_0000_0000_0000;
array[6134] <= 16'b0000_0000_0000_0000;
array[6135] <= 16'b0000_0000_0000_0000;
array[6136] <= 16'b0000_0000_0000_0000;
array[6137] <= 16'b0000_0000_0000_0000;
array[6138] <= 16'b0000_0000_0000_0000;
array[6139] <= 16'b0000_0000_0000_0000;
array[6140] <= 16'b0000_0000_0000_0000;
array[6141] <= 16'b0000_0000_0000_0000;
array[6142] <= 16'b0000_0000_0000_0000;
array[6143] <= 16'b0000_0000_0000_0000;
array[6144] <= 16'b0000_0000_0000_0000;
array[6145] <= 16'b0000_0000_0000_0000;
array[6146] <= 16'b0000_0000_0000_0000;
array[6147] <= 16'b0000_0000_0000_0000;
array[6148] <= 16'b0000_0000_0000_0000;
array[6149] <= 16'b0000_0000_0000_0000;
array[6150] <= 16'b0000_0000_0000_0000;
array[6151] <= 16'b0000_0000_0000_0000;
array[6152] <= 16'b0000_0000_0000_0000;
array[6153] <= 16'b0000_0000_0000_0000;
array[6154] <= 16'b0000_0000_0000_0000;
array[6155] <= 16'b0000_0000_0000_0000;
array[6156] <= 16'b0000_0000_0000_0000;
array[6157] <= 16'b0000_0000_0000_0000;
array[6158] <= 16'b0000_0000_0000_0000;
array[6159] <= 16'b0000_0000_0000_0000;
array[6160] <= 16'b0000_0000_0000_0000;
array[6161] <= 16'b0000_0000_0000_0000;
array[6162] <= 16'b0000_0000_0000_0000;
array[6163] <= 16'b0000_0000_0000_0000;
array[6164] <= 16'b0000_0000_0000_0000;
array[6165] <= 16'b0000_0000_0000_0000;
array[6166] <= 16'b0000_0000_0000_0000;
array[6167] <= 16'b0000_0000_0000_0000;
array[6168] <= 16'b0000_0000_0000_0000;
array[6169] <= 16'b0000_0000_0000_0000;
array[6170] <= 16'b0000_0000_0000_0000;
array[6171] <= 16'b0000_0000_0000_0000;
array[6172] <= 16'b0000_0000_0000_0000;
array[6173] <= 16'b0000_0000_0000_0000;
array[6174] <= 16'b0000_0000_0000_0000;
array[6175] <= 16'b0000_0000_0000_0000;
array[6176] <= 16'b0000_0000_0000_0000;
array[6177] <= 16'b0000_0000_0000_0000;
array[6178] <= 16'b0000_0000_0000_0000;
array[6179] <= 16'b0000_0000_0000_0000;
array[6180] <= 16'b0000_0000_0000_0000;
array[6181] <= 16'b0000_0000_0000_0000;
array[6182] <= 16'b0000_0000_0000_0000;
array[6183] <= 16'b0000_0000_0000_0000;
array[6184] <= 16'b0000_0000_0000_0000;
array[6185] <= 16'b0000_0000_0000_0000;
array[6186] <= 16'b0000_0000_0000_0000;
array[6187] <= 16'b0000_0000_0000_0000;
array[6188] <= 16'b0000_0000_0000_0000;
array[6189] <= 16'b0000_0000_0000_0000;
array[6190] <= 16'b0000_0000_0000_0000;
array[6191] <= 16'b0000_0000_0000_0000;
array[6192] <= 16'b0000_0000_0000_0000;
array[6193] <= 16'b0000_0000_0000_0000;
array[6194] <= 16'b0000_0000_0000_0000;
array[6195] <= 16'b0000_0000_0000_0000;
array[6196] <= 16'b0000_0000_0000_0000;
array[6197] <= 16'b0000_0000_0000_0000;
array[6198] <= 16'b0000_0000_0000_0000;
array[6199] <= 16'b0000_0000_0000_0000;
array[6200] <= 16'b0000_0000_0000_0000;
array[6201] <= 16'b0000_0000_0000_0000;
array[6202] <= 16'b0000_0000_0000_0000;
array[6203] <= 16'b0000_0000_0000_0000;
array[6204] <= 16'b0000_0000_0000_0000;
array[6205] <= 16'b0000_0000_0000_0000;
array[6206] <= 16'b0000_0000_0000_0000;
array[6207] <= 16'b0000_0000_0000_0000;
array[6208] <= 16'b0000_0000_0000_0000;
array[6209] <= 16'b0000_0000_0000_0000;
array[6210] <= 16'b0000_0000_0000_0000;
array[6211] <= 16'b0000_0000_0000_0000;
array[6212] <= 16'b0000_0000_0000_0000;
array[6213] <= 16'b0000_0000_0000_0000;
array[6214] <= 16'b0000_0000_0000_0000;
array[6215] <= 16'b0000_0000_0000_0000;
array[6216] <= 16'b0000_0000_0000_0000;
array[6217] <= 16'b0000_0000_0000_0000;
array[6218] <= 16'b0000_0000_0000_0000;
array[6219] <= 16'b0000_0000_0000_0000;
array[6220] <= 16'b0000_0000_0000_0000;
array[6221] <= 16'b0000_0000_0000_0000;
array[6222] <= 16'b0000_0000_0000_0000;
array[6223] <= 16'b0000_0000_0000_0000;
array[6224] <= 16'b0000_0000_0000_0000;
array[6225] <= 16'b0000_0000_0000_0000;
array[6226] <= 16'b0000_0000_0000_0000;
array[6227] <= 16'b0000_0000_0000_0000;
array[6228] <= 16'b0000_0000_0000_0000;
array[6229] <= 16'b0000_0000_0000_0000;
array[6230] <= 16'b0000_0000_0000_0000;
array[6231] <= 16'b0000_0000_0000_0000;
array[6232] <= 16'b0000_0000_0000_0000;
array[6233] <= 16'b0000_0000_0000_0000;
array[6234] <= 16'b0000_0000_0000_0000;
array[6235] <= 16'b0000_0000_0000_0000;
array[6236] <= 16'b0000_0000_0000_0000;
array[6237] <= 16'b0000_0000_0000_0000;
array[6238] <= 16'b0000_0000_0000_0000;
array[6239] <= 16'b0000_0000_0000_0000;
array[6240] <= 16'b0000_0000_0000_0000;
array[6241] <= 16'b0000_0000_0000_0000;
array[6242] <= 16'b0000_0000_0000_0000;
array[6243] <= 16'b0000_0000_0000_0000;
array[6244] <= 16'b0000_0000_0000_0000;
array[6245] <= 16'b0000_0000_0000_0000;
array[6246] <= 16'b0000_0000_0000_0000;
array[6247] <= 16'b0000_0000_0000_0000;
array[6248] <= 16'b0000_0000_0000_0000;
array[6249] <= 16'b0000_0000_0000_0000;
array[6250] <= 16'b0000_0000_0000_0000;
array[6251] <= 16'b0000_0000_0000_0000;
array[6252] <= 16'b0000_0000_0000_0000;
array[6253] <= 16'b0000_0000_0000_0000;
array[6254] <= 16'b0000_0000_0000_0000;
array[6255] <= 16'b0000_0000_0000_0000;
array[6256] <= 16'b0000_0000_0000_0000;
array[6257] <= 16'b0000_0000_0000_0000;
array[6258] <= 16'b0000_0000_0000_0000;
array[6259] <= 16'b0000_0000_0000_0000;
array[6260] <= 16'b0000_0000_0000_0000;
array[6261] <= 16'b0000_0000_0000_0000;
array[6262] <= 16'b0000_0000_0000_0000;
array[6263] <= 16'b0000_0000_0000_0000;
array[6264] <= 16'b0000_0000_0000_0000;
array[6265] <= 16'b0000_0000_0000_0000;
array[6266] <= 16'b0000_0000_0000_0000;
array[6267] <= 16'b0000_0000_0000_0000;
array[6268] <= 16'b0000_0000_0000_0000;
array[6269] <= 16'b0000_0000_0000_0000;
array[6270] <= 16'b0000_0000_0000_0000;
array[6271] <= 16'b0000_0000_0000_0000;
array[6272] <= 16'b0000_0000_0000_0000;
array[6273] <= 16'b0000_0000_0000_0000;
array[6274] <= 16'b0000_0000_0000_0000;
array[6275] <= 16'b0000_0000_0000_0000;
array[6276] <= 16'b0000_0000_0000_0000;
array[6277] <= 16'b0000_0000_0000_0000;
array[6278] <= 16'b0000_0000_0000_0000;
array[6279] <= 16'b0000_0000_0000_0000;
array[6280] <= 16'b0000_0000_0000_0000;
array[6281] <= 16'b0000_0000_0000_0000;
array[6282] <= 16'b0000_0000_0000_0000;
array[6283] <= 16'b0000_0000_0000_0000;
array[6284] <= 16'b0000_0000_0000_0000;
array[6285] <= 16'b0000_0000_0000_0000;
array[6286] <= 16'b0000_0000_0000_0000;
array[6287] <= 16'b0000_0000_0000_0000;
array[6288] <= 16'b0000_0000_0000_0000;
array[6289] <= 16'b0000_0000_0000_0000;
array[6290] <= 16'b0000_0000_0000_0000;
array[6291] <= 16'b0000_0000_0000_0000;
array[6292] <= 16'b0000_0000_0000_0000;
array[6293] <= 16'b0000_0000_0000_0000;
array[6294] <= 16'b0000_0000_0000_0000;
array[6295] <= 16'b0000_0000_0000_0000;
array[6296] <= 16'b0000_0000_0000_0000;
array[6297] <= 16'b0000_0000_0000_0000;
array[6298] <= 16'b0000_0000_0000_0000;
array[6299] <= 16'b0000_0000_0000_0000;
array[6300] <= 16'b0000_0000_0000_0000;
array[6301] <= 16'b0000_0000_0000_0000;
array[6302] <= 16'b0000_0000_0000_0000;
array[6303] <= 16'b0000_0000_0000_0000;
array[6304] <= 16'b0000_0000_0000_0000;
array[6305] <= 16'b0000_0000_0000_0000;
array[6306] <= 16'b0000_0000_0000_0000;
array[6307] <= 16'b0000_0000_0000_0000;
array[6308] <= 16'b0000_0000_0000_0000;
array[6309] <= 16'b0000_0000_0000_0000;
array[6310] <= 16'b0000_0000_0000_0000;
array[6311] <= 16'b0000_0000_0000_0000;
array[6312] <= 16'b0000_0000_0000_0000;
array[6313] <= 16'b0000_0000_0000_0000;
array[6314] <= 16'b0000_0000_0000_0000;
array[6315] <= 16'b0000_0000_0000_0000;
array[6316] <= 16'b0000_0000_0000_0000;
array[6317] <= 16'b0000_0000_0000_0000;
array[6318] <= 16'b0000_0000_0000_0000;
array[6319] <= 16'b0000_0000_0000_0000;
array[6320] <= 16'b0000_0000_0000_0000;
array[6321] <= 16'b0000_0000_0000_0000;
array[6322] <= 16'b0000_0000_0000_0000;
array[6323] <= 16'b0000_0000_0000_0000;
array[6324] <= 16'b0000_0000_0000_0000;
array[6325] <= 16'b0000_0000_0000_0000;
array[6326] <= 16'b0000_0000_0000_0000;
array[6327] <= 16'b0000_0000_0000_0000;
array[6328] <= 16'b0000_0000_0000_0000;
array[6329] <= 16'b0000_0000_0000_0000;
array[6330] <= 16'b0000_0000_0000_0000;
array[6331] <= 16'b0000_0000_0000_0000;
array[6332] <= 16'b0000_0000_0000_0000;
array[6333] <= 16'b0000_0000_0000_0000;
array[6334] <= 16'b0000_0000_0000_0000;
array[6335] <= 16'b0000_0000_0000_0000;
array[6336] <= 16'b0000_0000_0000_0000;
array[6337] <= 16'b0000_0000_0000_0000;
array[6338] <= 16'b0000_0000_0000_0000;
array[6339] <= 16'b0000_0000_0000_0000;
array[6340] <= 16'b0000_0000_0000_0000;
array[6341] <= 16'b0000_0000_0000_0000;
array[6342] <= 16'b0000_0000_0000_0000;
array[6343] <= 16'b0000_0000_0000_0000;
array[6344] <= 16'b0000_0000_0000_0000;
array[6345] <= 16'b0000_0000_0000_0000;
array[6346] <= 16'b0000_0000_0000_0000;
array[6347] <= 16'b0000_0000_0000_0000;
array[6348] <= 16'b0000_0000_0000_0000;
array[6349] <= 16'b0000_0000_0000_0000;
array[6350] <= 16'b0000_0000_0000_0000;
array[6351] <= 16'b0000_0000_0000_0000;
array[6352] <= 16'b0000_0000_0000_0000;
array[6353] <= 16'b0000_0000_0000_0000;
array[6354] <= 16'b0000_0000_0000_0000;
array[6355] <= 16'b0000_0000_0000_0000;
array[6356] <= 16'b0000_0000_0000_0000;
array[6357] <= 16'b0000_0000_0000_0000;
array[6358] <= 16'b0000_0000_0000_0000;
array[6359] <= 16'b0000_0000_0000_0000;
array[6360] <= 16'b0000_0000_0000_0000;
array[6361] <= 16'b0000_0000_0000_0000;
array[6362] <= 16'b0000_0000_0000_0000;
array[6363] <= 16'b0000_0000_0000_0000;
array[6364] <= 16'b0000_0000_0000_0000;
array[6365] <= 16'b0000_0000_0000_0000;
array[6366] <= 16'b0000_0000_0000_0000;
array[6367] <= 16'b0000_0000_0000_0000;
array[6368] <= 16'b0000_0000_0000_0000;
array[6369] <= 16'b0000_0000_0000_0000;
array[6370] <= 16'b0000_0000_0000_0000;
array[6371] <= 16'b0000_0000_0000_0000;
array[6372] <= 16'b0000_0000_0000_0000;
array[6373] <= 16'b0000_0000_0000_0000;
array[6374] <= 16'b0000_0000_0000_0000;
array[6375] <= 16'b0000_0000_0000_0000;
array[6376] <= 16'b0000_0000_0000_0000;
array[6377] <= 16'b0000_0000_0000_0000;
array[6378] <= 16'b0000_0000_0000_0000;
array[6379] <= 16'b0000_0000_0000_0000;
array[6380] <= 16'b0000_0000_0000_0000;
array[6381] <= 16'b0000_0000_0000_0000;
array[6382] <= 16'b0000_0000_0000_0000;
array[6383] <= 16'b0000_0000_0000_0000;
array[6384] <= 16'b0000_0000_0000_0000;
array[6385] <= 16'b0000_0000_0000_0000;
array[6386] <= 16'b0000_0000_0000_0000;
array[6387] <= 16'b0000_0000_0000_0000;
array[6388] <= 16'b0000_0000_0000_0000;
array[6389] <= 16'b0000_0000_0000_0000;
array[6390] <= 16'b0000_0000_0000_0000;
array[6391] <= 16'b0000_0000_0000_0000;
array[6392] <= 16'b0000_0000_0000_0000;
array[6393] <= 16'b0000_0000_0000_0000;
array[6394] <= 16'b0000_0000_0000_0000;
array[6395] <= 16'b0000_0000_0000_0000;
array[6396] <= 16'b0000_0000_0000_0000;
array[6397] <= 16'b0000_0000_0000_0000;
array[6398] <= 16'b0000_0000_0000_0000;
array[6399] <= 16'b0000_0000_0000_0000;
array[6400] <= 16'b0000_0000_0000_0000;
array[6401] <= 16'b0000_0000_0000_0000;
array[6402] <= 16'b0000_0000_0000_0000;
array[6403] <= 16'b0000_0000_0000_0000;
array[6404] <= 16'b0000_0000_0000_0000;
array[6405] <= 16'b0000_0000_0000_0000;
array[6406] <= 16'b0000_0000_0000_0000;
array[6407] <= 16'b0000_0000_0000_0000;
array[6408] <= 16'b0000_0000_0000_0000;
array[6409] <= 16'b0000_0000_0000_0000;
array[6410] <= 16'b0000_0000_0000_0000;
array[6411] <= 16'b0000_0000_0000_0000;
array[6412] <= 16'b0000_0000_0000_0000;
array[6413] <= 16'b0000_0000_0000_0000;
array[6414] <= 16'b0000_0000_0000_0000;
array[6415] <= 16'b0000_0000_0000_0000;
array[6416] <= 16'b0000_0000_0000_0000;
array[6417] <= 16'b0000_0000_0000_0000;
array[6418] <= 16'b0000_0000_0000_0000;
array[6419] <= 16'b0000_0000_0000_0000;
array[6420] <= 16'b0000_0000_0000_0000;
array[6421] <= 16'b0000_0000_0000_0000;
array[6422] <= 16'b0000_0000_0000_0000;
array[6423] <= 16'b0000_0000_0000_0000;
array[6424] <= 16'b0000_0000_0000_0000;
array[6425] <= 16'b0000_0000_0000_0000;
array[6426] <= 16'b0000_0000_0000_0000;
array[6427] <= 16'b0000_0000_0000_0000;
array[6428] <= 16'b0000_0000_0000_0000;
array[6429] <= 16'b0000_0000_0000_0000;
array[6430] <= 16'b0000_0000_0000_0000;
array[6431] <= 16'b0000_0000_0000_0000;
array[6432] <= 16'b0000_0000_0000_0000;
array[6433] <= 16'b0000_0000_0000_0000;
array[6434] <= 16'b0000_0000_0000_0000;
array[6435] <= 16'b0000_0000_0000_0000;
array[6436] <= 16'b0000_0000_0000_0000;
array[6437] <= 16'b0000_0000_0000_0000;
array[6438] <= 16'b0000_0000_0000_0000;
array[6439] <= 16'b0000_0000_0000_0000;
array[6440] <= 16'b0000_0000_0000_0000;
array[6441] <= 16'b0000_0000_0000_0000;
array[6442] <= 16'b0000_0000_0000_0000;
array[6443] <= 16'b0000_0000_0000_0000;
array[6444] <= 16'b0000_0000_0000_0000;
array[6445] <= 16'b0000_0000_0000_0000;
array[6446] <= 16'b0000_0000_0000_0000;
array[6447] <= 16'b0000_0000_0000_0000;
array[6448] <= 16'b0000_0000_0000_0000;
array[6449] <= 16'b0000_0000_0000_0000;
array[6450] <= 16'b0000_0000_0000_0000;
array[6451] <= 16'b0000_0000_0000_0000;
array[6452] <= 16'b0000_0000_0000_0000;
array[6453] <= 16'b0000_0000_0000_0000;
array[6454] <= 16'b0000_0000_0000_0000;
array[6455] <= 16'b0000_0000_0000_0000;
array[6456] <= 16'b0000_0000_0000_0000;
array[6457] <= 16'b0000_0000_0000_0000;
array[6458] <= 16'b0000_0000_0000_0000;
array[6459] <= 16'b0000_0000_0000_0000;
array[6460] <= 16'b0000_0000_0000_0000;
array[6461] <= 16'b0000_0000_0000_0000;
array[6462] <= 16'b0000_0000_0000_0000;
array[6463] <= 16'b0000_0000_0000_0000;
array[6464] <= 16'b0000_0000_0000_0000;
array[6465] <= 16'b0000_0000_0000_0000;
array[6466] <= 16'b0000_0000_0000_0000;
array[6467] <= 16'b0000_0000_0000_0000;
array[6468] <= 16'b0000_0000_0000_0000;
array[6469] <= 16'b0000_0000_0000_0000;
array[6470] <= 16'b0000_0000_0000_0000;
array[6471] <= 16'b0000_0000_0000_0000;
array[6472] <= 16'b0000_0000_0000_0000;
array[6473] <= 16'b0000_0000_0000_0000;
array[6474] <= 16'b0000_0000_0000_0000;
array[6475] <= 16'b0000_0000_0000_0000;
array[6476] <= 16'b0000_0000_0000_0000;
array[6477] <= 16'b0000_0000_0000_0000;
array[6478] <= 16'b0000_0000_0000_0000;
array[6479] <= 16'b0000_0000_0000_0000;
array[6480] <= 16'b0000_0000_0000_0000;
array[6481] <= 16'b0000_0000_0000_0000;
array[6482] <= 16'b0000_0000_0000_0000;
array[6483] <= 16'b0000_0000_0000_0000;
array[6484] <= 16'b0000_0000_0000_0000;
array[6485] <= 16'b0000_0000_0000_0000;
array[6486] <= 16'b0000_0000_0000_0000;
array[6487] <= 16'b0000_0000_0000_0000;
array[6488] <= 16'b0000_0000_0000_0000;
array[6489] <= 16'b0000_0000_0000_0000;
array[6490] <= 16'b0000_0000_0000_0000;
array[6491] <= 16'b0000_0000_0000_0000;
array[6492] <= 16'b0000_0000_0000_0000;
array[6493] <= 16'b0000_0000_0000_0000;
array[6494] <= 16'b0000_0000_0000_0000;
array[6495] <= 16'b0000_0000_0000_0000;
array[6496] <= 16'b0000_0000_0000_0000;
array[6497] <= 16'b0000_0000_0000_0000;
array[6498] <= 16'b0000_0000_0000_0000;
array[6499] <= 16'b0000_0000_0000_0000;
array[6500] <= 16'b0000_0000_0000_0000;
array[6501] <= 16'b0000_0000_0000_0000;
array[6502] <= 16'b0000_0000_0000_0000;
array[6503] <= 16'b0000_0000_0000_0000;
array[6504] <= 16'b0000_0000_0000_0000;
array[6505] <= 16'b0000_0000_0000_0000;
array[6506] <= 16'b0000_0000_0000_0000;
array[6507] <= 16'b0000_0000_0000_0000;
array[6508] <= 16'b0000_0000_0000_0000;
array[6509] <= 16'b0000_0000_0000_0000;
array[6510] <= 16'b0000_0000_0000_0000;
array[6511] <= 16'b0000_0000_0000_0000;
array[6512] <= 16'b0000_0000_0000_0000;
array[6513] <= 16'b0000_0000_0000_0000;
array[6514] <= 16'b0000_0000_0000_0000;
array[6515] <= 16'b0000_0000_0000_0000;
array[6516] <= 16'b0000_0000_0000_0000;
array[6517] <= 16'b0000_0000_0000_0000;
array[6518] <= 16'b0000_0000_0000_0000;
array[6519] <= 16'b0000_0000_0000_0000;
array[6520] <= 16'b0000_0000_0000_0000;
array[6521] <= 16'b0000_0000_0000_0000;
array[6522] <= 16'b0000_0000_0000_0000;
array[6523] <= 16'b0000_0000_0000_0000;
array[6524] <= 16'b0000_0000_0000_0000;
array[6525] <= 16'b0000_0000_0000_0000;
array[6526] <= 16'b0000_0000_0000_0000;
array[6527] <= 16'b0000_0000_0000_0000;
array[6528] <= 16'b0000_0000_0000_0000;
array[6529] <= 16'b0000_0000_0000_0000;
array[6530] <= 16'b0000_0000_0000_0000;
array[6531] <= 16'b0000_0000_0000_0000;
array[6532] <= 16'b0000_0000_0000_0000;
array[6533] <= 16'b0000_0000_0000_0000;
array[6534] <= 16'b0000_0000_0000_0000;
array[6535] <= 16'b0000_0000_0000_0000;
array[6536] <= 16'b0000_0000_0000_0000;
array[6537] <= 16'b0000_0000_0000_0000;
array[6538] <= 16'b0000_0000_0000_0000;
array[6539] <= 16'b0000_0000_0000_0000;
array[6540] <= 16'b0000_0000_0000_0000;
array[6541] <= 16'b0000_0000_0000_0000;
array[6542] <= 16'b0000_0000_0000_0000;
array[6543] <= 16'b0000_0000_0000_0000;
array[6544] <= 16'b0000_0000_0000_0000;
array[6545] <= 16'b0000_0000_0000_0000;
array[6546] <= 16'b0000_0000_0000_0000;
array[6547] <= 16'b0000_0000_0000_0000;
array[6548] <= 16'b0000_0000_0000_0000;
array[6549] <= 16'b0000_0000_0000_0000;
array[6550] <= 16'b0000_0000_0000_0000;
array[6551] <= 16'b0000_0000_0000_0000;
array[6552] <= 16'b0000_0000_0000_0000;
array[6553] <= 16'b0000_0000_0000_0000;
array[6554] <= 16'b0000_0000_0000_0000;
array[6555] <= 16'b0000_0000_0000_0000;
array[6556] <= 16'b0000_0000_0000_0000;
array[6557] <= 16'b0000_0000_0000_0000;
array[6558] <= 16'b0000_0000_0000_0000;
array[6559] <= 16'b0000_0000_0000_0000;
array[6560] <= 16'b0000_0000_0000_0000;
array[6561] <= 16'b0000_0000_0000_0000;
array[6562] <= 16'b0000_0000_0000_0000;
array[6563] <= 16'b0000_0000_0000_0000;
array[6564] <= 16'b0000_0000_0000_0000;
array[6565] <= 16'b0000_0000_0000_0000;
array[6566] <= 16'b0000_0000_0000_0000;
array[6567] <= 16'b0000_0000_0000_0000;
array[6568] <= 16'b0000_0000_0000_0000;
array[6569] <= 16'b0000_0000_0000_0000;
array[6570] <= 16'b0000_0000_0000_0000;
array[6571] <= 16'b0000_0000_0000_0000;
array[6572] <= 16'b0000_0000_0000_0000;
array[6573] <= 16'b0000_0000_0000_0000;
array[6574] <= 16'b0000_0000_0000_0000;
array[6575] <= 16'b0000_0000_0000_0000;
array[6576] <= 16'b0000_0000_0000_0000;
array[6577] <= 16'b0000_0000_0000_0000;
array[6578] <= 16'b0000_0000_0000_0000;
array[6579] <= 16'b0000_0000_0000_0000;
array[6580] <= 16'b0000_0000_0000_0000;
array[6581] <= 16'b0000_0000_0000_0000;
array[6582] <= 16'b0000_0000_0000_0000;
array[6583] <= 16'b0000_0000_0000_0000;
array[6584] <= 16'b0000_0000_0000_0000;
array[6585] <= 16'b0000_0000_0000_0000;
array[6586] <= 16'b0000_0000_0000_0000;
array[6587] <= 16'b0000_0000_0000_0000;
array[6588] <= 16'b0000_0000_0000_0000;
array[6589] <= 16'b0000_0000_0000_0000;
array[6590] <= 16'b0000_0000_0000_0000;
array[6591] <= 16'b0000_0000_0000_0000;
array[6592] <= 16'b0000_0000_0000_0000;
array[6593] <= 16'b0000_0000_0000_0000;
array[6594] <= 16'b0000_0000_0000_0000;
array[6595] <= 16'b0000_0000_0000_0000;
array[6596] <= 16'b0000_0000_0000_0000;
array[6597] <= 16'b0000_0000_0000_0000;
array[6598] <= 16'b0000_0000_0000_0000;
array[6599] <= 16'b0000_0000_0000_0000;
array[6600] <= 16'b0000_0000_0000_0000;
array[6601] <= 16'b0000_0000_0000_0000;
array[6602] <= 16'b0000_0000_0000_0000;
array[6603] <= 16'b0000_0000_0000_0000;
array[6604] <= 16'b0000_0000_0000_0000;
array[6605] <= 16'b0000_0000_0000_0000;
array[6606] <= 16'b0000_0000_0000_0000;
array[6607] <= 16'b0000_0000_0000_0000;
array[6608] <= 16'b0000_0000_0000_0000;
array[6609] <= 16'b0000_0000_0000_0000;
array[6610] <= 16'b0000_0000_0000_0000;
array[6611] <= 16'b0000_0000_0000_0000;
array[6612] <= 16'b0000_0000_0000_0000;
array[6613] <= 16'b0000_0000_0000_0000;
array[6614] <= 16'b0000_0000_0000_0000;
array[6615] <= 16'b0000_0000_0000_0000;
array[6616] <= 16'b0000_0000_0000_0000;
array[6617] <= 16'b0000_0000_0000_0000;
array[6618] <= 16'b0000_0000_0000_0000;
array[6619] <= 16'b0000_0000_0000_0000;
array[6620] <= 16'b0000_0000_0000_0000;
array[6621] <= 16'b0000_0000_0000_0000;
array[6622] <= 16'b0000_0000_0000_0000;
array[6623] <= 16'b0000_0000_0000_0000;
array[6624] <= 16'b0000_0000_0000_0000;
array[6625] <= 16'b0000_0000_0000_0000;
array[6626] <= 16'b0000_0000_0000_0000;
array[6627] <= 16'b0000_0000_0000_0000;
array[6628] <= 16'b0000_0000_0000_0000;
array[6629] <= 16'b0000_0000_0000_0000;
array[6630] <= 16'b0000_0000_0000_0000;
array[6631] <= 16'b0000_0000_0000_0000;
array[6632] <= 16'b0000_0000_0000_0000;
array[6633] <= 16'b0000_0000_0000_0000;
array[6634] <= 16'b0000_0000_0000_0000;
array[6635] <= 16'b0000_0000_0000_0000;
array[6636] <= 16'b0000_0000_0000_0000;
array[6637] <= 16'b0000_0000_0000_0000;
array[6638] <= 16'b0000_0000_0000_0000;
array[6639] <= 16'b0000_0000_0000_0000;
array[6640] <= 16'b0000_0000_0000_0000;
array[6641] <= 16'b0000_0000_0000_0000;
array[6642] <= 16'b0000_0000_0000_0000;
array[6643] <= 16'b0000_0000_0000_0000;
array[6644] <= 16'b0000_0000_0000_0000;
array[6645] <= 16'b0000_0000_0000_0000;
array[6646] <= 16'b0000_0000_0000_0000;
array[6647] <= 16'b0000_0000_0000_0000;
array[6648] <= 16'b0000_0000_0000_0000;
array[6649] <= 16'b0000_0000_0000_0000;
array[6650] <= 16'b0000_0000_0000_0000;
array[6651] <= 16'b0000_0000_0000_0000;
array[6652] <= 16'b0000_0000_0000_0000;
array[6653] <= 16'b0000_0000_0000_0000;
array[6654] <= 16'b0000_0000_0000_0000;
array[6655] <= 16'b0000_0000_0000_0000;
array[6656] <= 16'b0000_0000_0000_0000;
array[6657] <= 16'b0000_0000_0000_0000;
array[6658] <= 16'b0000_0000_0000_0000;
array[6659] <= 16'b0000_0000_0000_0000;
array[6660] <= 16'b0000_0000_0000_0000;
array[6661] <= 16'b0000_0000_0000_0000;
array[6662] <= 16'b0000_0000_0000_0000;
array[6663] <= 16'b0000_0000_0000_0000;
array[6664] <= 16'b0000_0000_0000_0000;
array[6665] <= 16'b0000_0000_0000_0000;
array[6666] <= 16'b0000_0000_0000_0000;
array[6667] <= 16'b0000_0000_0000_0000;
array[6668] <= 16'b0000_0000_0000_0000;
array[6669] <= 16'b0000_0000_0000_0000;
array[6670] <= 16'b0000_0000_0000_0000;
array[6671] <= 16'b0000_0000_0000_0000;
array[6672] <= 16'b0000_0000_0000_0000;
array[6673] <= 16'b0000_0000_0000_0000;
array[6674] <= 16'b0000_0000_0000_0000;
array[6675] <= 16'b0000_0000_0000_0000;
array[6676] <= 16'b0000_0000_0000_0000;
array[6677] <= 16'b0000_0000_0000_0000;
array[6678] <= 16'b0000_0000_0000_0000;
array[6679] <= 16'b0000_0000_0000_0000;
array[6680] <= 16'b0000_0000_0000_0000;
array[6681] <= 16'b0000_0000_0000_0000;
array[6682] <= 16'b0000_0000_0000_0000;
array[6683] <= 16'b0000_0000_0000_0000;
array[6684] <= 16'b0000_0000_0000_0000;
array[6685] <= 16'b0000_0000_0000_0000;
array[6686] <= 16'b0000_0000_0000_0000;
array[6687] <= 16'b0000_0000_0000_0000;
array[6688] <= 16'b0000_0000_0000_0000;
array[6689] <= 16'b0000_0000_0000_0000;
array[6690] <= 16'b0000_0000_0000_0000;
array[6691] <= 16'b0000_0000_0000_0000;
array[6692] <= 16'b0000_0000_0000_0000;
array[6693] <= 16'b0000_0000_0000_0000;
array[6694] <= 16'b0000_0000_0000_0000;
array[6695] <= 16'b0000_0000_0000_0000;
array[6696] <= 16'b0000_0000_0000_0000;
array[6697] <= 16'b0000_0000_0000_0000;
array[6698] <= 16'b0000_0000_0000_0000;
array[6699] <= 16'b0000_0000_0000_0000;
array[6700] <= 16'b0000_0000_0000_0000;
array[6701] <= 16'b0000_0000_0000_0000;
array[6702] <= 16'b0000_0000_0000_0000;
array[6703] <= 16'b0000_0000_0000_0000;
array[6704] <= 16'b0000_0000_0000_0000;
array[6705] <= 16'b0000_0000_0000_0000;
array[6706] <= 16'b0000_0000_0000_0000;
array[6707] <= 16'b0000_0000_0000_0000;
array[6708] <= 16'b0000_0000_0000_0000;
array[6709] <= 16'b0000_0000_0000_0000;
array[6710] <= 16'b0000_0000_0000_0000;
array[6711] <= 16'b0000_0000_0000_0000;
array[6712] <= 16'b0000_0000_0000_0000;
array[6713] <= 16'b0000_0000_0000_0000;
array[6714] <= 16'b0000_0000_0000_0000;
array[6715] <= 16'b0000_0000_0000_0000;
array[6716] <= 16'b0000_0000_0000_0000;
array[6717] <= 16'b0000_0000_0000_0000;
array[6718] <= 16'b0000_0000_0000_0000;
array[6719] <= 16'b0000_0000_0000_0000;
array[6720] <= 16'b0000_0000_0000_0000;
array[6721] <= 16'b0000_0000_0000_0000;
array[6722] <= 16'b0000_0000_0000_0000;
array[6723] <= 16'b0000_0000_0000_0000;
array[6724] <= 16'b0000_0000_0000_0000;
array[6725] <= 16'b0000_0000_0000_0000;
array[6726] <= 16'b0000_0000_0000_0000;
array[6727] <= 16'b0000_0000_0000_0000;
array[6728] <= 16'b0000_0000_0000_0000;
array[6729] <= 16'b0000_0000_0000_0000;
array[6730] <= 16'b0000_0000_0000_0000;
array[6731] <= 16'b0000_0000_0000_0000;
array[6732] <= 16'b0000_0000_0000_0000;
array[6733] <= 16'b0000_0000_0000_0000;
array[6734] <= 16'b0000_0000_0000_0000;
array[6735] <= 16'b0000_0000_0000_0000;
array[6736] <= 16'b0000_0000_0000_0000;
array[6737] <= 16'b0000_0000_0000_0000;
array[6738] <= 16'b0000_0000_0000_0000;
array[6739] <= 16'b0000_0000_0000_0000;
array[6740] <= 16'b0000_0000_0000_0000;
array[6741] <= 16'b0000_0000_0000_0000;
array[6742] <= 16'b0000_0000_0000_0000;
array[6743] <= 16'b0000_0000_0000_0000;
array[6744] <= 16'b0000_0000_0000_0000;
array[6745] <= 16'b0000_0000_0000_0000;
array[6746] <= 16'b0000_0000_0000_0000;
array[6747] <= 16'b0000_0000_0000_0000;
array[6748] <= 16'b0000_0000_0000_0000;
array[6749] <= 16'b0000_0000_0000_0000;
array[6750] <= 16'b0000_0000_0000_0000;
array[6751] <= 16'b0000_0000_0000_0000;
array[6752] <= 16'b0000_0000_0000_0000;
array[6753] <= 16'b0000_0000_0000_0000;
array[6754] <= 16'b0000_0000_0000_0000;
array[6755] <= 16'b0000_0000_0000_0000;
array[6756] <= 16'b0000_0000_0000_0000;
array[6757] <= 16'b0000_0000_0000_0000;
array[6758] <= 16'b0000_0000_0000_0000;
array[6759] <= 16'b0000_0000_0000_0000;
array[6760] <= 16'b0000_0000_0000_0000;
array[6761] <= 16'b0000_0000_0000_0000;
array[6762] <= 16'b0000_0000_0000_0000;
array[6763] <= 16'b0000_0000_0000_0000;
array[6764] <= 16'b0000_0000_0000_0000;
array[6765] <= 16'b0000_0000_0000_0000;
array[6766] <= 16'b0000_0000_0000_0000;
array[6767] <= 16'b0000_0000_0000_0000;
array[6768] <= 16'b0000_0000_0000_0000;
array[6769] <= 16'b0000_0000_0000_0000;
array[6770] <= 16'b0000_0000_0000_0000;
array[6771] <= 16'b0000_0000_0000_0000;
array[6772] <= 16'b0000_0000_0000_0000;
array[6773] <= 16'b0000_0000_0000_0000;
array[6774] <= 16'b0000_0000_0000_0000;
array[6775] <= 16'b0000_0000_0000_0000;
array[6776] <= 16'b0000_0000_0000_0000;
array[6777] <= 16'b0000_0000_0000_0000;
array[6778] <= 16'b0000_0000_0000_0000;
array[6779] <= 16'b0000_0000_0000_0000;
array[6780] <= 16'b0000_0000_0000_0000;
array[6781] <= 16'b0000_0000_0000_0000;
array[6782] <= 16'b0000_0000_0000_0000;
array[6783] <= 16'b0000_0000_0000_0000;
array[6784] <= 16'b0000_0000_0000_0000;
array[6785] <= 16'b0000_0000_0000_0000;
array[6786] <= 16'b0000_0000_0000_0000;
array[6787] <= 16'b0000_0000_0000_0000;
array[6788] <= 16'b0000_0000_0000_0000;
array[6789] <= 16'b0000_0000_0000_0000;
array[6790] <= 16'b0000_0000_0000_0000;
array[6791] <= 16'b0000_0000_0000_0000;
array[6792] <= 16'b0000_0000_0000_0000;
array[6793] <= 16'b0000_0000_0000_0000;
array[6794] <= 16'b0000_0000_0000_0000;
array[6795] <= 16'b0000_0000_0000_0000;
array[6796] <= 16'b0000_0000_0000_0000;
array[6797] <= 16'b0000_0000_0000_0000;
array[6798] <= 16'b0000_0000_0000_0000;
array[6799] <= 16'b0000_0000_0000_0000;
array[6800] <= 16'b0000_0000_0000_0000;
array[6801] <= 16'b0000_0000_0000_0000;
array[6802] <= 16'b0000_0000_0000_0000;
array[6803] <= 16'b0000_0000_0000_0000;
array[6804] <= 16'b0000_0000_0000_0000;
array[6805] <= 16'b0000_0000_0000_0000;
array[6806] <= 16'b0000_0000_0000_0000;
array[6807] <= 16'b0000_0000_0000_0000;
array[6808] <= 16'b0000_0000_0000_0000;
array[6809] <= 16'b0000_0000_0000_0000;
array[6810] <= 16'b0000_0000_0000_0000;
array[6811] <= 16'b0000_0000_0000_0000;
array[6812] <= 16'b0000_0000_0000_0000;
array[6813] <= 16'b0000_0000_0000_0000;
array[6814] <= 16'b0000_0000_0000_0000;
array[6815] <= 16'b0000_0000_0000_0000;
array[6816] <= 16'b0000_0000_0000_0000;
array[6817] <= 16'b0000_0000_0000_0000;
array[6818] <= 16'b0000_0000_0000_0000;
array[6819] <= 16'b0000_0000_0000_0000;
array[6820] <= 16'b0000_0000_0000_0000;
array[6821] <= 16'b0000_0000_0000_0000;
array[6822] <= 16'b0000_0000_0000_0000;
array[6823] <= 16'b0000_0000_0000_0000;
array[6824] <= 16'b0000_0000_0000_0000;
array[6825] <= 16'b0000_0000_0000_0000;
array[6826] <= 16'b0000_0000_0000_0000;
array[6827] <= 16'b0000_0000_0000_0000;
array[6828] <= 16'b0000_0000_0000_0000;
array[6829] <= 16'b0000_0000_0000_0000;
array[6830] <= 16'b0000_0000_0000_0000;
array[6831] <= 16'b0000_0000_0000_0000;
array[6832] <= 16'b0000_0000_0000_0000;
array[6833] <= 16'b0000_0000_0000_0000;
array[6834] <= 16'b0000_0000_0000_0000;
array[6835] <= 16'b0000_0000_0000_0000;
array[6836] <= 16'b0000_0000_0000_0000;
array[6837] <= 16'b0000_0000_0000_0000;
array[6838] <= 16'b0000_0000_0000_0000;
array[6839] <= 16'b0000_0000_0000_0000;
array[6840] <= 16'b0000_0000_0000_0000;
array[6841] <= 16'b0000_0000_0000_0000;
array[6842] <= 16'b0000_0000_0000_0000;
array[6843] <= 16'b0000_0000_0000_0000;
array[6844] <= 16'b0000_0000_0000_0000;
array[6845] <= 16'b0000_0000_0000_0000;
array[6846] <= 16'b0000_0000_0000_0000;
array[6847] <= 16'b0000_0000_0000_0000;
array[6848] <= 16'b0000_0000_0000_0000;
array[6849] <= 16'b0000_0000_0000_0000;
array[6850] <= 16'b0000_0000_0000_0000;
array[6851] <= 16'b0000_0000_0000_0000;
array[6852] <= 16'b0000_0000_0000_0000;
array[6853] <= 16'b0000_0000_0000_0000;
array[6854] <= 16'b0000_0000_0000_0000;
array[6855] <= 16'b0000_0000_0000_0000;
array[6856] <= 16'b0000_0000_0000_0000;
array[6857] <= 16'b0000_0000_0000_0000;
array[6858] <= 16'b0000_0000_0000_0000;
array[6859] <= 16'b0000_0000_0000_0000;
array[6860] <= 16'b0000_0000_0000_0000;
array[6861] <= 16'b0000_0000_0000_0000;
array[6862] <= 16'b0000_0000_0000_0000;
array[6863] <= 16'b0000_0000_0000_0000;
array[6864] <= 16'b0000_0000_0000_0000;
array[6865] <= 16'b0000_0000_0000_0000;
array[6866] <= 16'b0000_0000_0000_0000;
array[6867] <= 16'b0000_0000_0000_0000;
array[6868] <= 16'b0000_0000_0000_0000;
array[6869] <= 16'b0000_0000_0000_0000;
array[6870] <= 16'b0000_0000_0000_0000;
array[6871] <= 16'b0000_0000_0000_0000;
array[6872] <= 16'b0000_0000_0000_0000;
array[6873] <= 16'b0000_0000_0000_0000;
array[6874] <= 16'b0000_0000_0000_0000;
array[6875] <= 16'b0000_0000_0000_0000;
array[6876] <= 16'b0000_0000_0000_0000;
array[6877] <= 16'b0000_0000_0000_0000;
array[6878] <= 16'b0000_0000_0000_0000;
array[6879] <= 16'b0000_0000_0000_0000;
array[6880] <= 16'b0000_0000_0000_0000;
array[6881] <= 16'b0000_0000_0000_0000;
array[6882] <= 16'b0000_0000_0000_0000;
array[6883] <= 16'b0000_0000_0000_0000;
array[6884] <= 16'b0000_0000_0000_0000;
array[6885] <= 16'b0000_0000_0000_0000;
array[6886] <= 16'b0000_0000_0000_0000;
array[6887] <= 16'b0000_0000_0000_0000;
array[6888] <= 16'b0000_0000_0000_0000;
array[6889] <= 16'b0000_0000_0000_0000;
array[6890] <= 16'b0000_0000_0000_0000;
array[6891] <= 16'b0000_0000_0000_0000;
array[6892] <= 16'b0000_0000_0000_0000;
array[6893] <= 16'b0000_0000_0000_0000;
array[6894] <= 16'b0000_0000_0000_0000;
array[6895] <= 16'b0000_0000_0000_0000;
array[6896] <= 16'b0000_0000_0000_0000;
array[6897] <= 16'b0000_0000_0000_0000;
array[6898] <= 16'b0000_0000_0000_0000;
array[6899] <= 16'b0000_0000_0000_0000;
array[6900] <= 16'b0000_0000_0000_0000;
array[6901] <= 16'b0000_0000_0000_0000;
array[6902] <= 16'b0000_0000_0000_0000;
array[6903] <= 16'b0000_0000_0000_0000;
array[6904] <= 16'b0000_0000_0000_0000;
array[6905] <= 16'b0000_0000_0000_0000;
array[6906] <= 16'b0000_0000_0000_0000;
array[6907] <= 16'b0000_0000_0000_0000;
array[6908] <= 16'b0000_0000_0000_0000;
array[6909] <= 16'b0000_0000_0000_0000;
array[6910] <= 16'b0000_0000_0000_0000;
array[6911] <= 16'b0000_0000_0000_0000;
array[6912] <= 16'b0000_0000_0000_0000;
array[6913] <= 16'b0000_0000_0000_0000;
array[6914] <= 16'b0000_0000_0000_0000;
array[6915] <= 16'b0000_0000_0000_0000;
array[6916] <= 16'b0000_0000_0000_0000;
array[6917] <= 16'b0000_0000_0000_0000;
array[6918] <= 16'b0000_0000_0000_0000;
array[6919] <= 16'b0000_0000_0000_0000;
array[6920] <= 16'b0000_0000_0000_0000;
array[6921] <= 16'b0000_0000_0000_0000;
array[6922] <= 16'b0000_0000_0000_0000;
array[6923] <= 16'b0000_0000_0000_0000;
array[6924] <= 16'b0000_0000_0000_0000;
array[6925] <= 16'b0000_0000_0000_0000;
array[6926] <= 16'b0000_0000_0000_0000;
array[6927] <= 16'b0000_0000_0000_0000;
array[6928] <= 16'b0000_0000_0000_0000;
array[6929] <= 16'b0000_0000_0000_0000;
array[6930] <= 16'b0000_0000_0000_0000;
array[6931] <= 16'b0000_0000_0000_0000;
array[6932] <= 16'b0000_0000_0000_0000;
array[6933] <= 16'b0000_0000_0000_0000;
array[6934] <= 16'b0000_0000_0000_0000;
array[6935] <= 16'b0000_0000_0000_0000;
array[6936] <= 16'b0000_0000_0000_0000;
array[6937] <= 16'b0000_0000_0000_0000;
array[6938] <= 16'b0000_0000_0000_0000;
array[6939] <= 16'b0000_0000_0000_0000;
array[6940] <= 16'b0000_0000_0000_0000;
array[6941] <= 16'b0000_0000_0000_0000;
array[6942] <= 16'b0000_0000_0000_0000;
array[6943] <= 16'b0000_0000_0000_0000;
array[6944] <= 16'b0000_0000_0000_0000;
array[6945] <= 16'b0000_0000_0000_0000;
array[6946] <= 16'b0000_0000_0000_0000;
array[6947] <= 16'b0000_0000_0000_0000;
array[6948] <= 16'b0000_0000_0000_0000;
array[6949] <= 16'b0000_0000_0000_0000;
array[6950] <= 16'b0000_0000_0000_0000;
array[6951] <= 16'b0000_0000_0000_0000;
array[6952] <= 16'b0000_0000_0000_0000;
array[6953] <= 16'b0000_0000_0000_0000;
array[6954] <= 16'b0000_0000_0000_0000;
array[6955] <= 16'b0000_0000_0000_0000;
array[6956] <= 16'b0000_0000_0000_0000;
array[6957] <= 16'b0000_0000_0000_0000;
array[6958] <= 16'b0000_0000_0000_0000;
array[6959] <= 16'b0000_0000_0000_0000;
array[6960] <= 16'b0000_0000_0000_0000;
array[6961] <= 16'b0000_0000_0000_0000;
array[6962] <= 16'b0000_0000_0000_0000;
array[6963] <= 16'b0000_0000_0000_0000;
array[6964] <= 16'b0000_0000_0000_0000;
array[6965] <= 16'b0000_0000_0000_0000;
array[6966] <= 16'b0000_0000_0000_0000;
array[6967] <= 16'b0000_0000_0000_0000;
array[6968] <= 16'b0000_0000_0000_0000;
array[6969] <= 16'b0000_0000_0000_0000;
array[6970] <= 16'b0000_0000_0000_0000;
array[6971] <= 16'b0000_0000_0000_0000;
array[6972] <= 16'b0000_0000_0000_0000;
array[6973] <= 16'b0000_0000_0000_0000;
array[6974] <= 16'b0000_0000_0000_0000;
array[6975] <= 16'b0000_0000_0000_0000;
array[6976] <= 16'b0000_0000_0000_0000;
array[6977] <= 16'b0000_0000_0000_0000;
array[6978] <= 16'b0000_0000_0000_0000;
array[6979] <= 16'b0000_0000_0000_0000;
array[6980] <= 16'b0000_0000_0000_0000;
array[6981] <= 16'b0000_0000_0000_0000;
array[6982] <= 16'b0000_0000_0000_0000;
array[6983] <= 16'b0000_0000_0000_0000;
array[6984] <= 16'b0000_0000_0000_0000;
array[6985] <= 16'b0000_0000_0000_0000;
array[6986] <= 16'b0000_0000_0000_0000;
array[6987] <= 16'b0000_0000_0000_0000;
array[6988] <= 16'b0000_0000_0000_0000;
array[6989] <= 16'b0000_0000_0000_0000;
array[6990] <= 16'b0000_0000_0000_0000;
array[6991] <= 16'b0000_0000_0000_0000;
array[6992] <= 16'b0000_0000_0000_0000;
array[6993] <= 16'b0000_0000_0000_0000;
array[6994] <= 16'b0000_0000_0000_0000;
array[6995] <= 16'b0000_0000_0000_0000;
array[6996] <= 16'b0000_0000_0000_0000;
array[6997] <= 16'b0000_0000_0000_0000;
array[6998] <= 16'b0000_0000_0000_0000;
array[6999] <= 16'b0000_0000_0000_0000;
array[7000] <= 16'b0000_0000_0000_0000;
array[7001] <= 16'b0000_0000_0000_0000;
array[7002] <= 16'b0000_0000_0000_0000;
array[7003] <= 16'b0000_0000_0000_0000;
array[7004] <= 16'b0000_0000_0000_0000;
array[7005] <= 16'b0000_0000_0000_0000;
array[7006] <= 16'b0000_0000_0000_0000;
array[7007] <= 16'b0000_0000_0000_0000;
array[7008] <= 16'b0000_0000_0000_0000;
array[7009] <= 16'b0000_0000_0000_0000;
array[7010] <= 16'b0000_0000_0000_0000;
array[7011] <= 16'b0000_0000_0000_0000;
array[7012] <= 16'b0000_0000_0000_0000;
array[7013] <= 16'b0000_0000_0000_0000;
array[7014] <= 16'b0000_0000_0000_0000;
array[7015] <= 16'b0000_0000_0000_0000;
array[7016] <= 16'b0000_0000_0000_0000;
array[7017] <= 16'b0000_0000_0000_0000;
array[7018] <= 16'b0000_0000_0000_0000;
array[7019] <= 16'b0000_0000_0000_0000;
array[7020] <= 16'b0000_0000_0000_0000;
array[7021] <= 16'b0000_0000_0000_0000;
array[7022] <= 16'b0000_0000_0000_0000;
array[7023] <= 16'b0000_0000_0000_0000;
array[7024] <= 16'b0000_0000_0000_0000;
array[7025] <= 16'b0000_0000_0000_0000;
array[7026] <= 16'b0000_0000_0000_0000;
array[7027] <= 16'b0000_0000_0000_0000;
array[7028] <= 16'b0000_0000_0000_0000;
array[7029] <= 16'b0000_0000_0000_0000;
array[7030] <= 16'b0000_0000_0000_0000;
array[7031] <= 16'b0000_0000_0000_0000;
array[7032] <= 16'b0000_0000_0000_0000;
array[7033] <= 16'b0000_0000_0000_0000;
array[7034] <= 16'b0000_0000_0000_0000;
array[7035] <= 16'b0000_0000_0000_0000;
array[7036] <= 16'b0000_0000_0000_0000;
array[7037] <= 16'b0000_0000_0000_0000;
array[7038] <= 16'b0000_0000_0000_0000;
array[7039] <= 16'b0000_0000_0000_0000;
array[7040] <= 16'b0000_0000_0000_0000;
array[7041] <= 16'b0000_0000_0000_0000;
array[7042] <= 16'b0000_0000_0000_0000;
array[7043] <= 16'b0000_0000_0000_0000;
array[7044] <= 16'b0000_0000_0000_0000;
array[7045] <= 16'b0000_0000_0000_0000;
array[7046] <= 16'b0000_0000_0000_0000;
array[7047] <= 16'b0000_0000_0000_0000;
array[7048] <= 16'b0000_0000_0000_0000;
array[7049] <= 16'b0000_0000_0000_0000;
array[7050] <= 16'b0000_0000_0000_0000;
array[7051] <= 16'b0000_0000_0000_0000;
array[7052] <= 16'b0000_0000_0000_0000;
array[7053] <= 16'b0000_0000_0000_0000;
array[7054] <= 16'b0000_0000_0000_0000;
array[7055] <= 16'b0000_0000_0000_0000;
array[7056] <= 16'b0000_0000_0000_0000;
array[7057] <= 16'b0000_0000_0000_0000;
array[7058] <= 16'b0000_0000_0000_0000;
array[7059] <= 16'b0000_0000_0000_0000;
array[7060] <= 16'b0000_0000_0000_0000;
array[7061] <= 16'b0000_0000_0000_0000;
array[7062] <= 16'b0000_0000_0000_0000;
array[7063] <= 16'b0000_0000_0000_0000;
array[7064] <= 16'b0000_0000_0000_0000;
array[7065] <= 16'b0000_0000_0000_0000;
array[7066] <= 16'b0000_0000_0000_0000;
array[7067] <= 16'b0000_0000_0000_0000;
array[7068] <= 16'b0000_0000_0000_0000;
array[7069] <= 16'b0000_0000_0000_0000;
array[7070] <= 16'b0000_0000_0000_0000;
array[7071] <= 16'b0000_0000_0000_0000;
array[7072] <= 16'b0000_0000_0000_0000;
array[7073] <= 16'b0000_0000_0000_0000;
array[7074] <= 16'b0000_0000_0000_0000;
array[7075] <= 16'b0000_0000_0000_0000;
array[7076] <= 16'b0000_0000_0000_0000;
array[7077] <= 16'b0000_0000_0000_0000;
array[7078] <= 16'b0000_0000_0000_0000;
array[7079] <= 16'b0000_0000_0000_0000;
array[7080] <= 16'b0000_0000_0000_0000;
array[7081] <= 16'b0000_0000_0000_0000;
array[7082] <= 16'b0000_0000_0000_0000;
array[7083] <= 16'b0000_0000_0000_0000;
array[7084] <= 16'b0000_0000_0000_0000;
array[7085] <= 16'b0000_0000_0000_0000;
array[7086] <= 16'b0000_0000_0000_0000;
array[7087] <= 16'b0000_0000_0000_0000;
array[7088] <= 16'b0000_0000_0000_0000;
array[7089] <= 16'b0000_0000_0000_0000;
array[7090] <= 16'b0000_0000_0000_0000;
array[7091] <= 16'b0000_0000_0000_0000;
array[7092] <= 16'b0000_0000_0000_0000;
array[7093] <= 16'b0000_0000_0000_0000;
array[7094] <= 16'b0000_0000_0000_0000;
array[7095] <= 16'b0000_0000_0000_0000;
array[7096] <= 16'b0000_0000_0000_0000;
array[7097] <= 16'b0000_0000_0000_0000;
array[7098] <= 16'b0000_0000_0000_0000;
array[7099] <= 16'b0000_0000_0000_0000;
array[7100] <= 16'b0000_0000_0000_0000;
array[7101] <= 16'b0000_0000_0000_0000;
array[7102] <= 16'b0000_0000_0000_0000;
array[7103] <= 16'b0000_0000_0000_0000;
array[7104] <= 16'b0000_0000_0000_0000;
array[7105] <= 16'b0000_0000_0000_0000;
array[7106] <= 16'b0000_0000_0000_0000;
array[7107] <= 16'b0000_0000_0000_0000;
array[7108] <= 16'b0000_0000_0000_0000;
array[7109] <= 16'b0000_0000_0000_0000;
array[7110] <= 16'b0000_0000_0000_0000;
array[7111] <= 16'b0000_0000_0000_0000;
array[7112] <= 16'b0000_0000_0000_0000;
array[7113] <= 16'b0000_0000_0000_0000;
array[7114] <= 16'b0000_0000_0000_0000;
array[7115] <= 16'b0000_0000_0000_0000;
array[7116] <= 16'b0000_0000_0000_0000;
array[7117] <= 16'b0000_0000_0000_0000;
array[7118] <= 16'b0000_0000_0000_0000;
array[7119] <= 16'b0000_0000_0000_0000;
array[7120] <= 16'b0000_0000_0000_0000;
array[7121] <= 16'b0000_0000_0000_0000;
array[7122] <= 16'b0000_0000_0000_0000;
array[7123] <= 16'b0000_0000_0000_0000;
array[7124] <= 16'b0000_0000_0000_0000;
array[7125] <= 16'b0000_0000_0000_0000;
array[7126] <= 16'b0000_0000_0000_0000;
array[7127] <= 16'b0000_0000_0000_0000;
array[7128] <= 16'b0000_0000_0000_0000;
array[7129] <= 16'b0000_0000_0000_0000;
array[7130] <= 16'b0000_0000_0000_0000;
array[7131] <= 16'b0000_0000_0000_0000;
array[7132] <= 16'b0000_0000_0000_0000;
array[7133] <= 16'b0000_0000_0000_0000;
array[7134] <= 16'b0000_0000_0000_0000;
array[7135] <= 16'b0000_0000_0000_0000;
array[7136] <= 16'b0000_0000_0000_0000;
array[7137] <= 16'b0000_0000_0000_0000;
array[7138] <= 16'b0000_0000_0000_0000;
array[7139] <= 16'b0000_0000_0000_0000;
array[7140] <= 16'b0000_0000_0000_0000;
array[7141] <= 16'b0000_0000_0000_0000;
array[7142] <= 16'b0000_0000_0000_0000;
array[7143] <= 16'b0000_0000_0000_0000;
array[7144] <= 16'b0000_0000_0000_0000;
array[7145] <= 16'b0000_0000_0000_0000;
array[7146] <= 16'b0000_0000_0000_0000;
array[7147] <= 16'b0000_0000_0000_0000;
array[7148] <= 16'b0000_0000_0000_0000;
array[7149] <= 16'b0000_0000_0000_0000;
array[7150] <= 16'b0000_0000_0000_0000;
array[7151] <= 16'b0000_0000_0000_0000;
array[7152] <= 16'b0000_0000_0000_0000;
array[7153] <= 16'b0000_0000_0000_0000;
array[7154] <= 16'b0000_0000_0000_0000;
array[7155] <= 16'b0000_0000_0000_0000;
array[7156] <= 16'b0000_0000_0000_0000;
array[7157] <= 16'b0000_0000_0000_0000;
array[7158] <= 16'b0000_0000_0000_0000;
array[7159] <= 16'b0000_0000_0000_0000;
array[7160] <= 16'b0000_0000_0000_0000;
array[7161] <= 16'b0000_0000_0000_0000;
array[7162] <= 16'b0000_0000_0000_0000;
array[7163] <= 16'b0000_0000_0000_0000;
array[7164] <= 16'b0000_0000_0000_0000;
array[7165] <= 16'b0000_0000_0000_0000;
array[7166] <= 16'b0000_0000_0000_0000;
array[7167] <= 16'b0000_0000_0000_0000;
array[7168] <= 16'b0000_0000_0000_0000;
array[7169] <= 16'b0000_0000_0000_0000;
array[7170] <= 16'b0000_0000_0000_0000;
array[7171] <= 16'b0000_0000_0000_0000;
array[7172] <= 16'b0000_0000_0000_0000;
array[7173] <= 16'b0000_0000_0000_0000;
array[7174] <= 16'b0000_0000_0000_0000;
array[7175] <= 16'b0000_0000_0000_0000;
array[7176] <= 16'b0000_0000_0000_0000;
array[7177] <= 16'b0000_0000_0000_0000;
array[7178] <= 16'b0000_0000_0000_0000;
array[7179] <= 16'b0000_0000_0000_0000;
array[7180] <= 16'b0000_0000_0000_0000;
array[7181] <= 16'b0000_0000_0000_0000;
array[7182] <= 16'b0000_0000_0000_0000;
array[7183] <= 16'b0000_0000_0000_0000;
array[7184] <= 16'b0000_0000_0000_0000;
array[7185] <= 16'b0000_0000_0000_0000;
array[7186] <= 16'b0000_0000_0000_0000;
array[7187] <= 16'b0000_0000_0000_0000;
array[7188] <= 16'b0000_0000_0000_0000;
array[7189] <= 16'b0000_0000_0000_0000;
array[7190] <= 16'b0000_0000_0000_0000;
array[7191] <= 16'b0000_0000_0000_0000;
array[7192] <= 16'b0000_0000_0000_0000;
array[7193] <= 16'b0000_0000_0000_0000;
array[7194] <= 16'b0000_0000_0000_0000;
array[7195] <= 16'b0000_0000_0000_0000;
array[7196] <= 16'b0000_0000_0000_0000;
array[7197] <= 16'b0000_0000_0000_0000;
array[7198] <= 16'b0000_0000_0000_0000;
array[7199] <= 16'b0000_0000_0000_0000;
array[7200] <= 16'b0000_0000_0000_0000;
array[7201] <= 16'b0000_0000_0000_0000;
array[7202] <= 16'b0000_0000_0000_0000;
array[7203] <= 16'b0000_0000_0000_0000;
array[7204] <= 16'b0000_0000_0000_0000;
array[7205] <= 16'b0000_0000_0000_0000;
array[7206] <= 16'b0000_0000_0000_0000;
array[7207] <= 16'b0000_0000_0000_0000;
array[7208] <= 16'b0000_0000_0000_0000;
array[7209] <= 16'b0000_0000_0000_0000;
array[7210] <= 16'b0000_0000_0000_0000;
array[7211] <= 16'b0000_0000_0000_0000;
array[7212] <= 16'b0000_0000_0000_0000;
array[7213] <= 16'b0000_0000_0000_0000;
array[7214] <= 16'b0000_0000_0000_0000;
array[7215] <= 16'b0000_0000_0000_0000;
array[7216] <= 16'b0000_0000_0000_0000;
array[7217] <= 16'b0000_0000_0000_0000;
array[7218] <= 16'b0000_0000_0000_0000;
array[7219] <= 16'b0000_0000_0000_0000;
array[7220] <= 16'b0000_0000_0000_0000;
array[7221] <= 16'b0000_0000_0000_0000;
array[7222] <= 16'b0000_0000_0000_0000;
array[7223] <= 16'b0000_0000_0000_0000;
array[7224] <= 16'b0000_0000_0000_0000;
array[7225] <= 16'b0000_0000_0000_0000;
array[7226] <= 16'b0000_0000_0000_0000;
array[7227] <= 16'b0000_0000_0000_0000;
array[7228] <= 16'b0000_0000_0000_0000;
array[7229] <= 16'b0000_0000_0000_0000;
array[7230] <= 16'b0000_0000_0000_0000;
array[7231] <= 16'b0000_0000_0000_0000;
array[7232] <= 16'b0000_0000_0000_0000;
array[7233] <= 16'b0000_0000_0000_0000;
array[7234] <= 16'b0000_0000_0000_0000;
array[7235] <= 16'b0000_0000_0000_0000;
array[7236] <= 16'b0000_0000_0000_0000;
array[7237] <= 16'b0000_0000_0000_0000;
array[7238] <= 16'b0000_0000_0000_0000;
array[7239] <= 16'b0000_0000_0000_0000;
array[7240] <= 16'b0000_0000_0000_0000;
array[7241] <= 16'b0000_0000_0000_0000;
array[7242] <= 16'b0000_0000_0000_0000;
array[7243] <= 16'b0000_0000_0000_0000;
array[7244] <= 16'b0000_0000_0000_0000;
array[7245] <= 16'b0000_0000_0000_0000;
array[7246] <= 16'b0000_0000_0000_0000;
array[7247] <= 16'b0000_0000_0000_0000;
array[7248] <= 16'b0000_0000_0000_0000;
array[7249] <= 16'b0000_0000_0000_0000;
array[7250] <= 16'b0000_0000_0000_0000;
array[7251] <= 16'b0000_0000_0000_0000;
array[7252] <= 16'b0000_0000_0000_0000;
array[7253] <= 16'b0000_0000_0000_0000;
array[7254] <= 16'b0000_0000_0000_0000;
array[7255] <= 16'b0000_0000_0000_0000;
array[7256] <= 16'b0000_0000_0000_0000;
array[7257] <= 16'b0000_0000_0000_0000;
array[7258] <= 16'b0000_0000_0000_0000;
array[7259] <= 16'b0000_0000_0000_0000;
array[7260] <= 16'b0000_0000_0000_0000;
array[7261] <= 16'b0000_0000_0000_0000;
array[7262] <= 16'b0000_0000_0000_0000;
array[7263] <= 16'b0000_0000_0000_0000;
array[7264] <= 16'b0000_0000_0000_0000;
array[7265] <= 16'b0000_0000_0000_0000;
array[7266] <= 16'b0000_0000_0000_0000;
array[7267] <= 16'b0000_0000_0000_0000;
array[7268] <= 16'b0000_0000_0000_0000;
array[7269] <= 16'b0000_0000_0000_0000;
array[7270] <= 16'b0000_0000_0000_0000;
array[7271] <= 16'b0000_0000_0000_0000;
array[7272] <= 16'b0000_0000_0000_0000;
array[7273] <= 16'b0000_0000_0000_0000;
array[7274] <= 16'b0000_0000_0000_0000;
array[7275] <= 16'b0000_0000_0000_0000;
array[7276] <= 16'b0000_0000_0000_0000;
array[7277] <= 16'b0000_0000_0000_0000;
array[7278] <= 16'b0000_0000_0000_0000;
array[7279] <= 16'b0000_0000_0000_0000;
array[7280] <= 16'b0000_0000_0000_0000;
array[7281] <= 16'b0000_0000_0000_0000;
array[7282] <= 16'b0000_0000_0000_0000;
array[7283] <= 16'b0000_0000_0000_0000;
array[7284] <= 16'b0000_0000_0000_0000;
array[7285] <= 16'b0000_0000_0000_0000;
array[7286] <= 16'b0000_0000_0000_0000;
array[7287] <= 16'b0000_0000_0000_0000;
array[7288] <= 16'b0000_0000_0000_0000;
array[7289] <= 16'b0000_0000_0000_0000;
array[7290] <= 16'b0000_0000_0000_0000;
array[7291] <= 16'b0000_0000_0000_0000;
array[7292] <= 16'b0000_0000_0000_0000;
array[7293] <= 16'b0000_0000_0000_0000;
array[7294] <= 16'b0000_0000_0000_0000;
array[7295] <= 16'b0000_0000_0000_0000;
array[7296] <= 16'b0000_0000_0000_0000;
array[7297] <= 16'b0000_0000_0000_0000;
array[7298] <= 16'b0000_0000_0000_0000;
array[7299] <= 16'b0000_0000_0000_0000;
array[7300] <= 16'b0000_0000_0000_0000;
array[7301] <= 16'b0000_0000_0000_0000;
array[7302] <= 16'b0000_0000_0000_0000;
array[7303] <= 16'b0000_0000_0000_0000;
array[7304] <= 16'b0000_0000_0000_0000;
array[7305] <= 16'b0000_0000_0000_0000;
array[7306] <= 16'b0000_0000_0000_0000;
array[7307] <= 16'b0000_0000_0000_0000;
array[7308] <= 16'b0000_0000_0000_0000;
array[7309] <= 16'b0000_0000_0000_0000;
array[7310] <= 16'b0000_0000_0000_0000;
array[7311] <= 16'b0000_0000_0000_0000;
array[7312] <= 16'b0000_0000_0000_0000;
array[7313] <= 16'b0000_0000_0000_0000;
array[7314] <= 16'b0000_0000_0000_0000;
array[7315] <= 16'b0000_0000_0000_0000;
array[7316] <= 16'b0000_0000_0000_0000;
array[7317] <= 16'b0000_0000_0000_0000;
array[7318] <= 16'b0000_0000_0000_0000;
array[7319] <= 16'b0000_0000_0000_0000;
array[7320] <= 16'b0000_0000_0000_0000;
array[7321] <= 16'b0000_0000_0000_0000;
array[7322] <= 16'b0000_0000_0000_0000;
array[7323] <= 16'b0000_0000_0000_0000;
array[7324] <= 16'b0000_0000_0000_0000;
array[7325] <= 16'b0000_0000_0000_0000;
array[7326] <= 16'b0000_0000_0000_0000;
array[7327] <= 16'b0000_0000_0000_0000;
array[7328] <= 16'b0000_0000_0000_0000;
array[7329] <= 16'b0000_0000_0000_0000;
array[7330] <= 16'b0000_0000_0000_0000;
array[7331] <= 16'b0000_0000_0000_0000;
array[7332] <= 16'b0000_0000_0000_0000;
array[7333] <= 16'b0000_0000_0000_0000;
array[7334] <= 16'b0000_0000_0000_0000;
array[7335] <= 16'b0000_0000_0000_0000;
array[7336] <= 16'b0000_0000_0000_0000;
array[7337] <= 16'b0000_0000_0000_0000;
array[7338] <= 16'b0000_0000_0000_0000;
array[7339] <= 16'b0000_0000_0000_0000;
array[7340] <= 16'b0000_0000_0000_0000;
array[7341] <= 16'b0000_0000_0000_0000;
array[7342] <= 16'b0000_0000_0000_0000;
array[7343] <= 16'b0000_0000_0000_0000;
array[7344] <= 16'b0000_0000_0000_0000;
array[7345] <= 16'b0000_0000_0000_0000;
array[7346] <= 16'b0000_0000_0000_0000;
array[7347] <= 16'b0000_0000_0000_0000;
array[7348] <= 16'b0000_0000_0000_0000;
array[7349] <= 16'b0000_0000_0000_0000;
array[7350] <= 16'b0000_0000_0000_0000;
array[7351] <= 16'b0000_0000_0000_0000;
array[7352] <= 16'b0000_0000_0000_0000;
array[7353] <= 16'b0000_0000_0000_0000;
array[7354] <= 16'b0000_0000_0000_0000;
array[7355] <= 16'b0000_0000_0000_0000;
array[7356] <= 16'b0000_0000_0000_0000;
array[7357] <= 16'b0000_0000_0000_0000;
array[7358] <= 16'b0000_0000_0000_0000;
array[7359] <= 16'b0000_0000_0000_0000;
array[7360] <= 16'b0000_0000_0000_0000;
array[7361] <= 16'b0000_0000_0000_0000;
array[7362] <= 16'b0000_0000_0000_0000;
array[7363] <= 16'b0000_0000_0000_0000;
array[7364] <= 16'b0000_0000_0000_0000;
array[7365] <= 16'b0000_0000_0000_0000;
array[7366] <= 16'b0000_0000_0000_0000;
array[7367] <= 16'b0000_0000_0000_0000;
array[7368] <= 16'b0000_0000_0000_0000;
array[7369] <= 16'b0000_0000_0000_0000;
array[7370] <= 16'b0000_0000_0000_0000;
array[7371] <= 16'b0000_0000_0000_0000;
array[7372] <= 16'b0000_0000_0000_0000;
array[7373] <= 16'b0000_0000_0000_0000;
array[7374] <= 16'b0000_0000_0000_0000;
array[7375] <= 16'b0000_0000_0000_0000;
array[7376] <= 16'b0000_0000_0000_0000;
array[7377] <= 16'b0000_0000_0000_0000;
array[7378] <= 16'b0000_0000_0000_0000;
array[7379] <= 16'b0000_0000_0000_0000;
array[7380] <= 16'b0000_0000_0000_0000;
array[7381] <= 16'b0000_0000_0000_0000;
array[7382] <= 16'b0000_0000_0000_0000;
array[7383] <= 16'b0000_0000_0000_0000;
array[7384] <= 16'b0000_0000_0000_0000;
array[7385] <= 16'b0000_0000_0000_0000;
array[7386] <= 16'b0000_0000_0000_0000;
array[7387] <= 16'b0000_0000_0000_0000;
array[7388] <= 16'b0000_0000_0000_0000;
array[7389] <= 16'b0000_0000_0000_0000;
array[7390] <= 16'b0000_0000_0000_0000;
array[7391] <= 16'b0000_0000_0000_0000;
array[7392] <= 16'b0000_0000_0000_0000;
array[7393] <= 16'b0000_0000_0000_0000;
array[7394] <= 16'b0000_0000_0000_0000;
array[7395] <= 16'b0000_0000_0000_0000;
array[7396] <= 16'b0000_0000_0000_0000;
array[7397] <= 16'b0000_0000_0000_0000;
array[7398] <= 16'b0000_0000_0000_0000;
array[7399] <= 16'b0000_0000_0000_0000;
array[7400] <= 16'b0000_0000_0000_0000;
array[7401] <= 16'b0000_0000_0000_0000;
array[7402] <= 16'b0000_0000_0000_0000;
array[7403] <= 16'b0000_0000_0000_0000;
array[7404] <= 16'b0000_0000_0000_0000;
array[7405] <= 16'b0000_0000_0000_0000;
array[7406] <= 16'b0000_0000_0000_0000;
array[7407] <= 16'b0000_0000_0000_0000;
array[7408] <= 16'b0000_0000_0000_0000;
array[7409] <= 16'b0000_0000_0000_0000;
array[7410] <= 16'b0000_0000_0000_0000;
array[7411] <= 16'b0000_0000_0000_0000;
array[7412] <= 16'b0000_0000_0000_0000;
array[7413] <= 16'b0000_0000_0000_0000;
array[7414] <= 16'b0000_0000_0000_0000;
array[7415] <= 16'b0000_0000_0000_0000;
array[7416] <= 16'b0000_0000_0000_0000;
array[7417] <= 16'b0000_0000_0000_0000;
array[7418] <= 16'b0000_0000_0000_0000;
array[7419] <= 16'b0000_0000_0000_0000;
array[7420] <= 16'b0000_0000_0000_0000;
array[7421] <= 16'b0000_0000_0000_0000;
array[7422] <= 16'b0000_0000_0000_0000;
array[7423] <= 16'b0000_0000_0000_0000;
array[7424] <= 16'b0000_0000_0000_0000;
array[7425] <= 16'b0000_0000_0000_0000;
array[7426] <= 16'b0000_0000_0000_0000;
array[7427] <= 16'b0000_0000_0000_0000;
array[7428] <= 16'b0000_0000_0000_0000;
array[7429] <= 16'b0000_0000_0000_0000;
array[7430] <= 16'b0000_0000_0000_0000;
array[7431] <= 16'b0000_0000_0000_0000;
array[7432] <= 16'b0000_0000_0000_0000;
array[7433] <= 16'b0000_0000_0000_0000;
array[7434] <= 16'b0000_0000_0000_0000;
array[7435] <= 16'b0000_0000_0000_0000;
array[7436] <= 16'b0000_0000_0000_0000;
array[7437] <= 16'b0000_0000_0000_0000;
array[7438] <= 16'b0000_0000_0000_0000;
array[7439] <= 16'b0000_0000_0000_0000;
array[7440] <= 16'b0000_0000_0000_0000;
array[7441] <= 16'b0000_0000_0000_0000;
array[7442] <= 16'b0000_0000_0000_0000;
array[7443] <= 16'b0000_0000_0000_0000;
array[7444] <= 16'b0000_0000_0000_0000;
array[7445] <= 16'b0000_0000_0000_0000;
array[7446] <= 16'b0000_0000_0000_0000;
array[7447] <= 16'b0000_0000_0000_0000;
array[7448] <= 16'b0000_0000_0000_0000;
array[7449] <= 16'b0000_0000_0000_0000;
array[7450] <= 16'b0000_0000_0000_0000;
array[7451] <= 16'b0000_0000_0000_0000;
array[7452] <= 16'b0000_0000_0000_0000;
array[7453] <= 16'b0000_0000_0000_0000;
array[7454] <= 16'b0000_0000_0000_0000;
array[7455] <= 16'b0000_0000_0000_0000;
array[7456] <= 16'b0000_0000_0000_0000;
array[7457] <= 16'b0000_0000_0000_0000;
array[7458] <= 16'b0000_0000_0000_0000;
array[7459] <= 16'b0000_0000_0000_0000;
array[7460] <= 16'b0000_0000_0000_0000;
array[7461] <= 16'b0000_0000_0000_0000;
array[7462] <= 16'b0000_0000_0000_0000;
array[7463] <= 16'b0000_0000_0000_0000;
array[7464] <= 16'b0000_0000_0000_0000;
array[7465] <= 16'b0000_0000_0000_0000;
array[7466] <= 16'b0000_0000_0000_0000;
array[7467] <= 16'b0000_0000_0000_0000;
array[7468] <= 16'b0000_0000_0000_0000;
array[7469] <= 16'b0000_0000_0000_0000;
array[7470] <= 16'b0000_0000_0000_0000;
array[7471] <= 16'b0000_0000_0000_0000;
array[7472] <= 16'b0000_0000_0000_0000;
array[7473] <= 16'b0000_0000_0000_0000;
array[7474] <= 16'b0000_0000_0000_0000;
array[7475] <= 16'b0000_0000_0000_0000;
array[7476] <= 16'b0000_0000_0000_0000;
array[7477] <= 16'b0000_0000_0000_0000;
array[7478] <= 16'b0000_0000_0000_0000;
array[7479] <= 16'b0000_0000_0000_0000;
array[7480] <= 16'b0000_0000_0000_0000;
array[7481] <= 16'b0000_0000_0000_0000;
array[7482] <= 16'b0000_0000_0000_0000;
array[7483] <= 16'b0000_0000_0000_0000;
array[7484] <= 16'b0000_0000_0000_0000;
array[7485] <= 16'b0000_0000_0000_0000;
array[7486] <= 16'b0000_0000_0000_0000;
array[7487] <= 16'b0000_0000_0000_0000;
array[7488] <= 16'b0000_0000_0000_0000;
array[7489] <= 16'b0000_0000_0000_0000;
array[7490] <= 16'b0000_0000_0000_0000;
array[7491] <= 16'b0000_0000_0000_0000;
array[7492] <= 16'b0000_0000_0000_0000;
array[7493] <= 16'b0000_0000_0000_0000;
array[7494] <= 16'b0000_0000_0000_0000;
array[7495] <= 16'b0000_0000_0000_0000;
array[7496] <= 16'b0000_0000_0000_0000;
array[7497] <= 16'b0000_0000_0000_0000;
array[7498] <= 16'b0000_0000_0000_0000;
array[7499] <= 16'b0000_0000_0000_0000;
array[7500] <= 16'b0000_0000_0000_0000;
array[7501] <= 16'b0000_0000_0000_0000;
array[7502] <= 16'b0000_0000_0000_0000;
array[7503] <= 16'b0000_0000_0000_0000;
array[7504] <= 16'b0000_0000_0000_0000;
array[7505] <= 16'b0000_0000_0000_0000;
array[7506] <= 16'b0000_0000_0000_0000;
array[7507] <= 16'b0000_0000_0000_0000;
array[7508] <= 16'b0000_0000_0000_0000;
array[7509] <= 16'b0000_0000_0000_0000;
array[7510] <= 16'b0000_0000_0000_0000;
array[7511] <= 16'b0000_0000_0000_0000;
array[7512] <= 16'b0000_0000_0000_0000;
array[7513] <= 16'b0000_0000_0000_0000;
array[7514] <= 16'b0000_0000_0000_0000;
array[7515] <= 16'b0000_0000_0000_0000;
array[7516] <= 16'b0000_0000_0000_0000;
array[7517] <= 16'b0000_0000_0000_0000;
array[7518] <= 16'b0000_0000_0000_0000;
array[7519] <= 16'b0000_0000_0000_0000;
array[7520] <= 16'b0000_0000_0000_0000;
array[7521] <= 16'b0000_0000_0000_0000;
array[7522] <= 16'b0000_0000_0000_0000;
array[7523] <= 16'b0000_0000_0000_0000;
array[7524] <= 16'b0000_0000_0000_0000;
array[7525] <= 16'b0000_0000_0000_0000;
array[7526] <= 16'b0000_0000_0000_0000;
array[7527] <= 16'b0000_0000_0000_0000;
array[7528] <= 16'b0000_0000_0000_0000;
array[7529] <= 16'b0000_0000_0000_0000;
array[7530] <= 16'b0000_0000_0000_0000;
array[7531] <= 16'b0000_0000_0000_0000;
array[7532] <= 16'b0000_0000_0000_0000;
array[7533] <= 16'b0000_0000_0000_0000;
array[7534] <= 16'b0000_0000_0000_0000;
array[7535] <= 16'b0000_0000_0000_0000;
array[7536] <= 16'b0000_0000_0000_0000;
array[7537] <= 16'b0000_0000_0000_0000;
array[7538] <= 16'b0000_0000_0000_0000;
array[7539] <= 16'b0000_0000_0000_0000;
array[7540] <= 16'b0000_0000_0000_0000;
array[7541] <= 16'b0000_0000_0000_0000;
array[7542] <= 16'b0000_0000_0000_0000;
array[7543] <= 16'b0000_0000_0000_0000;
array[7544] <= 16'b0000_0000_0000_0000;
array[7545] <= 16'b0000_0000_0000_0000;
array[7546] <= 16'b0000_0000_0000_0000;
array[7547] <= 16'b0000_0000_0000_0000;
array[7548] <= 16'b0000_0000_0000_0000;
array[7549] <= 16'b0000_0000_0000_0000;
array[7550] <= 16'b0000_0000_0000_0000;
array[7551] <= 16'b0000_0000_0000_0000;
array[7552] <= 16'b0000_0000_0000_0000;
array[7553] <= 16'b0000_0000_0000_0000;
array[7554] <= 16'b0000_0000_0000_0000;
array[7555] <= 16'b0000_0000_0000_0000;
array[7556] <= 16'b0000_0000_0000_0000;
array[7557] <= 16'b0000_0000_0000_0000;
array[7558] <= 16'b0000_0000_0000_0000;
array[7559] <= 16'b0000_0000_0000_0000;
array[7560] <= 16'b0000_0000_0000_0000;
array[7561] <= 16'b0000_0000_0000_0000;
array[7562] <= 16'b0000_0000_0000_0000;
array[7563] <= 16'b0000_0000_0000_0000;
array[7564] <= 16'b0000_0000_0000_0000;
array[7565] <= 16'b0000_0000_0000_0000;
array[7566] <= 16'b0000_0000_0000_0000;
array[7567] <= 16'b0000_0000_0000_0000;
array[7568] <= 16'b0000_0000_0000_0000;
array[7569] <= 16'b0000_0000_0000_0000;
array[7570] <= 16'b0000_0000_0000_0000;
array[7571] <= 16'b0000_0000_0000_0000;
array[7572] <= 16'b0000_0000_0000_0000;
array[7573] <= 16'b0000_0000_0000_0000;
array[7574] <= 16'b0000_0000_0000_0000;
array[7575] <= 16'b0000_0000_0000_0000;
array[7576] <= 16'b0000_0000_0000_0000;
array[7577] <= 16'b0000_0000_0000_0000;
array[7578] <= 16'b0000_0000_0000_0000;
array[7579] <= 16'b0000_0000_0000_0000;
array[7580] <= 16'b0000_0000_0000_0000;
array[7581] <= 16'b0000_0000_0000_0000;
array[7582] <= 16'b0000_0000_0000_0000;
array[7583] <= 16'b0000_0000_0000_0000;
array[7584] <= 16'b0000_0000_0000_0000;
array[7585] <= 16'b0000_0000_0000_0000;
array[7586] <= 16'b0000_0000_0000_0000;
array[7587] <= 16'b0000_0000_0000_0000;
array[7588] <= 16'b0000_0000_0000_0000;
array[7589] <= 16'b0000_0000_0000_0000;
array[7590] <= 16'b0000_0000_0000_0000;
array[7591] <= 16'b0000_0000_0000_0000;
array[7592] <= 16'b0000_0000_0000_0000;
array[7593] <= 16'b0000_0000_0000_0000;
array[7594] <= 16'b0000_0000_0000_0000;
array[7595] <= 16'b0000_0000_0000_0000;
array[7596] <= 16'b0000_0000_0000_0000;
array[7597] <= 16'b0000_0000_0000_0000;
array[7598] <= 16'b0000_0000_0000_0000;
array[7599] <= 16'b0000_0000_0000_0000;
array[7600] <= 16'b0000_0000_0000_0000;
array[7601] <= 16'b0000_0000_0000_0000;
array[7602] <= 16'b0000_0000_0000_0000;
array[7603] <= 16'b0000_0000_0000_0000;
array[7604] <= 16'b0000_0000_0000_0000;
array[7605] <= 16'b0000_0000_0000_0000;
array[7606] <= 16'b0000_0000_0000_0000;
array[7607] <= 16'b0000_0000_0000_0000;
array[7608] <= 16'b0000_0000_0000_0000;
array[7609] <= 16'b0000_0000_0000_0000;
array[7610] <= 16'b0000_0000_0000_0000;
array[7611] <= 16'b0000_0000_0000_0000;
array[7612] <= 16'b0000_0000_0000_0000;
array[7613] <= 16'b0000_0000_0000_0000;
array[7614] <= 16'b0000_0000_0000_0000;
array[7615] <= 16'b0000_0000_0000_0000;
array[7616] <= 16'b0000_0000_0000_0000;
array[7617] <= 16'b0000_0000_0000_0000;
array[7618] <= 16'b0000_0000_0000_0000;
array[7619] <= 16'b0000_0000_0000_0000;
array[7620] <= 16'b0000_0000_0000_0000;
array[7621] <= 16'b0000_0000_0000_0000;
array[7622] <= 16'b0000_0000_0000_0000;
array[7623] <= 16'b0000_0000_0000_0000;
array[7624] <= 16'b0000_0000_0000_0000;
array[7625] <= 16'b0000_0000_0000_0000;
array[7626] <= 16'b0000_0000_0000_0000;
array[7627] <= 16'b0000_0000_0000_0000;
array[7628] <= 16'b0000_0000_0000_0000;
array[7629] <= 16'b0000_0000_0000_0000;
array[7630] <= 16'b0000_0000_0000_0000;
array[7631] <= 16'b0000_0000_0000_0000;
array[7632] <= 16'b0000_0000_0000_0000;
array[7633] <= 16'b0000_0000_0000_0000;
array[7634] <= 16'b0000_0000_0000_0000;
array[7635] <= 16'b0000_0000_0000_0000;
array[7636] <= 16'b0000_0000_0000_0000;
array[7637] <= 16'b0000_0000_0000_0000;
array[7638] <= 16'b0000_0000_0000_0000;
array[7639] <= 16'b0000_0000_0000_0000;
array[7640] <= 16'b0000_0000_0000_0000;
array[7641] <= 16'b0000_0000_0000_0000;
array[7642] <= 16'b0000_0000_0000_0000;
array[7643] <= 16'b0000_0000_0000_0000;
array[7644] <= 16'b0000_0000_0000_0000;
array[7645] <= 16'b0000_0000_0000_0000;
array[7646] <= 16'b0000_0000_0000_0000;
array[7647] <= 16'b0000_0000_0000_0000;
array[7648] <= 16'b0000_0000_0000_0000;
array[7649] <= 16'b0000_0000_0000_0000;
array[7650] <= 16'b0000_0000_0000_0000;
array[7651] <= 16'b0000_0000_0000_0000;
array[7652] <= 16'b0000_0000_0000_0000;
array[7653] <= 16'b0000_0000_0000_0000;
array[7654] <= 16'b0000_0000_0000_0000;
array[7655] <= 16'b0000_0000_0000_0000;
array[7656] <= 16'b0000_0000_0000_0000;
array[7657] <= 16'b0000_0000_0000_0000;
array[7658] <= 16'b0000_0000_0000_0000;
array[7659] <= 16'b0000_0000_0000_0000;
array[7660] <= 16'b0000_0000_0000_0000;
array[7661] <= 16'b0000_0000_0000_0000;
array[7662] <= 16'b0000_0000_0000_0000;
array[7663] <= 16'b0000_0000_0000_0000;
array[7664] <= 16'b0000_0000_0000_0000;
array[7665] <= 16'b0000_0000_0000_0000;
array[7666] <= 16'b0000_0000_0000_0000;
array[7667] <= 16'b0000_0000_0000_0000;
array[7668] <= 16'b0000_0000_0000_0000;
array[7669] <= 16'b0000_0000_0000_0000;
array[7670] <= 16'b0000_0000_0000_0000;
array[7671] <= 16'b0000_0000_0000_0000;
array[7672] <= 16'b0000_0000_0000_0000;
array[7673] <= 16'b0000_0000_0000_0000;
array[7674] <= 16'b0000_0000_0000_0000;
array[7675] <= 16'b0000_0000_0000_0000;
array[7676] <= 16'b0000_0000_0000_0000;
array[7677] <= 16'b0000_0000_0000_0000;
array[7678] <= 16'b0000_0000_0000_0000;
array[7679] <= 16'b0000_0000_0000_0000;
array[7680] <= 16'b0000_0000_0000_0000;
array[7681] <= 16'b0000_0000_0000_0000;
array[7682] <= 16'b0000_0000_0000_0000;
array[7683] <= 16'b0000_0000_0000_0000;
array[7684] <= 16'b0000_0000_0000_0000;
array[7685] <= 16'b0000_0000_0000_0000;
array[7686] <= 16'b0000_0000_0000_0000;
array[7687] <= 16'b0000_0000_0000_0000;
array[7688] <= 16'b0000_0000_0000_0000;
array[7689] <= 16'b0000_0000_0000_0000;
array[7690] <= 16'b0000_0000_0000_0000;
array[7691] <= 16'b0000_0000_0000_0000;
array[7692] <= 16'b0000_0000_0000_0000;
array[7693] <= 16'b0000_0000_0000_0000;
array[7694] <= 16'b0000_0000_0000_0000;
array[7695] <= 16'b0000_0000_0000_0000;
array[7696] <= 16'b0000_0000_0000_0000;
array[7697] <= 16'b0000_0000_0000_0000;
array[7698] <= 16'b0000_0000_0000_0000;
array[7699] <= 16'b0000_0000_0000_0000;
array[7700] <= 16'b0000_0000_0000_0000;
array[7701] <= 16'b0000_0000_0000_0000;
array[7702] <= 16'b0000_0000_0000_0000;
array[7703] <= 16'b0000_0000_0000_0000;
array[7704] <= 16'b0000_0000_0000_0000;
array[7705] <= 16'b0000_0000_0000_0000;
array[7706] <= 16'b0000_0000_0000_0000;
array[7707] <= 16'b0000_0000_0000_0000;
array[7708] <= 16'b0000_0000_0000_0000;
array[7709] <= 16'b0000_0000_0000_0000;
array[7710] <= 16'b0000_0000_0000_0000;
array[7711] <= 16'b0000_0000_0000_0000;
array[7712] <= 16'b0000_0000_0000_0000;
array[7713] <= 16'b0000_0000_0000_0000;
array[7714] <= 16'b0000_0000_0000_0000;
array[7715] <= 16'b0000_0000_0000_0000;
array[7716] <= 16'b0000_0000_0000_0000;
array[7717] <= 16'b0000_0000_0000_0000;
array[7718] <= 16'b0000_0000_0000_0000;
array[7719] <= 16'b0000_0000_0000_0000;
array[7720] <= 16'b0000_0000_0000_0000;
array[7721] <= 16'b0000_0000_0000_0000;
array[7722] <= 16'b0000_0000_0000_0000;
array[7723] <= 16'b0000_0000_0000_0000;
array[7724] <= 16'b0000_0000_0000_0000;
array[7725] <= 16'b0000_0000_0000_0000;
array[7726] <= 16'b0000_0000_0000_0000;
array[7727] <= 16'b0000_0000_0000_0000;
array[7728] <= 16'b0000_0000_0000_0000;
array[7729] <= 16'b0000_0000_0000_0000;
array[7730] <= 16'b0000_0000_0000_0000;
array[7731] <= 16'b0000_0000_0000_0000;
array[7732] <= 16'b0000_0000_0000_0000;
array[7733] <= 16'b0000_0000_0000_0000;
array[7734] <= 16'b0000_0000_0000_0000;
array[7735] <= 16'b0000_0000_0000_0000;
array[7736] <= 16'b0000_0000_0000_0000;
array[7737] <= 16'b0000_0000_0000_0000;
array[7738] <= 16'b0000_0000_0000_0000;
array[7739] <= 16'b0000_0000_0000_0000;
array[7740] <= 16'b0000_0000_0000_0000;
array[7741] <= 16'b0000_0000_0000_0000;
array[7742] <= 16'b0000_0000_0000_0000;
array[7743] <= 16'b0000_0000_0000_0000;
array[7744] <= 16'b0000_0000_0000_0000;
array[7745] <= 16'b0000_0000_0000_0000;
array[7746] <= 16'b0000_0000_0000_0000;
array[7747] <= 16'b0000_0000_0000_0000;
array[7748] <= 16'b0000_0000_0000_0000;
array[7749] <= 16'b0000_0000_0000_0000;
array[7750] <= 16'b0000_0000_0000_0000;
array[7751] <= 16'b0000_0000_0000_0000;
array[7752] <= 16'b0000_0000_0000_0000;
array[7753] <= 16'b0000_0000_0000_0000;
array[7754] <= 16'b0000_0000_0000_0000;
array[7755] <= 16'b0000_0000_0000_0000;
array[7756] <= 16'b0000_0000_0000_0000;
array[7757] <= 16'b0000_0000_0000_0000;
array[7758] <= 16'b0000_0000_0000_0000;
array[7759] <= 16'b0000_0000_0000_0000;
array[7760] <= 16'b0000_0000_0000_0000;
array[7761] <= 16'b0000_0000_0000_0000;
array[7762] <= 16'b0000_0000_0000_0000;
array[7763] <= 16'b0000_0000_0000_0000;
array[7764] <= 16'b0000_0000_0000_0000;
array[7765] <= 16'b0000_0000_0000_0000;
array[7766] <= 16'b0000_0000_0000_0000;
array[7767] <= 16'b0000_0000_0000_0000;
array[7768] <= 16'b0000_0000_0000_0000;
array[7769] <= 16'b0000_0000_0000_0000;
array[7770] <= 16'b0000_0000_0000_0000;
array[7771] <= 16'b0000_0000_0000_0000;
array[7772] <= 16'b0000_0000_0000_0000;
array[7773] <= 16'b0000_0000_0000_0000;
array[7774] <= 16'b0000_0000_0000_0000;
array[7775] <= 16'b0000_0000_0000_0000;
array[7776] <= 16'b0000_0000_0000_0000;
array[7777] <= 16'b0000_0000_0000_0000;
array[7778] <= 16'b0000_0000_0000_0000;
array[7779] <= 16'b0000_0000_0000_0000;
array[7780] <= 16'b0000_0000_0000_0000;
array[7781] <= 16'b0000_0000_0000_0000;
array[7782] <= 16'b0000_0000_0000_0000;
array[7783] <= 16'b0000_0000_0000_0000;
array[7784] <= 16'b0000_0000_0000_0000;
array[7785] <= 16'b0000_0000_0000_0000;
array[7786] <= 16'b0000_0000_0000_0000;
array[7787] <= 16'b0000_0000_0000_0000;
array[7788] <= 16'b0000_0000_0000_0000;
array[7789] <= 16'b0000_0000_0000_0000;
array[7790] <= 16'b0000_0000_0000_0000;
array[7791] <= 16'b0000_0000_0000_0000;
array[7792] <= 16'b0000_0000_0000_0000;
array[7793] <= 16'b0000_0000_0000_0000;
array[7794] <= 16'b0000_0000_0000_0000;
array[7795] <= 16'b0000_0000_0000_0000;
array[7796] <= 16'b0000_0000_0000_0000;
array[7797] <= 16'b0000_0000_0000_0000;
array[7798] <= 16'b0000_0000_0000_0000;
array[7799] <= 16'b0000_0000_0000_0000;
array[7800] <= 16'b0000_0000_0000_0000;
array[7801] <= 16'b0000_0000_0000_0000;
array[7802] <= 16'b0000_0000_0000_0000;
array[7803] <= 16'b0000_0000_0000_0000;
array[7804] <= 16'b0000_0000_0000_0000;
array[7805] <= 16'b0000_0000_0000_0000;
array[7806] <= 16'b0000_0000_0000_0000;
array[7807] <= 16'b0000_0000_0000_0000;
array[7808] <= 16'b0000_0000_0000_0000;
array[7809] <= 16'b0000_0000_0000_0000;
array[7810] <= 16'b0000_0000_0000_0000;
array[7811] <= 16'b0000_0000_0000_0000;
array[7812] <= 16'b0000_0000_0000_0000;
array[7813] <= 16'b0000_0000_0000_0000;
array[7814] <= 16'b0000_0000_0000_0000;
array[7815] <= 16'b0000_0000_0000_0000;
array[7816] <= 16'b0000_0000_0000_0000;
array[7817] <= 16'b0000_0000_0000_0000;
array[7818] <= 16'b0000_0000_0000_0000;
array[7819] <= 16'b0000_0000_0000_0000;
array[7820] <= 16'b0000_0000_0000_0000;
array[7821] <= 16'b0000_0000_0000_0000;
array[7822] <= 16'b0000_0000_0000_0000;
array[7823] <= 16'b0000_0000_0000_0000;
array[7824] <= 16'b0000_0000_0000_0000;
array[7825] <= 16'b0000_0000_0000_0000;
array[7826] <= 16'b0000_0000_0000_0000;
array[7827] <= 16'b0000_0000_0000_0000;
array[7828] <= 16'b0000_0000_0000_0000;
array[7829] <= 16'b0000_0000_0000_0000;
array[7830] <= 16'b0000_0000_0000_0000;
array[7831] <= 16'b0000_0000_0000_0000;
array[7832] <= 16'b0000_0000_0000_0000;
array[7833] <= 16'b0000_0000_0000_0000;
array[7834] <= 16'b0000_0000_0000_0000;
array[7835] <= 16'b0000_0000_0000_0000;
array[7836] <= 16'b0000_0000_0000_0000;
array[7837] <= 16'b0000_0000_0000_0000;
array[7838] <= 16'b0000_0000_0000_0000;
array[7839] <= 16'b0000_0000_0000_0000;
array[7840] <= 16'b0000_0000_0000_0000;
array[7841] <= 16'b0000_0000_0000_0000;
array[7842] <= 16'b0000_0000_0000_0000;
array[7843] <= 16'b0000_0000_0000_0000;
array[7844] <= 16'b0000_0000_0000_0000;
array[7845] <= 16'b0000_0000_0000_0000;
array[7846] <= 16'b0000_0000_0000_0000;
array[7847] <= 16'b0000_0000_0000_0000;
array[7848] <= 16'b0000_0000_0000_0000;
array[7849] <= 16'b0000_0000_0000_0000;
array[7850] <= 16'b0000_0000_0000_0000;
array[7851] <= 16'b0000_0000_0000_0000;
array[7852] <= 16'b0000_0000_0000_0000;
array[7853] <= 16'b0000_0000_0000_0000;
array[7854] <= 16'b0000_0000_0000_0000;
array[7855] <= 16'b0000_0000_0000_0000;
array[7856] <= 16'b0000_0000_0000_0000;
array[7857] <= 16'b0000_0000_0000_0000;
array[7858] <= 16'b0000_0000_0000_0000;
array[7859] <= 16'b0000_0000_0000_0000;
array[7860] <= 16'b0000_0000_0000_0000;
array[7861] <= 16'b0000_0000_0000_0000;
array[7862] <= 16'b0000_0000_0000_0000;
array[7863] <= 16'b0000_0000_0000_0000;
array[7864] <= 16'b0000_0000_0000_0000;
array[7865] <= 16'b0000_0000_0000_0000;
array[7866] <= 16'b0000_0000_0000_0000;
array[7867] <= 16'b0000_0000_0000_0000;
array[7868] <= 16'b0000_0000_0000_0000;
array[7869] <= 16'b0000_0000_0000_0000;
array[7870] <= 16'b0000_0000_0000_0000;
array[7871] <= 16'b0000_0000_0000_0000;
array[7872] <= 16'b0000_0000_0000_0000;
array[7873] <= 16'b0000_0000_0000_0000;
array[7874] <= 16'b0000_0000_0000_0000;
array[7875] <= 16'b0000_0000_0000_0000;
array[7876] <= 16'b0000_0000_0000_0000;
array[7877] <= 16'b0000_0000_0000_0000;
array[7878] <= 16'b0000_0000_0000_0000;
array[7879] <= 16'b0000_0000_0000_0000;
array[7880] <= 16'b0000_0000_0000_0000;
array[7881] <= 16'b0000_0000_0000_0000;
array[7882] <= 16'b0000_0000_0000_0000;
array[7883] <= 16'b0000_0000_0000_0000;
array[7884] <= 16'b0000_0000_0000_0000;
array[7885] <= 16'b0000_0000_0000_0000;
array[7886] <= 16'b0000_0000_0000_0000;
array[7887] <= 16'b0000_0000_0000_0000;
array[7888] <= 16'b0000_0000_0000_0000;
array[7889] <= 16'b0000_0000_0000_0000;
array[7890] <= 16'b0000_0000_0000_0000;
array[7891] <= 16'b0000_0000_0000_0000;
array[7892] <= 16'b0000_0000_0000_0000;
array[7893] <= 16'b0000_0000_0000_0000;
array[7894] <= 16'b0000_0000_0000_0000;
array[7895] <= 16'b0000_0000_0000_0000;
array[7896] <= 16'b0000_0000_0000_0000;
array[7897] <= 16'b0000_0000_0000_0000;
array[7898] <= 16'b0000_0000_0000_0000;
array[7899] <= 16'b0000_0000_0000_0000;
array[7900] <= 16'b0000_0000_0000_0000;
array[7901] <= 16'b0000_0000_0000_0000;
array[7902] <= 16'b0000_0000_0000_0000;
array[7903] <= 16'b0000_0000_0000_0000;
array[7904] <= 16'b0000_0000_0000_0000;
array[7905] <= 16'b0000_0000_0000_0000;
array[7906] <= 16'b0000_0000_0000_0000;
array[7907] <= 16'b0000_0000_0000_0000;
array[7908] <= 16'b0000_0000_0000_0000;
array[7909] <= 16'b0000_0000_0000_0000;
array[7910] <= 16'b0000_0000_0000_0000;
array[7911] <= 16'b0000_0000_0000_0000;
array[7912] <= 16'b0000_0000_0000_0000;
array[7913] <= 16'b0000_0000_0000_0000;
array[7914] <= 16'b0000_0000_0000_0000;
array[7915] <= 16'b0000_0000_0000_0000;
array[7916] <= 16'b0000_0000_0000_0000;
array[7917] <= 16'b0000_0000_0000_0000;
array[7918] <= 16'b0000_0000_0000_0000;
array[7919] <= 16'b0000_0000_0000_0000;
array[7920] <= 16'b0000_0000_0000_0000;
array[7921] <= 16'b0000_0000_0000_0000;
array[7922] <= 16'b0000_0000_0000_0000;
array[7923] <= 16'b0000_0000_0000_0000;
array[7924] <= 16'b0000_0000_0000_0000;
array[7925] <= 16'b0000_0000_0000_0000;
array[7926] <= 16'b0000_0000_0000_0000;
array[7927] <= 16'b0000_0000_0000_0000;
array[7928] <= 16'b0000_0000_0000_0000;
array[7929] <= 16'b0000_0000_0000_0000;
array[7930] <= 16'b0000_0000_0000_0000;
array[7931] <= 16'b0000_0000_0000_0000;
array[7932] <= 16'b0000_0000_0000_0000;
array[7933] <= 16'b0000_0000_0000_0000;
array[7934] <= 16'b0000_0000_0000_0000;
array[7935] <= 16'b0000_0000_0000_0000;
array[7936] <= 16'b0000_0000_0000_0000;
array[7937] <= 16'b0000_0000_0000_0000;
array[7938] <= 16'b0000_0000_0000_0000;
array[7939] <= 16'b0000_0000_0000_0000;
array[7940] <= 16'b0000_0000_0000_0000;
array[7941] <= 16'b0000_0000_0000_0000;
array[7942] <= 16'b0000_0000_0000_0000;
array[7943] <= 16'b0000_0000_0000_0000;
array[7944] <= 16'b0000_0000_0000_0000;
array[7945] <= 16'b0000_0000_0000_0000;
array[7946] <= 16'b0000_0000_0000_0000;
array[7947] <= 16'b0000_0000_0000_0000;
array[7948] <= 16'b0000_0000_0000_0000;
array[7949] <= 16'b0000_0000_0000_0000;
array[7950] <= 16'b0000_0000_0000_0000;
array[7951] <= 16'b0000_0000_0000_0000;
array[7952] <= 16'b0000_0000_0000_0000;
array[7953] <= 16'b0000_0000_0000_0000;
array[7954] <= 16'b0000_0000_0000_0000;
array[7955] <= 16'b0000_0000_0000_0000;
array[7956] <= 16'b0000_0000_0000_0000;
array[7957] <= 16'b0000_0000_0000_0000;
array[7958] <= 16'b0000_0000_0000_0000;
array[7959] <= 16'b0000_0000_0000_0000;
array[7960] <= 16'b0000_0000_0000_0000;
array[7961] <= 16'b0000_0000_0000_0000;
array[7962] <= 16'b0000_0000_0000_0000;
array[7963] <= 16'b0000_0000_0000_0000;
array[7964] <= 16'b0000_0000_0000_0000;
array[7965] <= 16'b0000_0000_0000_0000;
array[7966] <= 16'b0000_0000_0000_0000;
array[7967] <= 16'b0000_0000_0000_0000;
array[7968] <= 16'b0000_0000_0000_0000;
array[7969] <= 16'b0000_0000_0000_0000;
array[7970] <= 16'b0000_0000_0000_0000;
array[7971] <= 16'b0000_0000_0000_0000;
array[7972] <= 16'b0000_0000_0000_0000;
array[7973] <= 16'b0000_0000_0000_0000;
array[7974] <= 16'b0000_0000_0000_0000;
array[7975] <= 16'b0000_0000_0000_0000;
array[7976] <= 16'b0000_0000_0000_0000;
array[7977] <= 16'b0000_0000_0000_0000;
array[7978] <= 16'b0000_0000_0000_0000;
array[7979] <= 16'b0000_0000_0000_0000;
array[7980] <= 16'b0000_0000_0000_0000;
array[7981] <= 16'b0000_0000_0000_0000;
array[7982] <= 16'b0000_0000_0000_0000;
array[7983] <= 16'b0000_0000_0000_0000;
array[7984] <= 16'b0000_0000_0000_0000;
array[7985] <= 16'b0000_0000_0000_0000;
array[7986] <= 16'b0000_0000_0000_0000;
array[7987] <= 16'b0000_0000_0000_0000;
array[7988] <= 16'b0000_0000_0000_0000;
array[7989] <= 16'b0000_0000_0000_0000;
array[7990] <= 16'b0000_0000_0000_0000;
array[7991] <= 16'b0000_0000_0000_0000;
array[7992] <= 16'b0000_0000_0000_0000;
array[7993] <= 16'b0000_0000_0000_0000;
array[7994] <= 16'b0000_0000_0000_0000;
array[7995] <= 16'b0000_0000_0000_0000;
array[7996] <= 16'b0000_0000_0000_0000;
array[7997] <= 16'b0000_0000_0000_0000;
array[7998] <= 16'b0000_0000_0000_0000;
array[7999] <= 16'b0000_0000_0000_0000;
array[8000] <= 16'b0000_0000_0000_0000;
array[8001] <= 16'b0000_0000_0000_0000;
array[8002] <= 16'b0000_0000_0000_0000;
array[8003] <= 16'b0000_0000_0000_0000;
array[8004] <= 16'b0000_0000_0000_0000;
array[8005] <= 16'b0000_0000_0000_0000;
array[8006] <= 16'b0000_0000_0000_0000;
array[8007] <= 16'b0000_0000_0000_0000;
array[8008] <= 16'b0000_0000_0000_0000;
array[8009] <= 16'b0000_0000_0000_0000;
array[8010] <= 16'b0000_0000_0000_0000;
array[8011] <= 16'b0000_0000_0000_0000;
array[8012] <= 16'b0000_0000_0000_0000;
array[8013] <= 16'b0000_0000_0000_0000;
array[8014] <= 16'b0000_0000_0000_0000;
array[8015] <= 16'b0000_0000_0000_0000;
array[8016] <= 16'b0000_0000_0000_0000;
array[8017] <= 16'b0000_0000_0000_0000;
array[8018] <= 16'b0000_0000_0000_0000;
array[8019] <= 16'b0000_0000_0000_0000;
array[8020] <= 16'b0000_0000_0000_0000;
array[8021] <= 16'b0000_0000_0000_0000;
array[8022] <= 16'b0000_0000_0000_0000;
array[8023] <= 16'b0000_0000_0000_0000;
array[8024] <= 16'b0000_0000_0000_0000;
array[8025] <= 16'b0000_0000_0000_0000;
array[8026] <= 16'b0000_0000_0000_0000;
array[8027] <= 16'b0000_0000_0000_0000;
array[8028] <= 16'b0000_0000_0000_0000;
array[8029] <= 16'b0000_0000_0000_0000;
array[8030] <= 16'b0000_0000_0000_0000;
array[8031] <= 16'b0000_0000_0000_0000;
array[8032] <= 16'b0000_0000_0000_0000;
array[8033] <= 16'b0000_0000_0000_0000;
array[8034] <= 16'b0000_0000_0000_0000;
array[8035] <= 16'b0000_0000_0000_0000;
array[8036] <= 16'b0000_0000_0000_0000;
array[8037] <= 16'b0000_0000_0000_0000;
array[8038] <= 16'b0000_0000_0000_0000;
array[8039] <= 16'b0000_0000_0000_0000;
array[8040] <= 16'b0000_0000_0000_0000;
array[8041] <= 16'b0000_0000_0000_0000;
array[8042] <= 16'b0000_0000_0000_0000;
array[8043] <= 16'b0000_0000_0000_0000;
array[8044] <= 16'b0000_0000_0000_0000;
array[8045] <= 16'b0000_0000_0000_0000;
array[8046] <= 16'b0000_0000_0000_0000;
array[8047] <= 16'b0000_0000_0000_0000;
array[8048] <= 16'b0000_0000_0000_0000;
array[8049] <= 16'b0000_0000_0000_0000;
array[8050] <= 16'b0000_0000_0000_0000;
array[8051] <= 16'b0000_0000_0000_0000;
array[8052] <= 16'b0000_0000_0000_0000;
array[8053] <= 16'b0000_0000_0000_0000;
array[8054] <= 16'b0000_0000_0000_0000;
array[8055] <= 16'b0000_0000_0000_0000;
array[8056] <= 16'b0000_0000_0000_0000;
array[8057] <= 16'b0000_0000_0000_0000;
array[8058] <= 16'b0000_0000_0000_0000;
array[8059] <= 16'b0000_0000_0000_0000;
array[8060] <= 16'b0000_0000_0000_0000;
array[8061] <= 16'b0000_0000_0000_0000;
array[8062] <= 16'b0000_0000_0000_0000;
array[8063] <= 16'b0000_0000_0000_0000;
array[8064] <= 16'b0000_0000_0000_0000;
array[8065] <= 16'b0000_0000_0000_0000;
array[8066] <= 16'b0000_0000_0000_0000;
array[8067] <= 16'b0000_0000_0000_0000;
array[8068] <= 16'b0000_0000_0000_0000;
array[8069] <= 16'b0000_0000_0000_0000;
array[8070] <= 16'b0000_0000_0000_0000;
array[8071] <= 16'b0000_0000_0000_0000;
array[8072] <= 16'b0000_0000_0000_0000;
array[8073] <= 16'b0000_0000_0000_0000;
array[8074] <= 16'b0000_0000_0000_0000;
array[8075] <= 16'b0000_0000_0000_0000;
array[8076] <= 16'b0000_0000_0000_0000;
array[8077] <= 16'b0000_0000_0000_0000;
array[8078] <= 16'b0000_0000_0000_0000;
array[8079] <= 16'b0000_0000_0000_0000;
array[8080] <= 16'b0000_0000_0000_0000;
array[8081] <= 16'b0000_0000_0000_0000;
array[8082] <= 16'b0000_0000_0000_0000;
array[8083] <= 16'b0000_0000_0000_0000;
array[8084] <= 16'b0000_0000_0000_0000;
array[8085] <= 16'b0000_0000_0000_0000;
array[8086] <= 16'b0000_0000_0000_0000;
array[8087] <= 16'b0000_0000_0000_0000;
array[8088] <= 16'b0000_0000_0000_0000;
array[8089] <= 16'b0000_0000_0000_0000;
array[8090] <= 16'b0000_0000_0000_0000;
array[8091] <= 16'b0000_0000_0000_0000;
array[8092] <= 16'b0000_0000_0000_0000;
array[8093] <= 16'b0000_0000_0000_0000;
array[8094] <= 16'b0000_0000_0000_0000;
array[8095] <= 16'b0000_0000_0000_0000;
array[8096] <= 16'b0000_0000_0000_0000;
array[8097] <= 16'b0000_0000_0000_0000;
array[8098] <= 16'b0000_0000_0000_0000;
array[8099] <= 16'b0000_0000_0000_0000;
array[8100] <= 16'b0000_0000_0000_0000;
array[8101] <= 16'b0000_0000_0000_0000;
array[8102] <= 16'b0000_0000_0000_0000;
array[8103] <= 16'b0000_0000_0000_0000;
array[8104] <= 16'b0000_0000_0000_0000;
array[8105] <= 16'b0000_0000_0000_0000;
array[8106] <= 16'b0000_0000_0000_0000;
array[8107] <= 16'b0000_0000_0000_0000;
array[8108] <= 16'b0000_0000_0000_0000;
array[8109] <= 16'b0000_0000_0000_0000;
array[8110] <= 16'b0000_0000_0000_0000;
array[8111] <= 16'b0000_0000_0000_0000;
array[8112] <= 16'b0000_0000_0000_0000;
array[8113] <= 16'b0000_0000_0000_0000;
array[8114] <= 16'b0000_0000_0000_0000;
array[8115] <= 16'b0000_0000_0000_0000;
array[8116] <= 16'b0000_0000_0000_0000;
array[8117] <= 16'b0000_0000_0000_0000;
array[8118] <= 16'b0000_0000_0000_0000;
array[8119] <= 16'b0000_0000_0000_0000;
array[8120] <= 16'b0000_0000_0000_0000;
array[8121] <= 16'b0000_0000_0000_0000;
array[8122] <= 16'b0000_0000_0000_0000;
array[8123] <= 16'b0000_0000_0000_0000;
array[8124] <= 16'b0000_0000_0000_0000;
array[8125] <= 16'b0000_0000_0000_0000;
array[8126] <= 16'b0000_0000_0000_0000;
array[8127] <= 16'b0000_0000_0000_0000;
array[8128] <= 16'b0000_0000_0000_0000;
array[8129] <= 16'b0000_0000_0000_0000;
array[8130] <= 16'b0000_0000_0000_0000;
array[8131] <= 16'b0000_0000_0000_0000;
array[8132] <= 16'b0000_0000_0000_0000;
array[8133] <= 16'b0000_0000_0000_0000;
array[8134] <= 16'b0000_0000_0000_0000;
array[8135] <= 16'b0000_0000_0000_0000;
array[8136] <= 16'b0000_0000_0000_0000;
array[8137] <= 16'b0000_0000_0000_0000;
array[8138] <= 16'b0000_0000_0000_0000;
array[8139] <= 16'b0000_0000_0000_0000;
array[8140] <= 16'b0000_0000_0000_0000;
array[8141] <= 16'b0000_0000_0000_0000;
array[8142] <= 16'b0000_0000_0000_0000;
array[8143] <= 16'b0000_0000_0000_0000;
array[8144] <= 16'b0000_0000_0000_0000;
array[8145] <= 16'b0000_0000_0000_0000;
array[8146] <= 16'b0000_0000_0000_0000;
array[8147] <= 16'b0000_0000_0000_0000;
array[8148] <= 16'b0000_0000_0000_0000;
array[8149] <= 16'b0000_0000_0000_0000;
array[8150] <= 16'b0000_0000_0000_0000;
array[8151] <= 16'b0000_0000_0000_0000;
array[8152] <= 16'b0000_0000_0000_0000;
array[8153] <= 16'b0000_0000_0000_0000;
array[8154] <= 16'b0000_0000_0000_0000;
array[8155] <= 16'b0000_0000_0000_0000;
array[8156] <= 16'b0000_0000_0000_0000;
array[8157] <= 16'b0000_0000_0000_0000;
array[8158] <= 16'b0000_0000_0000_0000;
array[8159] <= 16'b0000_0000_0000_0000;
array[8160] <= 16'b0000_0000_0000_0000;
array[8161] <= 16'b0000_0000_0000_0000;
array[8162] <= 16'b0000_0000_0000_0000;
array[8163] <= 16'b0000_0000_0000_0000;
array[8164] <= 16'b0000_0000_0000_0000;
array[8165] <= 16'b0000_0000_0000_0000;
array[8166] <= 16'b0000_0000_0000_0000;
array[8167] <= 16'b0000_0000_0000_0000;
array[8168] <= 16'b0000_0000_0000_0000;
array[8169] <= 16'b0000_0000_0000_0000;
array[8170] <= 16'b0000_0000_0000_0000;
array[8171] <= 16'b0000_0000_0000_0000;
array[8172] <= 16'b0000_0000_0000_0000;
array[8173] <= 16'b0000_0000_0000_0000;
array[8174] <= 16'b0000_0000_0000_0000;
array[8175] <= 16'b0000_0000_0000_0000;
array[8176] <= 16'b0000_0000_0000_0000;
array[8177] <= 16'b0000_0000_0000_0000;
array[8178] <= 16'b0000_0000_0000_0000;
array[8179] <= 16'b0000_0000_0000_0000;
array[8180] <= 16'b0000_0000_0000_0000;
array[8181] <= 16'b0000_0000_0000_0000;
array[8182] <= 16'b0000_0000_0000_0000;
array[8183] <= 16'b0000_0000_0000_0000;
array[8184] <= 16'b0000_0000_0000_0000;
array[8185] <= 16'b0000_0000_0000_0000;
array[8186] <= 16'b0000_0000_0000_0000;
array[8187] <= 16'b0000_0000_0000_0000;
array[8188] <= 16'b0000_0000_0000_0000;
array[8189] <= 16'b0000_0000_0000_0000;
array[8190] <= 16'b0000_0000_0000_0000;
array[8191] <= 16'b0000_0000_0000_0000;
array[8192] <= 16'b0000_0000_0000_0000;
array[8193] <= 16'b0000_0000_0000_0000;
array[8194] <= 16'b0000_0000_0000_0000;
array[8195] <= 16'b0000_0000_0000_0000;
array[8196] <= 16'b0000_0000_0000_0000;
array[8197] <= 16'b0000_0000_0000_0000;
array[8198] <= 16'b0000_0000_0000_0000;
array[8199] <= 16'b0000_0000_0000_0000;
array[8200] <= 16'b0000_0000_0000_0000;
array[8201] <= 16'b0000_0000_0000_0000;
array[8202] <= 16'b0000_0000_0000_0000;
array[8203] <= 16'b0000_0000_0000_0000;
array[8204] <= 16'b0000_0000_0000_0000;
array[8205] <= 16'b0000_0000_0000_0000;
array[8206] <= 16'b0000_0000_0000_0000;
array[8207] <= 16'b0000_0000_0000_0000;
array[8208] <= 16'b0000_0000_0000_0000;
array[8209] <= 16'b0000_0000_0000_0000;
array[8210] <= 16'b0000_0000_0000_0000;
array[8211] <= 16'b0000_0000_0000_0000;
array[8212] <= 16'b0000_0000_0000_0000;
array[8213] <= 16'b0000_0000_0000_0000;
array[8214] <= 16'b0000_0000_0000_0000;
array[8215] <= 16'b0000_0000_0000_0000;
array[8216] <= 16'b0000_0000_0000_0000;
array[8217] <= 16'b0000_0000_0000_0000;
array[8218] <= 16'b0000_0000_0000_0000;
array[8219] <= 16'b0000_0000_0000_0000;
array[8220] <= 16'b0000_0000_0000_0000;
array[8221] <= 16'b0000_0000_0000_0000;
array[8222] <= 16'b0000_0000_0000_0000;
array[8223] <= 16'b0000_0000_0000_0000;
array[8224] <= 16'b0000_0000_0000_0000;
array[8225] <= 16'b0000_0000_0000_0000;
array[8226] <= 16'b0000_0000_0000_0000;
array[8227] <= 16'b0000_0000_0000_0000;
array[8228] <= 16'b0000_0000_0000_0000;
array[8229] <= 16'b0000_0000_0000_0000;
array[8230] <= 16'b0000_0000_0000_0000;
array[8231] <= 16'b0000_0000_0000_0000;
array[8232] <= 16'b0000_0000_0000_0000;
array[8233] <= 16'b0000_0000_0000_0000;
array[8234] <= 16'b0000_0000_0000_0000;
array[8235] <= 16'b0000_0000_0000_0000;
array[8236] <= 16'b0000_0000_0000_0000;
array[8237] <= 16'b0000_0000_0000_0000;
array[8238] <= 16'b0000_0000_0000_0000;
array[8239] <= 16'b0000_0000_0000_0000;
array[8240] <= 16'b0000_0000_0000_0000;
array[8241] <= 16'b0000_0000_0000_0000;
array[8242] <= 16'b0000_0000_0000_0000;
array[8243] <= 16'b0000_0000_0000_0000;
array[8244] <= 16'b0000_0000_0000_0000;
array[8245] <= 16'b0000_0000_0000_0000;
array[8246] <= 16'b0000_0000_0000_0000;
array[8247] <= 16'b0000_0000_0000_0000;
array[8248] <= 16'b0000_0000_0000_0000;
array[8249] <= 16'b0000_0000_0000_0000;
array[8250] <= 16'b0000_0000_0000_0000;
array[8251] <= 16'b0000_0000_0000_0000;
array[8252] <= 16'b0000_0000_0000_0000;
array[8253] <= 16'b0000_0000_0000_0000;
array[8254] <= 16'b0000_0000_0000_0000;
array[8255] <= 16'b0000_0000_0000_0000;
array[8256] <= 16'b0000_0000_0000_0000;
array[8257] <= 16'b0000_0000_0000_0000;
array[8258] <= 16'b0000_0000_0000_0000;
array[8259] <= 16'b0000_0000_0000_0000;
array[8260] <= 16'b0000_0000_0000_0000;
array[8261] <= 16'b0000_0000_0000_0000;
array[8262] <= 16'b0000_0000_0000_0000;
array[8263] <= 16'b0000_0000_0000_0000;
array[8264] <= 16'b0000_0000_0000_0000;
array[8265] <= 16'b0000_0000_0000_0000;
array[8266] <= 16'b0000_0000_0000_0000;
array[8267] <= 16'b0000_0000_0000_0000;
array[8268] <= 16'b0000_0000_0000_0000;
array[8269] <= 16'b0000_0000_0000_0000;
array[8270] <= 16'b0000_0000_0000_0000;
array[8271] <= 16'b0000_0000_0000_0000;
array[8272] <= 16'b0000_0000_0000_0000;
array[8273] <= 16'b0000_0000_0000_0000;
array[8274] <= 16'b0000_0000_0000_0000;
array[8275] <= 16'b0000_0000_0000_0000;
array[8276] <= 16'b0000_0000_0000_0000;
array[8277] <= 16'b0000_0000_0000_0000;
array[8278] <= 16'b0000_0000_0000_0000;
array[8279] <= 16'b0000_0000_0000_0000;
array[8280] <= 16'b0000_0000_0000_0000;
array[8281] <= 16'b0000_0000_0000_0000;
array[8282] <= 16'b0000_0000_0000_0000;
array[8283] <= 16'b0000_0000_0000_0000;
array[8284] <= 16'b0000_0000_0000_0000;
array[8285] <= 16'b0000_0000_0000_0000;
array[8286] <= 16'b0000_0000_0000_0000;
array[8287] <= 16'b0000_0000_0000_0000;
array[8288] <= 16'b0000_0000_0000_0000;
array[8289] <= 16'b0000_0000_0000_0000;
array[8290] <= 16'b0000_0000_0000_0000;
array[8291] <= 16'b0000_0000_0000_0000;
array[8292] <= 16'b0000_0000_0000_0000;
array[8293] <= 16'b0000_0000_0000_0000;
array[8294] <= 16'b0000_0000_0000_0000;
array[8295] <= 16'b0000_0000_0000_0000;
array[8296] <= 16'b0000_0000_0000_0000;
array[8297] <= 16'b0000_0000_0000_0000;
array[8298] <= 16'b0000_0000_0000_0000;
array[8299] <= 16'b0000_0000_0000_0000;
array[8300] <= 16'b0000_0000_0000_0000;
array[8301] <= 16'b0000_0000_0000_0000;
array[8302] <= 16'b0000_0000_0000_0000;
array[8303] <= 16'b0000_0000_0000_0000;
array[8304] <= 16'b0000_0000_0000_0000;
array[8305] <= 16'b0000_0000_0000_0000;
array[8306] <= 16'b0000_0000_0000_0000;
array[8307] <= 16'b0000_0000_0000_0000;
array[8308] <= 16'b0000_0000_0000_0000;
array[8309] <= 16'b0000_0000_0000_0000;
array[8310] <= 16'b0000_0000_0000_0000;
array[8311] <= 16'b0000_0000_0000_0000;
array[8312] <= 16'b0000_0000_0000_0000;
array[8313] <= 16'b0000_0000_0000_0000;
array[8314] <= 16'b0000_0000_0000_0000;
array[8315] <= 16'b0000_0000_0000_0000;
array[8316] <= 16'b0000_0000_0000_0000;
array[8317] <= 16'b0000_0000_0000_0000;
array[8318] <= 16'b0000_0000_0000_0000;
array[8319] <= 16'b0000_0000_0000_0000;
array[8320] <= 16'b0000_0000_0000_0000;
array[8321] <= 16'b0000_0000_0000_0000;
array[8322] <= 16'b0000_0000_0000_0000;
array[8323] <= 16'b0000_0000_0000_0000;
array[8324] <= 16'b0000_0000_0000_0000;
array[8325] <= 16'b0000_0000_0000_0000;
array[8326] <= 16'b0000_0000_0000_0000;
array[8327] <= 16'b0000_0000_0000_0000;
array[8328] <= 16'b0000_0000_0000_0000;
array[8329] <= 16'b0000_0000_0000_0000;
array[8330] <= 16'b0000_0000_0000_0000;
array[8331] <= 16'b0000_0000_0000_0000;
array[8332] <= 16'b0000_0000_0000_0000;
array[8333] <= 16'b0000_0000_0000_0000;
array[8334] <= 16'b0000_0000_0000_0000;
array[8335] <= 16'b0000_0000_0000_0000;
array[8336] <= 16'b0000_0000_0000_0000;
array[8337] <= 16'b0000_0000_0000_0000;
array[8338] <= 16'b0000_0000_0000_0000;
array[8339] <= 16'b0000_0000_0000_0000;
array[8340] <= 16'b0000_0000_0000_0000;
array[8341] <= 16'b0000_0000_0000_0000;
array[8342] <= 16'b0000_0000_0000_0000;
array[8343] <= 16'b0000_0000_0000_0000;
array[8344] <= 16'b0000_0000_0000_0000;
array[8345] <= 16'b0000_0000_0000_0000;
array[8346] <= 16'b0000_0000_0000_0000;
array[8347] <= 16'b0000_0000_0000_0000;
array[8348] <= 16'b0000_0000_0000_0000;
array[8349] <= 16'b0000_0000_0000_0000;
array[8350] <= 16'b0000_0000_0000_0000;
array[8351] <= 16'b0000_0000_0000_0000;
array[8352] <= 16'b0000_0000_0000_0000;
array[8353] <= 16'b0000_0000_0000_0000;
array[8354] <= 16'b0000_0000_0000_0000;
array[8355] <= 16'b0000_0000_0000_0000;
array[8356] <= 16'b0000_0000_0000_0000;
array[8357] <= 16'b0000_0000_0000_0000;
array[8358] <= 16'b0000_0000_0000_0000;
array[8359] <= 16'b0000_0000_0000_0000;
array[8360] <= 16'b0000_0000_0000_0000;
array[8361] <= 16'b0000_0000_0000_0000;
array[8362] <= 16'b0000_0000_0000_0000;
array[8363] <= 16'b0000_0000_0000_0000;
array[8364] <= 16'b0000_0000_0000_0000;
array[8365] <= 16'b0000_0000_0000_0000;
array[8366] <= 16'b0000_0000_0000_0000;
array[8367] <= 16'b0000_0000_0000_0000;
array[8368] <= 16'b0000_0000_0000_0000;
array[8369] <= 16'b0000_0000_0000_0000;
array[8370] <= 16'b0000_0000_0000_0000;
array[8371] <= 16'b0000_0000_0000_0000;
array[8372] <= 16'b0000_0000_0000_0000;
array[8373] <= 16'b0000_0000_0000_0000;
array[8374] <= 16'b0000_0000_0000_0000;
array[8375] <= 16'b0000_0000_0000_0000;
array[8376] <= 16'b0000_0000_0000_0000;
array[8377] <= 16'b0000_0000_0000_0000;
array[8378] <= 16'b0000_0000_0000_0000;
array[8379] <= 16'b0000_0000_0000_0000;
array[8380] <= 16'b0000_0000_0000_0000;
array[8381] <= 16'b0000_0000_0000_0000;
array[8382] <= 16'b0000_0000_0000_0000;
array[8383] <= 16'b0000_0000_0000_0000;
array[8384] <= 16'b0000_0000_0000_0000;
array[8385] <= 16'b0000_0000_0000_0000;
array[8386] <= 16'b0000_0000_0000_0000;
array[8387] <= 16'b0000_0000_0000_0000;
array[8388] <= 16'b0000_0000_0000_0000;
array[8389] <= 16'b0000_0000_0000_0000;
array[8390] <= 16'b0000_0000_0000_0000;
array[8391] <= 16'b0000_0000_0000_0000;
array[8392] <= 16'b0000_0000_0000_0000;
array[8393] <= 16'b0000_0000_0000_0000;
array[8394] <= 16'b0000_0000_0000_0000;
array[8395] <= 16'b0000_0000_0000_0000;
array[8396] <= 16'b0000_0000_0000_0000;
array[8397] <= 16'b0000_0000_0000_0000;
array[8398] <= 16'b0000_0000_0000_0000;
array[8399] <= 16'b0000_0000_0000_0000;
array[8400] <= 16'b0000_0000_0000_0000;
array[8401] <= 16'b0000_0000_0000_0000;
array[8402] <= 16'b0000_0000_0000_0000;
array[8403] <= 16'b0000_0000_0000_0000;
array[8404] <= 16'b0000_0000_0000_0000;
array[8405] <= 16'b0000_0000_0000_0000;
array[8406] <= 16'b0000_0000_0000_0000;
array[8407] <= 16'b0000_0000_0000_0000;
array[8408] <= 16'b0000_0000_0000_0000;
array[8409] <= 16'b0000_0000_0000_0000;
array[8410] <= 16'b0000_0000_0000_0000;
array[8411] <= 16'b0000_0000_0000_0000;
array[8412] <= 16'b0000_0000_0000_0000;
array[8413] <= 16'b0000_0000_0000_0000;
array[8414] <= 16'b0000_0000_0000_0000;
array[8415] <= 16'b0000_0000_0000_0000;
array[8416] <= 16'b0000_0000_0000_0000;
array[8417] <= 16'b0000_0000_0000_0000;
array[8418] <= 16'b0000_0000_0000_0000;
array[8419] <= 16'b0000_0000_0000_0000;
array[8420] <= 16'b0000_0000_0000_0000;
array[8421] <= 16'b0000_0000_0000_0000;
array[8422] <= 16'b0000_0000_0000_0000;
array[8423] <= 16'b0000_0000_0000_0000;
array[8424] <= 16'b0000_0000_0000_0000;
array[8425] <= 16'b0000_0000_0000_0000;
array[8426] <= 16'b0000_0000_0000_0000;
array[8427] <= 16'b0000_0000_0000_0000;
array[8428] <= 16'b0000_0000_0000_0000;
array[8429] <= 16'b0000_0000_0000_0000;
array[8430] <= 16'b0000_0000_0000_0000;
array[8431] <= 16'b0000_0000_0000_0000;
array[8432] <= 16'b0000_0000_0000_0000;
array[8433] <= 16'b0000_0000_0000_0000;
array[8434] <= 16'b0000_0000_0000_0000;
array[8435] <= 16'b0000_0000_0000_0000;
array[8436] <= 16'b0000_0000_0000_0000;
array[8437] <= 16'b0000_0000_0000_0000;
array[8438] <= 16'b0000_0000_0000_0000;
array[8439] <= 16'b0000_0000_0000_0000;
array[8440] <= 16'b0000_0000_0000_0000;
array[8441] <= 16'b0000_0000_0000_0000;
array[8442] <= 16'b0000_0000_0000_0000;
array[8443] <= 16'b0000_0000_0000_0000;
array[8444] <= 16'b0000_0000_0000_0000;
array[8445] <= 16'b0000_0000_0000_0000;
array[8446] <= 16'b0000_0000_0000_0000;
array[8447] <= 16'b0000_0000_0000_0000;
array[8448] <= 16'b0000_0000_0000_0000;
array[8449] <= 16'b0000_0000_0000_0000;
array[8450] <= 16'b0000_0000_0000_0000;
array[8451] <= 16'b0000_0000_0000_0000;
array[8452] <= 16'b0000_0000_0000_0000;
array[8453] <= 16'b0000_0000_0000_0000;
array[8454] <= 16'b0000_0000_0000_0000;
array[8455] <= 16'b0000_0000_0000_0000;
array[8456] <= 16'b0000_0000_0000_0000;
array[8457] <= 16'b0000_0000_0000_0000;
array[8458] <= 16'b0000_0000_0000_0000;
array[8459] <= 16'b0000_0000_0000_0000;
array[8460] <= 16'b0000_0000_0000_0000;
array[8461] <= 16'b0000_0000_0000_0000;
array[8462] <= 16'b0000_0000_0000_0000;
array[8463] <= 16'b0000_0000_0000_0000;
array[8464] <= 16'b0000_0000_0000_0000;
array[8465] <= 16'b0000_0000_0000_0000;
array[8466] <= 16'b0000_0000_0000_0000;
array[8467] <= 16'b0000_0000_0000_0000;
array[8468] <= 16'b0000_0000_0000_0000;
array[8469] <= 16'b0000_0000_0000_0000;
array[8470] <= 16'b0000_0000_0000_0000;
array[8471] <= 16'b0000_0000_0000_0000;
array[8472] <= 16'b0000_0000_0000_0000;
array[8473] <= 16'b0000_0000_0000_0000;
array[8474] <= 16'b0000_0000_0000_0000;
array[8475] <= 16'b0000_0000_0000_0000;
array[8476] <= 16'b0000_0000_0000_0000;
array[8477] <= 16'b0000_0000_0000_0000;
array[8478] <= 16'b0000_0000_0000_0000;
array[8479] <= 16'b0000_0000_0000_0000;
array[8480] <= 16'b0000_0000_0000_0000;
array[8481] <= 16'b0000_0000_0000_0000;
array[8482] <= 16'b0000_0000_0000_0000;
array[8483] <= 16'b0000_0000_0000_0000;
array[8484] <= 16'b0000_0000_0000_0000;
array[8485] <= 16'b0000_0000_0000_0000;
array[8486] <= 16'b0000_0000_0000_0000;
array[8487] <= 16'b0000_0000_0000_0000;
array[8488] <= 16'b0000_0000_0000_0000;
array[8489] <= 16'b0000_0000_0000_0000;
array[8490] <= 16'b0000_0000_0000_0000;
array[8491] <= 16'b0000_0000_0000_0000;
array[8492] <= 16'b0000_0000_0000_0000;
array[8493] <= 16'b0000_0000_0000_0000;
array[8494] <= 16'b0000_0000_0000_0000;
array[8495] <= 16'b0000_0000_0000_0000;
array[8496] <= 16'b0000_0000_0000_0000;
array[8497] <= 16'b0000_0000_0000_0000;
array[8498] <= 16'b0000_0000_0000_0000;
array[8499] <= 16'b0000_0000_0000_0000;
array[8500] <= 16'b0000_0000_0000_0000;
array[8501] <= 16'b0000_0000_0000_0000;
array[8502] <= 16'b0000_0000_0000_0000;
array[8503] <= 16'b0000_0000_0000_0000;
array[8504] <= 16'b0000_0000_0000_0000;
array[8505] <= 16'b0000_0000_0000_0000;
array[8506] <= 16'b0000_0000_0000_0000;
array[8507] <= 16'b0000_0000_0000_0000;
array[8508] <= 16'b0000_0000_0000_0000;
array[8509] <= 16'b0000_0000_0000_0000;
array[8510] <= 16'b0000_0000_0000_0000;
array[8511] <= 16'b0000_0000_0000_0000;
array[8512] <= 16'b0000_0000_0000_0000;
array[8513] <= 16'b0000_0000_0000_0000;
array[8514] <= 16'b0000_0000_0000_0000;
array[8515] <= 16'b0000_0000_0000_0000;
array[8516] <= 16'b0000_0000_0000_0000;
array[8517] <= 16'b0000_0000_0000_0000;
array[8518] <= 16'b0000_0000_0000_0000;
array[8519] <= 16'b0000_0000_0000_0000;
array[8520] <= 16'b0000_0000_0000_0000;
array[8521] <= 16'b0000_0000_0000_0000;
array[8522] <= 16'b0000_0000_0000_0000;
array[8523] <= 16'b0000_0000_0000_0000;
array[8524] <= 16'b0000_0000_0000_0000;
array[8525] <= 16'b0000_0000_0000_0000;
array[8526] <= 16'b0000_0000_0000_0000;
array[8527] <= 16'b0000_0000_0000_0000;
array[8528] <= 16'b0000_0000_0000_0000;
array[8529] <= 16'b0000_0000_0000_0000;
array[8530] <= 16'b0000_0000_0000_0000;
array[8531] <= 16'b0000_0000_0000_0000;
array[8532] <= 16'b0000_0000_0000_0000;
array[8533] <= 16'b0000_0000_0000_0000;
array[8534] <= 16'b0000_0000_0000_0000;
array[8535] <= 16'b0000_0000_0000_0000;
array[8536] <= 16'b0000_0000_0000_0000;
array[8537] <= 16'b0000_0000_0000_0000;
array[8538] <= 16'b0000_0000_0000_0000;
array[8539] <= 16'b0000_0000_0000_0000;
array[8540] <= 16'b0000_0000_0000_0000;
array[8541] <= 16'b0000_0000_0000_0000;
array[8542] <= 16'b0000_0000_0000_0000;
array[8543] <= 16'b0000_0000_0000_0000;
array[8544] <= 16'b0000_0000_0000_0000;
array[8545] <= 16'b0000_0000_0000_0000;
array[8546] <= 16'b0000_0000_0000_0000;
array[8547] <= 16'b0000_0000_0000_0000;
array[8548] <= 16'b0000_0000_0000_0000;
array[8549] <= 16'b0000_0000_0000_0000;
array[8550] <= 16'b0000_0000_0000_0000;
array[8551] <= 16'b0000_0000_0000_0000;
array[8552] <= 16'b0000_0000_0000_0000;
array[8553] <= 16'b0000_0000_0000_0000;
array[8554] <= 16'b0000_0000_0000_0000;
array[8555] <= 16'b0000_0000_0000_0000;
array[8556] <= 16'b0000_0000_0000_0000;
array[8557] <= 16'b0000_0000_0000_0000;
array[8558] <= 16'b0000_0000_0000_0000;
array[8559] <= 16'b0000_0000_0000_0000;
array[8560] <= 16'b0000_0000_0000_0000;
array[8561] <= 16'b0000_0000_0000_0000;
array[8562] <= 16'b0000_0000_0000_0000;
array[8563] <= 16'b0000_0000_0000_0000;
array[8564] <= 16'b0000_0000_0000_0000;
array[8565] <= 16'b0000_0000_0000_0000;
array[8566] <= 16'b0000_0000_0000_0000;
array[8567] <= 16'b0000_0000_0000_0000;
array[8568] <= 16'b0000_0000_0000_0000;
array[8569] <= 16'b0000_0000_0000_0000;
array[8570] <= 16'b0000_0000_0000_0000;
array[8571] <= 16'b0000_0000_0000_0000;
array[8572] <= 16'b0000_0000_0000_0000;
array[8573] <= 16'b0000_0000_0000_0000;
array[8574] <= 16'b0000_0000_0000_0000;
array[8575] <= 16'b0000_0000_0000_0000;
array[8576] <= 16'b0000_0000_0000_0000;
array[8577] <= 16'b0000_0000_0000_0000;
array[8578] <= 16'b0000_0000_0000_0000;
array[8579] <= 16'b0000_0000_0000_0000;
array[8580] <= 16'b0000_0000_0000_0000;
array[8581] <= 16'b0000_0000_0000_0000;
array[8582] <= 16'b0000_0000_0000_0000;
array[8583] <= 16'b0000_0000_0000_0000;
array[8584] <= 16'b0000_0000_0000_0000;
array[8585] <= 16'b0000_0000_0000_0000;
array[8586] <= 16'b0000_0000_0000_0000;
array[8587] <= 16'b0000_0000_0000_0000;
array[8588] <= 16'b0000_0000_0000_0000;
array[8589] <= 16'b0000_0000_0000_0000;
array[8590] <= 16'b0000_0000_0000_0000;
array[8591] <= 16'b0000_0000_0000_0000;
array[8592] <= 16'b0000_0000_0000_0000;
array[8593] <= 16'b0000_0000_0000_0000;
array[8594] <= 16'b0000_0000_0000_0000;
array[8595] <= 16'b0000_0000_0000_0000;
array[8596] <= 16'b0000_0000_0000_0000;
array[8597] <= 16'b0000_0000_0000_0000;
array[8598] <= 16'b0000_0000_0000_0000;
array[8599] <= 16'b0000_0000_0000_0000;
array[8600] <= 16'b0000_0000_0000_0000;
array[8601] <= 16'b0000_0000_0000_0000;
array[8602] <= 16'b0000_0000_0000_0000;
array[8603] <= 16'b0000_0000_0000_0000;
array[8604] <= 16'b0000_0000_0000_0000;
array[8605] <= 16'b0000_0000_0000_0000;
array[8606] <= 16'b0000_0000_0000_0000;
array[8607] <= 16'b0000_0000_0000_0000;
array[8608] <= 16'b0000_0000_0000_0000;
array[8609] <= 16'b0000_0000_0000_0000;
array[8610] <= 16'b0000_0000_0000_0000;
array[8611] <= 16'b0000_0000_0000_0000;
array[8612] <= 16'b0000_0000_0000_0000;
array[8613] <= 16'b0000_0000_0000_0000;
array[8614] <= 16'b0000_0000_0000_0000;
array[8615] <= 16'b0000_0000_0000_0000;
array[8616] <= 16'b0000_0000_0000_0000;
array[8617] <= 16'b0000_0000_0000_0000;
array[8618] <= 16'b0000_0000_0000_0000;
array[8619] <= 16'b0000_0000_0000_0000;
array[8620] <= 16'b0000_0000_0000_0000;
array[8621] <= 16'b0000_0000_0000_0000;
array[8622] <= 16'b0000_0000_0000_0000;
array[8623] <= 16'b0000_0000_0000_0000;
array[8624] <= 16'b0000_0000_0000_0000;
array[8625] <= 16'b0000_0000_0000_0000;
array[8626] <= 16'b0000_0000_0000_0000;
array[8627] <= 16'b0000_0000_0000_0000;
array[8628] <= 16'b0000_0000_0000_0000;
array[8629] <= 16'b0000_0000_0000_0000;
array[8630] <= 16'b0000_0000_0000_0000;
array[8631] <= 16'b0000_0000_0000_0000;
array[8632] <= 16'b0000_0000_0000_0000;
array[8633] <= 16'b0000_0000_0000_0000;
array[8634] <= 16'b0000_0000_0000_0000;
array[8635] <= 16'b0000_0000_0000_0000;
array[8636] <= 16'b0000_0000_0000_0000;
array[8637] <= 16'b0000_0000_0000_0000;
array[8638] <= 16'b0000_0000_0000_0000;
array[8639] <= 16'b0000_0000_0000_0000;
array[8640] <= 16'b0000_0000_0000_0000;
array[8641] <= 16'b0000_0000_0000_0000;
array[8642] <= 16'b0000_0000_0000_0000;
array[8643] <= 16'b0000_0000_0000_0000;
array[8644] <= 16'b0000_0000_0000_0000;
array[8645] <= 16'b0000_0000_0000_0000;
array[8646] <= 16'b0000_0000_0000_0000;
array[8647] <= 16'b0000_0000_0000_0000;
array[8648] <= 16'b0000_0000_0000_0000;
array[8649] <= 16'b0000_0000_0000_0000;
array[8650] <= 16'b0000_0000_0000_0000;
array[8651] <= 16'b0000_0000_0000_0000;
array[8652] <= 16'b0000_0000_0000_0000;
array[8653] <= 16'b0000_0000_0000_0000;
array[8654] <= 16'b0000_0000_0000_0000;
array[8655] <= 16'b0000_0000_0000_0000;
array[8656] <= 16'b0000_0000_0000_0000;
array[8657] <= 16'b0000_0000_0000_0000;
array[8658] <= 16'b0000_0000_0000_0000;
array[8659] <= 16'b0000_0000_0000_0000;
array[8660] <= 16'b0000_0000_0000_0000;
array[8661] <= 16'b0000_0000_0000_0000;
array[8662] <= 16'b0000_0000_0000_0000;
array[8663] <= 16'b0000_0000_0000_0000;
array[8664] <= 16'b0000_0000_0000_0000;
array[8665] <= 16'b0000_0000_0000_0000;
array[8666] <= 16'b0000_0000_0000_0000;
array[8667] <= 16'b0000_0000_0000_0000;
array[8668] <= 16'b0000_0000_0000_0000;
array[8669] <= 16'b0000_0000_0000_0000;
array[8670] <= 16'b0000_0000_0000_0000;
array[8671] <= 16'b0000_0000_0000_0000;
array[8672] <= 16'b0000_0000_0000_0000;
array[8673] <= 16'b0000_0000_0000_0000;
array[8674] <= 16'b0000_0000_0000_0000;
array[8675] <= 16'b0000_0000_0000_0000;
array[8676] <= 16'b0000_0000_0000_0000;
array[8677] <= 16'b0000_0000_0000_0000;
array[8678] <= 16'b0000_0000_0000_0000;
array[8679] <= 16'b0000_0000_0000_0000;
array[8680] <= 16'b0000_0000_0000_0000;
array[8681] <= 16'b0000_0000_0000_0000;
array[8682] <= 16'b0000_0000_0000_0000;
array[8683] <= 16'b0000_0000_0000_0000;
array[8684] <= 16'b0000_0000_0000_0000;
array[8685] <= 16'b0000_0000_0000_0000;
array[8686] <= 16'b0000_0000_0000_0000;
array[8687] <= 16'b0000_0000_0000_0000;
array[8688] <= 16'b0000_0000_0000_0000;
array[8689] <= 16'b0000_0000_0000_0000;
array[8690] <= 16'b0000_0000_0000_0000;
array[8691] <= 16'b0000_0000_0000_0000;
array[8692] <= 16'b0000_0000_0000_0000;
array[8693] <= 16'b0000_0000_0000_0000;
array[8694] <= 16'b0000_0000_0000_0000;
array[8695] <= 16'b0000_0000_0000_0000;
array[8696] <= 16'b0000_0000_0000_0000;
array[8697] <= 16'b0000_0000_0000_0000;
array[8698] <= 16'b0000_0000_0000_0000;
array[8699] <= 16'b0000_0000_0000_0000;
array[8700] <= 16'b0000_0000_0000_0000;
array[8701] <= 16'b0000_0000_0000_0000;
array[8702] <= 16'b0000_0000_0000_0000;
array[8703] <= 16'b0000_0000_0000_0000;
array[8704] <= 16'b0000_0000_0000_0000;
array[8705] <= 16'b0000_0000_0000_0000;
array[8706] <= 16'b0000_0000_0000_0000;
array[8707] <= 16'b0000_0000_0000_0000;
array[8708] <= 16'b0000_0000_0000_0000;
array[8709] <= 16'b0000_0000_0000_0000;
array[8710] <= 16'b0000_0000_0000_0000;
array[8711] <= 16'b0000_0000_0000_0000;
array[8712] <= 16'b0000_0000_0000_0000;
array[8713] <= 16'b0000_0000_0000_0000;
array[8714] <= 16'b0000_0000_0000_0000;
array[8715] <= 16'b0000_0000_0000_0000;
array[8716] <= 16'b0000_0000_0000_0000;
array[8717] <= 16'b0000_0000_0000_0000;
array[8718] <= 16'b0000_0000_0000_0000;
array[8719] <= 16'b0000_0000_0000_0000;
array[8720] <= 16'b0000_0000_0000_0000;
array[8721] <= 16'b0000_0000_0000_0000;
array[8722] <= 16'b0000_0000_0000_0000;
array[8723] <= 16'b0000_0000_0000_0000;
array[8724] <= 16'b0000_0000_0000_0000;
array[8725] <= 16'b0000_0000_0000_0000;
array[8726] <= 16'b0000_0000_0000_0000;
array[8727] <= 16'b0000_0000_0000_0000;
array[8728] <= 16'b0000_0000_0000_0000;
array[8729] <= 16'b0000_0000_0000_0000;
array[8730] <= 16'b0000_0000_0000_0000;
array[8731] <= 16'b0000_0000_0000_0000;
array[8732] <= 16'b0000_0000_0000_0000;
array[8733] <= 16'b0000_0000_0000_0000;
array[8734] <= 16'b0000_0000_0000_0000;
array[8735] <= 16'b0000_0000_0000_0000;
array[8736] <= 16'b0000_0000_0000_0000;
array[8737] <= 16'b0000_0000_0000_0000;
array[8738] <= 16'b0000_0000_0000_0000;
array[8739] <= 16'b0000_0000_0000_0000;
array[8740] <= 16'b0000_0000_0000_0000;
array[8741] <= 16'b0000_0000_0000_0000;
array[8742] <= 16'b0000_0000_0000_0000;
array[8743] <= 16'b0000_0000_0000_0000;
array[8744] <= 16'b0000_0000_0000_0000;
array[8745] <= 16'b0000_0000_0000_0000;
array[8746] <= 16'b0000_0000_0000_0000;
array[8747] <= 16'b0000_0000_0000_0000;
array[8748] <= 16'b0000_0000_0000_0000;
array[8749] <= 16'b0000_0000_0000_0000;
array[8750] <= 16'b0000_0000_0000_0000;
array[8751] <= 16'b0000_0000_0000_0000;
array[8752] <= 16'b0000_0000_0000_0000;
array[8753] <= 16'b0000_0000_0000_0000;
array[8754] <= 16'b0000_0000_0000_0000;
array[8755] <= 16'b0000_0000_0000_0000;
array[8756] <= 16'b0000_0000_0000_0000;
array[8757] <= 16'b0000_0000_0000_0000;
array[8758] <= 16'b0000_0000_0000_0000;
array[8759] <= 16'b0000_0000_0000_0000;
array[8760] <= 16'b0000_0000_0000_0000;
array[8761] <= 16'b0000_0000_0000_0000;
array[8762] <= 16'b0000_0000_0000_0000;
array[8763] <= 16'b0000_0000_0000_0000;
array[8764] <= 16'b0000_0000_0000_0000;
array[8765] <= 16'b0000_0000_0000_0000;
array[8766] <= 16'b0000_0000_0000_0000;
array[8767] <= 16'b0000_0000_0000_0000;
array[8768] <= 16'b0000_0000_0000_0000;
array[8769] <= 16'b0000_0000_0000_0000;
array[8770] <= 16'b0000_0000_0000_0000;
array[8771] <= 16'b0000_0000_0000_0000;
array[8772] <= 16'b0000_0000_0000_0000;
array[8773] <= 16'b0000_0000_0000_0000;
array[8774] <= 16'b0000_0000_0000_0000;
array[8775] <= 16'b0000_0000_0000_0000;
array[8776] <= 16'b0000_0000_0000_0000;
array[8777] <= 16'b0000_0000_0000_0000;
array[8778] <= 16'b0000_0000_0000_0000;
array[8779] <= 16'b0000_0000_0000_0000;
array[8780] <= 16'b0000_0000_0000_0000;
array[8781] <= 16'b0000_0000_0000_0000;
array[8782] <= 16'b0000_0000_0000_0000;
array[8783] <= 16'b0000_0000_0000_0000;
array[8784] <= 16'b0000_0000_0000_0000;
array[8785] <= 16'b0000_0000_0000_0000;
array[8786] <= 16'b0000_0000_0000_0000;
array[8787] <= 16'b0000_0000_0000_0000;
array[8788] <= 16'b0000_0000_0000_0000;
array[8789] <= 16'b0000_0000_0000_0000;
array[8790] <= 16'b0000_0000_0000_0000;
array[8791] <= 16'b0000_0000_0000_0000;
array[8792] <= 16'b0000_0000_0000_0000;
array[8793] <= 16'b0000_0000_0000_0000;
array[8794] <= 16'b0000_0000_0000_0000;
array[8795] <= 16'b0000_0000_0000_0000;
array[8796] <= 16'b0000_0000_0000_0000;
array[8797] <= 16'b0000_0000_0000_0000;
array[8798] <= 16'b0000_0000_0000_0000;
array[8799] <= 16'b0000_0000_0000_0000;
array[8800] <= 16'b0000_0000_0000_0000;
array[8801] <= 16'b0000_0000_0000_0000;
array[8802] <= 16'b0000_0000_0000_0000;
array[8803] <= 16'b0000_0000_0000_0000;
array[8804] <= 16'b0000_0000_0000_0000;
array[8805] <= 16'b0000_0000_0000_0000;
array[8806] <= 16'b0000_0000_0000_0000;
array[8807] <= 16'b0000_0000_0000_0000;
array[8808] <= 16'b0000_0000_0000_0000;
array[8809] <= 16'b0000_0000_0000_0000;
array[8810] <= 16'b0000_0000_0000_0000;
array[8811] <= 16'b0000_0000_0000_0000;
array[8812] <= 16'b0000_0000_0000_0000;
array[8813] <= 16'b0000_0000_0000_0000;
array[8814] <= 16'b0000_0000_0000_0000;
array[8815] <= 16'b0000_0000_0000_0000;
array[8816] <= 16'b0000_0000_0000_0000;
array[8817] <= 16'b0000_0000_0000_0000;
array[8818] <= 16'b0000_0000_0000_0000;
array[8819] <= 16'b0000_0000_0000_0000;
array[8820] <= 16'b0000_0000_0000_0000;
array[8821] <= 16'b0000_0000_0000_0000;
array[8822] <= 16'b0000_0000_0000_0000;
array[8823] <= 16'b0000_0000_0000_0000;
array[8824] <= 16'b0000_0000_0000_0000;
array[8825] <= 16'b0000_0000_0000_0000;
array[8826] <= 16'b0000_0000_0000_0000;
array[8827] <= 16'b0000_0000_0000_0000;
array[8828] <= 16'b0000_0000_0000_0000;
array[8829] <= 16'b0000_0000_0000_0000;
array[8830] <= 16'b0000_0000_0000_0000;
array[8831] <= 16'b0000_0000_0000_0000;
array[8832] <= 16'b0000_0000_0000_0000;
array[8833] <= 16'b0000_0000_0000_0000;
array[8834] <= 16'b0000_0000_0000_0000;
array[8835] <= 16'b0000_0000_0000_0000;
array[8836] <= 16'b0000_0000_0000_0000;
array[8837] <= 16'b0000_0000_0000_0000;
array[8838] <= 16'b0000_0000_0000_0000;
array[8839] <= 16'b0000_0000_0000_0000;
array[8840] <= 16'b0000_0000_0000_0000;
array[8841] <= 16'b0000_0000_0000_0000;
array[8842] <= 16'b0000_0000_0000_0000;
array[8843] <= 16'b0000_0000_0000_0000;
array[8844] <= 16'b0000_0000_0000_0000;
array[8845] <= 16'b0000_0000_0000_0000;
array[8846] <= 16'b0000_0000_0000_0000;
array[8847] <= 16'b0000_0000_0000_0000;
array[8848] <= 16'b0000_0000_0000_0000;
array[8849] <= 16'b0000_0000_0000_0000;
array[8850] <= 16'b0000_0000_0000_0000;
array[8851] <= 16'b0000_0000_0000_0000;
array[8852] <= 16'b0000_0000_0000_0000;
array[8853] <= 16'b0000_0000_0000_0000;
array[8854] <= 16'b0000_0000_0000_0000;
array[8855] <= 16'b0000_0000_0000_0000;
array[8856] <= 16'b0000_0000_0000_0000;
array[8857] <= 16'b0000_0000_0000_0000;
array[8858] <= 16'b0000_0000_0000_0000;
array[8859] <= 16'b0000_0000_0000_0000;
array[8860] <= 16'b0000_0000_0000_0000;
array[8861] <= 16'b0000_0000_0000_0000;
array[8862] <= 16'b0000_0000_0000_0000;
array[8863] <= 16'b0000_0000_0000_0000;
array[8864] <= 16'b0000_0000_0000_0000;
array[8865] <= 16'b0000_0000_0000_0000;
array[8866] <= 16'b0000_0000_0000_0000;
array[8867] <= 16'b0000_0000_0000_0000;
array[8868] <= 16'b0000_0000_0000_0000;
array[8869] <= 16'b0000_0000_0000_0000;
array[8870] <= 16'b0000_0000_0000_0000;
array[8871] <= 16'b0000_0000_0000_0000;
array[8872] <= 16'b0000_0000_0000_0000;
array[8873] <= 16'b0000_0000_0000_0000;
array[8874] <= 16'b0000_0000_0000_0000;
array[8875] <= 16'b0000_0000_0000_0000;
array[8876] <= 16'b0000_0000_0000_0000;
array[8877] <= 16'b0000_0000_0000_0000;
array[8878] <= 16'b0000_0000_0000_0000;
array[8879] <= 16'b0000_0000_0000_0000;
array[8880] <= 16'b0000_0000_0000_0000;
array[8881] <= 16'b0000_0000_0000_0000;
array[8882] <= 16'b0000_0000_0000_0000;
array[8883] <= 16'b0000_0000_0000_0000;
array[8884] <= 16'b0000_0000_0000_0000;
array[8885] <= 16'b0000_0000_0000_0000;
array[8886] <= 16'b0000_0000_0000_0000;
array[8887] <= 16'b0000_0000_0000_0000;
array[8888] <= 16'b0000_0000_0000_0000;
array[8889] <= 16'b0000_0000_0000_0000;
array[8890] <= 16'b0000_0000_0000_0000;
array[8891] <= 16'b0000_0000_0000_0000;
array[8892] <= 16'b0000_0000_0000_0000;
array[8893] <= 16'b0000_0000_0000_0000;
array[8894] <= 16'b0000_0000_0000_0000;
array[8895] <= 16'b0000_0000_0000_0000;
array[8896] <= 16'b0000_0000_0000_0000;
array[8897] <= 16'b0000_0000_0000_0000;
array[8898] <= 16'b0000_0000_0000_0000;
array[8899] <= 16'b0000_0000_0000_0000;
array[8900] <= 16'b0000_0000_0000_0000;
array[8901] <= 16'b0000_0000_0000_0000;
array[8902] <= 16'b0000_0000_0000_0000;
array[8903] <= 16'b0000_0000_0000_0000;
array[8904] <= 16'b0000_0000_0000_0000;
array[8905] <= 16'b0000_0000_0000_0000;
array[8906] <= 16'b0000_0000_0000_0000;
array[8907] <= 16'b0000_0000_0000_0000;
array[8908] <= 16'b0000_0000_0000_0000;
array[8909] <= 16'b0000_0000_0000_0000;
array[8910] <= 16'b0000_0000_0000_0000;
array[8911] <= 16'b0000_0000_0000_0000;
array[8912] <= 16'b0000_0000_0000_0000;
array[8913] <= 16'b0000_0000_0000_0000;
array[8914] <= 16'b0000_0000_0000_0000;
array[8915] <= 16'b0000_0000_0000_0000;
array[8916] <= 16'b0000_0000_0000_0000;
array[8917] <= 16'b0000_0000_0000_0000;
array[8918] <= 16'b0000_0000_0000_0000;
array[8919] <= 16'b0000_0000_0000_0000;
array[8920] <= 16'b0000_0000_0000_0000;
array[8921] <= 16'b0000_0000_0000_0000;
array[8922] <= 16'b0000_0000_0000_0000;
array[8923] <= 16'b0000_0000_0000_0000;
array[8924] <= 16'b0000_0000_0000_0000;
array[8925] <= 16'b0000_0000_0000_0000;
array[8926] <= 16'b0000_0000_0000_0000;
array[8927] <= 16'b0000_0000_0000_0000;
array[8928] <= 16'b0000_0000_0000_0000;
array[8929] <= 16'b0000_0000_0000_0000;
array[8930] <= 16'b0000_0000_0000_0000;
array[8931] <= 16'b0000_0000_0000_0000;
array[8932] <= 16'b0000_0000_0000_0000;
array[8933] <= 16'b0000_0000_0000_0000;
array[8934] <= 16'b0000_0000_0000_0000;
array[8935] <= 16'b0000_0000_0000_0000;
array[8936] <= 16'b0000_0000_0000_0000;
array[8937] <= 16'b0000_0000_0000_0000;
array[8938] <= 16'b0000_0000_0000_0000;
array[8939] <= 16'b0000_0000_0000_0000;
array[8940] <= 16'b0000_0000_0000_0000;
array[8941] <= 16'b0000_0000_0000_0000;
array[8942] <= 16'b0000_0000_0000_0000;
array[8943] <= 16'b0000_0000_0000_0000;
array[8944] <= 16'b0000_0000_0000_0000;
array[8945] <= 16'b0000_0000_0000_0000;
array[8946] <= 16'b0000_0000_0000_0000;
array[8947] <= 16'b0000_0000_0000_0000;
array[8948] <= 16'b0000_0000_0000_0000;
array[8949] <= 16'b0000_0000_0000_0000;
array[8950] <= 16'b0000_0000_0000_0000;
array[8951] <= 16'b0000_0000_0000_0000;
array[8952] <= 16'b0000_0000_0000_0000;
array[8953] <= 16'b0000_0000_0000_0000;
array[8954] <= 16'b0000_0000_0000_0000;
array[8955] <= 16'b0000_0000_0000_0000;
array[8956] <= 16'b0000_0000_0000_0000;
array[8957] <= 16'b0000_0000_0000_0000;
array[8958] <= 16'b0000_0000_0000_0000;
array[8959] <= 16'b0000_0000_0000_0000;
array[8960] <= 16'b0000_0000_0000_0000;
array[8961] <= 16'b0000_0000_0000_0000;
array[8962] <= 16'b0000_0000_0000_0000;
array[8963] <= 16'b0000_0000_0000_0000;
array[8964] <= 16'b0000_0000_0000_0000;
array[8965] <= 16'b0000_0000_0000_0000;
array[8966] <= 16'b0000_0000_0000_0000;
array[8967] <= 16'b0000_0000_0000_0000;
array[8968] <= 16'b0000_0000_0000_0000;
array[8969] <= 16'b0000_0000_0000_0000;
array[8970] <= 16'b0000_0000_0000_0000;
array[8971] <= 16'b0000_0000_0000_0000;
array[8972] <= 16'b0000_0000_0000_0000;
array[8973] <= 16'b0000_0000_0000_0000;
array[8974] <= 16'b0000_0000_0000_0000;
array[8975] <= 16'b0000_0000_0000_0000;
array[8976] <= 16'b0000_0000_0000_0000;
array[8977] <= 16'b0000_0000_0000_0000;
array[8978] <= 16'b0000_0000_0000_0000;
array[8979] <= 16'b0000_0000_0000_0000;
array[8980] <= 16'b0000_0000_0000_0000;
array[8981] <= 16'b0000_0000_0000_0000;
array[8982] <= 16'b0000_0000_0000_0000;
array[8983] <= 16'b0000_0000_0000_0000;
array[8984] <= 16'b0000_0000_0000_0000;
array[8985] <= 16'b0000_0000_0000_0000;
array[8986] <= 16'b0000_0000_0000_0000;
array[8987] <= 16'b0000_0000_0000_0000;
array[8988] <= 16'b0000_0000_0000_0000;
array[8989] <= 16'b0000_0000_0000_0000;
array[8990] <= 16'b0000_0000_0000_0000;
array[8991] <= 16'b0000_0000_0000_0000;
array[8992] <= 16'b0000_0000_0000_0000;
array[8993] <= 16'b0000_0000_0000_0000;
array[8994] <= 16'b0000_0000_0000_0000;
array[8995] <= 16'b0000_0000_0000_0000;
array[8996] <= 16'b0000_0000_0000_0000;
array[8997] <= 16'b0000_0000_0000_0000;
array[8998] <= 16'b0000_0000_0000_0000;
array[8999] <= 16'b0000_0000_0000_0000;
array[9000] <= 16'b0000_0000_0000_0000;
array[9001] <= 16'b0000_0000_0000_0000;
array[9002] <= 16'b0000_0000_0000_0000;
array[9003] <= 16'b0000_0000_0000_0000;
array[9004] <= 16'b0000_0000_0000_0000;
array[9005] <= 16'b0000_0000_0000_0000;
array[9006] <= 16'b0000_0000_0000_0000;
array[9007] <= 16'b0000_0000_0000_0000;
array[9008] <= 16'b0000_0000_0000_0000;
array[9009] <= 16'b0000_0000_0000_0000;
array[9010] <= 16'b0000_0000_0000_0000;
array[9011] <= 16'b0000_0000_0000_0000;
array[9012] <= 16'b0000_0000_0000_0000;
array[9013] <= 16'b0000_0000_0000_0000;
array[9014] <= 16'b0000_0000_0000_0000;
array[9015] <= 16'b0000_0000_0000_0000;
array[9016] <= 16'b0000_0000_0000_0000;
array[9017] <= 16'b0000_0000_0000_0000;
array[9018] <= 16'b0000_0000_0000_0000;
array[9019] <= 16'b0000_0000_0000_0000;
array[9020] <= 16'b0000_0000_0000_0000;
array[9021] <= 16'b0000_0000_0000_0000;
array[9022] <= 16'b0000_0000_0000_0000;
array[9023] <= 16'b0000_0000_0000_0000;
array[9024] <= 16'b0000_0000_0000_0000;
array[9025] <= 16'b0000_0000_0000_0000;
array[9026] <= 16'b0000_0000_0000_0000;
array[9027] <= 16'b0000_0000_0000_0000;
array[9028] <= 16'b0000_0000_0000_0000;
array[9029] <= 16'b0000_0000_0000_0000;
array[9030] <= 16'b0000_0000_0000_0000;
array[9031] <= 16'b0000_0000_0000_0000;
array[9032] <= 16'b0000_0000_0000_0000;
array[9033] <= 16'b0000_0000_0000_0000;
array[9034] <= 16'b0000_0000_0000_0000;
array[9035] <= 16'b0000_0000_0000_0000;
array[9036] <= 16'b0000_0000_0000_0000;
array[9037] <= 16'b0000_0000_0000_0000;
array[9038] <= 16'b0000_0000_0000_0000;
array[9039] <= 16'b0000_0000_0000_0000;
array[9040] <= 16'b0000_0000_0000_0000;
array[9041] <= 16'b0000_0000_0000_0000;
array[9042] <= 16'b0000_0000_0000_0000;
array[9043] <= 16'b0000_0000_0000_0000;
array[9044] <= 16'b0000_0000_0000_0000;
array[9045] <= 16'b0000_0000_0000_0000;
array[9046] <= 16'b0000_0000_0000_0000;
array[9047] <= 16'b0000_0000_0000_0000;
array[9048] <= 16'b0000_0000_0000_0000;
array[9049] <= 16'b0000_0000_0000_0000;
array[9050] <= 16'b0000_0000_0000_0000;
array[9051] <= 16'b0000_0000_0000_0000;
array[9052] <= 16'b0000_0000_0000_0000;
array[9053] <= 16'b0000_0000_0000_0000;
array[9054] <= 16'b0000_0000_0000_0000;
array[9055] <= 16'b0000_0000_0000_0000;
array[9056] <= 16'b0000_0000_0000_0000;
array[9057] <= 16'b0000_0000_0000_0000;
array[9058] <= 16'b0000_0000_0000_0000;
array[9059] <= 16'b0000_0000_0000_0000;
array[9060] <= 16'b0000_0000_0000_0000;
array[9061] <= 16'b0000_0000_0000_0000;
array[9062] <= 16'b0000_0000_0000_0000;
array[9063] <= 16'b0000_0000_0000_0000;
array[9064] <= 16'b0000_0000_0000_0000;
array[9065] <= 16'b0000_0000_0000_0000;
array[9066] <= 16'b0000_0000_0000_0000;
array[9067] <= 16'b0000_0000_0000_0000;
array[9068] <= 16'b0000_0000_0000_0000;
array[9069] <= 16'b0000_0000_0000_0000;
array[9070] <= 16'b0000_0000_0000_0000;
array[9071] <= 16'b0000_0000_0000_0000;
array[9072] <= 16'b0000_0000_0000_0000;
array[9073] <= 16'b0000_0000_0000_0000;
array[9074] <= 16'b0000_0000_0000_0000;
array[9075] <= 16'b0000_0000_0000_0000;
array[9076] <= 16'b0000_0000_0000_0000;
array[9077] <= 16'b0000_0000_0000_0000;
array[9078] <= 16'b0000_0000_0000_0000;
array[9079] <= 16'b0000_0000_0000_0000;
array[9080] <= 16'b0000_0000_0000_0000;
array[9081] <= 16'b0000_0000_0000_0000;
array[9082] <= 16'b0000_0000_0000_0000;
array[9083] <= 16'b0000_0000_0000_0000;
array[9084] <= 16'b0000_0000_0000_0000;
array[9085] <= 16'b0000_0000_0000_0000;
array[9086] <= 16'b0000_0000_0000_0000;
array[9087] <= 16'b0000_0000_0000_0000;
array[9088] <= 16'b0000_0000_0000_0000;
array[9089] <= 16'b0000_0000_0000_0000;
array[9090] <= 16'b0000_0000_0000_0000;
array[9091] <= 16'b0000_0000_0000_0000;
array[9092] <= 16'b0000_0000_0000_0000;
array[9093] <= 16'b0000_0000_0000_0000;
array[9094] <= 16'b0000_0000_0000_0000;
array[9095] <= 16'b0000_0000_0000_0000;
array[9096] <= 16'b0000_0000_0000_0000;
array[9097] <= 16'b0000_0000_0000_0000;
array[9098] <= 16'b0000_0000_0000_0000;
array[9099] <= 16'b0000_0000_0000_0000;
array[9100] <= 16'b0000_0000_0000_0000;
array[9101] <= 16'b0000_0000_0000_0000;
array[9102] <= 16'b0000_0000_0000_0000;
array[9103] <= 16'b0000_0000_0000_0000;
array[9104] <= 16'b0000_0000_0000_0000;
array[9105] <= 16'b0000_0000_0000_0000;
array[9106] <= 16'b0000_0000_0000_0000;
array[9107] <= 16'b0000_0000_0000_0000;
array[9108] <= 16'b0000_0000_0000_0000;
array[9109] <= 16'b0000_0000_0000_0000;
array[9110] <= 16'b0000_0000_0000_0000;
array[9111] <= 16'b0000_0000_0000_0000;
array[9112] <= 16'b0000_0000_0000_0000;
array[9113] <= 16'b0000_0000_0000_0000;
array[9114] <= 16'b0000_0000_0000_0000;
array[9115] <= 16'b0000_0000_0000_0000;
array[9116] <= 16'b0000_0000_0000_0000;
array[9117] <= 16'b0000_0000_0000_0000;
array[9118] <= 16'b0000_0000_0000_0000;
array[9119] <= 16'b0000_0000_0000_0000;
array[9120] <= 16'b0000_0000_0000_0000;
array[9121] <= 16'b0000_0000_0000_0000;
array[9122] <= 16'b0000_0000_0000_0000;
array[9123] <= 16'b0000_0000_0000_0000;
array[9124] <= 16'b0000_0000_0000_0000;
array[9125] <= 16'b0000_0000_0000_0000;
array[9126] <= 16'b0000_0000_0000_0000;
array[9127] <= 16'b0000_0000_0000_0000;
array[9128] <= 16'b0000_0000_0000_0000;
array[9129] <= 16'b0000_0000_0000_0000;
array[9130] <= 16'b0000_0000_0000_0000;
array[9131] <= 16'b0000_0000_0000_0000;
array[9132] <= 16'b0000_0000_0000_0000;
array[9133] <= 16'b0000_0000_0000_0000;
array[9134] <= 16'b0000_0000_0000_0000;
array[9135] <= 16'b0000_0000_0000_0000;
array[9136] <= 16'b0000_0000_0000_0000;
array[9137] <= 16'b0000_0000_0000_0000;
array[9138] <= 16'b0000_0000_0000_0000;
array[9139] <= 16'b0000_0000_0000_0000;
array[9140] <= 16'b0000_0000_0000_0000;
array[9141] <= 16'b0000_0000_0000_0000;
array[9142] <= 16'b0000_0000_0000_0000;
array[9143] <= 16'b0000_0000_0000_0000;
array[9144] <= 16'b0000_0000_0000_0000;
array[9145] <= 16'b0000_0000_0000_0000;
array[9146] <= 16'b0000_0000_0000_0000;
array[9147] <= 16'b0000_0000_0000_0000;
array[9148] <= 16'b0000_0000_0000_0000;
array[9149] <= 16'b0000_0000_0000_0000;
array[9150] <= 16'b0000_0000_0000_0000;
array[9151] <= 16'b0000_0000_0000_0000;
array[9152] <= 16'b0000_0000_0000_0000;
array[9153] <= 16'b0000_0000_0000_0000;
array[9154] <= 16'b0000_0000_0000_0000;
array[9155] <= 16'b0000_0000_0000_0000;
array[9156] <= 16'b0000_0000_0000_0000;
array[9157] <= 16'b0000_0000_0000_0000;
array[9158] <= 16'b0000_0000_0000_0000;
array[9159] <= 16'b0000_0000_0000_0000;
array[9160] <= 16'b0000_0000_0000_0000;
array[9161] <= 16'b0000_0000_0000_0000;
array[9162] <= 16'b0000_0000_0000_0000;
array[9163] <= 16'b0000_0000_0000_0000;
array[9164] <= 16'b0000_0000_0000_0000;
array[9165] <= 16'b0000_0000_0000_0000;
array[9166] <= 16'b0000_0000_0000_0000;
array[9167] <= 16'b0000_0000_0000_0000;
array[9168] <= 16'b0000_0000_0000_0000;
array[9169] <= 16'b0000_0000_0000_0000;
array[9170] <= 16'b0000_0000_0000_0000;
array[9171] <= 16'b0000_0000_0000_0000;
array[9172] <= 16'b0000_0000_0000_0000;
array[9173] <= 16'b0000_0000_0000_0000;
array[9174] <= 16'b0000_0000_0000_0000;
array[9175] <= 16'b0000_0000_0000_0000;
array[9176] <= 16'b0000_0000_0000_0000;
array[9177] <= 16'b0000_0000_0000_0000;
array[9178] <= 16'b0000_0000_0000_0000;
array[9179] <= 16'b0000_0000_0000_0000;
array[9180] <= 16'b0000_0000_0000_0000;
array[9181] <= 16'b0000_0000_0000_0000;
array[9182] <= 16'b0000_0000_0000_0000;
array[9183] <= 16'b0000_0000_0000_0000;
array[9184] <= 16'b0000_0000_0000_0000;
array[9185] <= 16'b0000_0000_0000_0000;
array[9186] <= 16'b0000_0000_0000_0000;
array[9187] <= 16'b0000_0000_0000_0000;
array[9188] <= 16'b0000_0000_0000_0000;
array[9189] <= 16'b0000_0000_0000_0000;
array[9190] <= 16'b0000_0000_0000_0000;
array[9191] <= 16'b0000_0000_0000_0000;
array[9192] <= 16'b0000_0000_0000_0000;
array[9193] <= 16'b0000_0000_0000_0000;
array[9194] <= 16'b0000_0000_0000_0000;
array[9195] <= 16'b0000_0000_0000_0000;
array[9196] <= 16'b0000_0000_0000_0000;
array[9197] <= 16'b0000_0000_0000_0000;
array[9198] <= 16'b0000_0000_0000_0000;
array[9199] <= 16'b0000_0000_0000_0000;
array[9200] <= 16'b0000_0000_0000_0000;
array[9201] <= 16'b0000_0000_0000_0000;
array[9202] <= 16'b0000_0000_0000_0000;
array[9203] <= 16'b0000_0000_0000_0000;
array[9204] <= 16'b0000_0000_0000_0000;
array[9205] <= 16'b0000_0000_0000_0000;
array[9206] <= 16'b0000_0000_0000_0000;
array[9207] <= 16'b0000_0000_0000_0000;
array[9208] <= 16'b0000_0000_0000_0000;
array[9209] <= 16'b0000_0000_0000_0000;
array[9210] <= 16'b0000_0000_0000_0000;
array[9211] <= 16'b0000_0000_0000_0000;
array[9212] <= 16'b0000_0000_0000_0000;
array[9213] <= 16'b0000_0000_0000_0000;
array[9214] <= 16'b0000_0000_0000_0000;
array[9215] <= 16'b0000_0000_0000_0000;
array[9216] <= 16'b0000_0000_0000_0000;
array[9217] <= 16'b0000_0000_0000_0000;
array[9218] <= 16'b0000_0000_0000_0000;
array[9219] <= 16'b0000_0000_0000_0000;
array[9220] <= 16'b0000_0000_0000_0000;
array[9221] <= 16'b0000_0000_0000_0000;
array[9222] <= 16'b0000_0000_0000_0000;
array[9223] <= 16'b0000_0000_0000_0000;
array[9224] <= 16'b0000_0000_0000_0000;
array[9225] <= 16'b0000_0000_0000_0000;
array[9226] <= 16'b0000_0000_0000_0000;
array[9227] <= 16'b0000_0000_0000_0000;
array[9228] <= 16'b0000_0000_0000_0000;
array[9229] <= 16'b0000_0000_0000_0000;
array[9230] <= 16'b0000_0000_0000_0000;
array[9231] <= 16'b0000_0000_0000_0000;
array[9232] <= 16'b0000_0000_0000_0000;
array[9233] <= 16'b0000_0000_0000_0000;
array[9234] <= 16'b0000_0000_0000_0000;
array[9235] <= 16'b0000_0000_0000_0000;
array[9236] <= 16'b0000_0000_0000_0000;
array[9237] <= 16'b0000_0000_0000_0000;
array[9238] <= 16'b0000_0000_0000_0000;
array[9239] <= 16'b0000_0000_0000_0000;
array[9240] <= 16'b0000_0000_0000_0000;
array[9241] <= 16'b0000_0000_0000_0000;
array[9242] <= 16'b0000_0000_0000_0000;
array[9243] <= 16'b0000_0000_0000_0000;
array[9244] <= 16'b0000_0000_0000_0000;
array[9245] <= 16'b0000_0000_0000_0000;
array[9246] <= 16'b0000_0000_0000_0000;
array[9247] <= 16'b0000_0000_0000_0000;
array[9248] <= 16'b0000_0000_0000_0000;
array[9249] <= 16'b0000_0000_0000_0000;
array[9250] <= 16'b0000_0000_0000_0000;
array[9251] <= 16'b0000_0000_0000_0000;
array[9252] <= 16'b0000_0000_0000_0000;
array[9253] <= 16'b0000_0000_0000_0000;
array[9254] <= 16'b0000_0000_0000_0000;
array[9255] <= 16'b0000_0000_0000_0000;
array[9256] <= 16'b0000_0000_0000_0000;
array[9257] <= 16'b0000_0000_0000_0000;
array[9258] <= 16'b0000_0000_0000_0000;
array[9259] <= 16'b0000_0000_0000_0000;
array[9260] <= 16'b0000_0000_0000_0000;
array[9261] <= 16'b0000_0000_0000_0000;
array[9262] <= 16'b0000_0000_0000_0000;
array[9263] <= 16'b0000_0000_0000_0000;
array[9264] <= 16'b0000_0000_0000_0000;
array[9265] <= 16'b0000_0000_0000_0000;
array[9266] <= 16'b0000_0000_0000_0000;
array[9267] <= 16'b0000_0000_0000_0000;
array[9268] <= 16'b0000_0000_0000_0000;
array[9269] <= 16'b0000_0000_0000_0000;
array[9270] <= 16'b0000_0000_0000_0000;
array[9271] <= 16'b0000_0000_0000_0000;
array[9272] <= 16'b0000_0000_0000_0000;
array[9273] <= 16'b0000_0000_0000_0000;
array[9274] <= 16'b0000_0000_0000_0000;
array[9275] <= 16'b0000_0000_0000_0000;
array[9276] <= 16'b0000_0000_0000_0000;
array[9277] <= 16'b0000_0000_0000_0000;
array[9278] <= 16'b0000_0000_0000_0000;
array[9279] <= 16'b0000_0000_0000_0000;
array[9280] <= 16'b0000_0000_0000_0000;
array[9281] <= 16'b0000_0000_0000_0000;
array[9282] <= 16'b0000_0000_0000_0000;
array[9283] <= 16'b0000_0000_0000_0000;
array[9284] <= 16'b0000_0000_0000_0000;
array[9285] <= 16'b0000_0000_0000_0000;
array[9286] <= 16'b0000_0000_0000_0000;
array[9287] <= 16'b0000_0000_0000_0000;
array[9288] <= 16'b0000_0000_0000_0000;
array[9289] <= 16'b0000_0000_0000_0000;
array[9290] <= 16'b0000_0000_0000_0000;
array[9291] <= 16'b0000_0000_0000_0000;
array[9292] <= 16'b0000_0000_0000_0000;
array[9293] <= 16'b0000_0000_0000_0000;
array[9294] <= 16'b0000_0000_0000_0000;
array[9295] <= 16'b0000_0000_0000_0000;
array[9296] <= 16'b0000_0000_0000_0000;
array[9297] <= 16'b0000_0000_0000_0000;
array[9298] <= 16'b0000_0000_0000_0000;
array[9299] <= 16'b0000_0000_0000_0000;
array[9300] <= 16'b0000_0000_0000_0000;
array[9301] <= 16'b0000_0000_0000_0000;
array[9302] <= 16'b0000_0000_0000_0000;
array[9303] <= 16'b0000_0000_0000_0000;
array[9304] <= 16'b0000_0000_0000_0000;
array[9305] <= 16'b0000_0000_0000_0000;
array[9306] <= 16'b0000_0000_0000_0000;
array[9307] <= 16'b0000_0000_0000_0000;
array[9308] <= 16'b0000_0000_0000_0000;
array[9309] <= 16'b0000_0000_0000_0000;
array[9310] <= 16'b0000_0000_0000_0000;
array[9311] <= 16'b0000_0000_0000_0000;
array[9312] <= 16'b0000_0000_0000_0000;
array[9313] <= 16'b0000_0000_0000_0000;
array[9314] <= 16'b0000_0000_0000_0000;
array[9315] <= 16'b0000_0000_0000_0000;
array[9316] <= 16'b0000_0000_0000_0000;
array[9317] <= 16'b0000_0000_0000_0000;
array[9318] <= 16'b0000_0000_0000_0000;
array[9319] <= 16'b0000_0000_0000_0000;
array[9320] <= 16'b0000_0000_0000_0000;
array[9321] <= 16'b0000_0000_0000_0000;
array[9322] <= 16'b0000_0000_0000_0000;
array[9323] <= 16'b0000_0000_0000_0000;
array[9324] <= 16'b0000_0000_0000_0000;
array[9325] <= 16'b0000_0000_0000_0000;
array[9326] <= 16'b0000_0000_0000_0000;
array[9327] <= 16'b0000_0000_0000_0000;
array[9328] <= 16'b0000_0000_0000_0000;
array[9329] <= 16'b0000_0000_0000_0000;
array[9330] <= 16'b0000_0000_0000_0000;
array[9331] <= 16'b0000_0000_0000_0000;
array[9332] <= 16'b0000_0000_0000_0000;
array[9333] <= 16'b0000_0000_0000_0000;
array[9334] <= 16'b0000_0000_0000_0000;
array[9335] <= 16'b0000_0000_0000_0000;
array[9336] <= 16'b0000_0000_0000_0000;
array[9337] <= 16'b0000_0000_0000_0000;
array[9338] <= 16'b0000_0000_0000_0000;
array[9339] <= 16'b0000_0000_0000_0000;
array[9340] <= 16'b0000_0000_0000_0000;
array[9341] <= 16'b0000_0000_0000_0000;
array[9342] <= 16'b0000_0000_0000_0000;
array[9343] <= 16'b0000_0000_0000_0000;
array[9344] <= 16'b0000_0000_0000_0000;
array[9345] <= 16'b0000_0000_0000_0000;
array[9346] <= 16'b0000_0000_0000_0000;
array[9347] <= 16'b0000_0000_0000_0000;
array[9348] <= 16'b0000_0000_0000_0000;
array[9349] <= 16'b0000_0000_0000_0000;
array[9350] <= 16'b0000_0000_0000_0000;
array[9351] <= 16'b0000_0000_0000_0000;
array[9352] <= 16'b0000_0000_0000_0000;
array[9353] <= 16'b0000_0000_0000_0000;
array[9354] <= 16'b0000_0000_0000_0000;
array[9355] <= 16'b0000_0000_0000_0000;
array[9356] <= 16'b0000_0000_0000_0000;
array[9357] <= 16'b0000_0000_0000_0000;
array[9358] <= 16'b0000_0000_0000_0000;
array[9359] <= 16'b0000_0000_0000_0000;
array[9360] <= 16'b0000_0000_0000_0000;
array[9361] <= 16'b0000_0000_0000_0000;
array[9362] <= 16'b0000_0000_0000_0000;
array[9363] <= 16'b0000_0000_0000_0000;
array[9364] <= 16'b0000_0000_0000_0000;
array[9365] <= 16'b0000_0000_0000_0000;
array[9366] <= 16'b0000_0000_0000_0000;
array[9367] <= 16'b0000_0000_0000_0000;
array[9368] <= 16'b0000_0000_0000_0000;
array[9369] <= 16'b0000_0000_0000_0000;
array[9370] <= 16'b0000_0000_0000_0000;
array[9371] <= 16'b0000_0000_0000_0000;
array[9372] <= 16'b0000_0000_0000_0000;
array[9373] <= 16'b0000_0000_0000_0000;
array[9374] <= 16'b0000_0000_0000_0000;
array[9375] <= 16'b0000_0000_0000_0000;
array[9376] <= 16'b0000_0000_0000_0000;
array[9377] <= 16'b0000_0000_0000_0000;
array[9378] <= 16'b0000_0000_0000_0000;
array[9379] <= 16'b0000_0000_0000_0000;
array[9380] <= 16'b0000_0000_0000_0000;
array[9381] <= 16'b0000_0000_0000_0000;
array[9382] <= 16'b0000_0000_0000_0000;
array[9383] <= 16'b0000_0000_0000_0000;
array[9384] <= 16'b0000_0000_0000_0000;
array[9385] <= 16'b0000_0000_0000_0000;
array[9386] <= 16'b0000_0000_0000_0000;
array[9387] <= 16'b0000_0000_0000_0000;
array[9388] <= 16'b0000_0000_0000_0000;
array[9389] <= 16'b0000_0000_0000_0000;
array[9390] <= 16'b0000_0000_0000_0000;
array[9391] <= 16'b0000_0000_0000_0000;
array[9392] <= 16'b0000_0000_0000_0000;
array[9393] <= 16'b0000_0000_0000_0000;
array[9394] <= 16'b0000_0000_0000_0000;
array[9395] <= 16'b0000_0000_0000_0000;
array[9396] <= 16'b0000_0000_0000_0000;
array[9397] <= 16'b0000_0000_0000_0000;
array[9398] <= 16'b0000_0000_0000_0000;
array[9399] <= 16'b0000_0000_0000_0000;
array[9400] <= 16'b0000_0000_0000_0000;
array[9401] <= 16'b0000_0000_0000_0000;
array[9402] <= 16'b0000_0000_0000_0000;
array[9403] <= 16'b0000_0000_0000_0000;
array[9404] <= 16'b0000_0000_0000_0000;
array[9405] <= 16'b0000_0000_0000_0000;
array[9406] <= 16'b0000_0000_0000_0000;
array[9407] <= 16'b0000_0000_0000_0000;
array[9408] <= 16'b0000_0000_0000_0000;
array[9409] <= 16'b0000_0000_0000_0000;
array[9410] <= 16'b0000_0000_0000_0000;
array[9411] <= 16'b0000_0000_0000_0000;
array[9412] <= 16'b0000_0000_0000_0000;
array[9413] <= 16'b0000_0000_0000_0000;
array[9414] <= 16'b0000_0000_0000_0000;
array[9415] <= 16'b0000_0000_0000_0000;
array[9416] <= 16'b0000_0000_0000_0000;
array[9417] <= 16'b0000_0000_0000_0000;
array[9418] <= 16'b0000_0000_0000_0000;
array[9419] <= 16'b0000_0000_0000_0000;
array[9420] <= 16'b0000_0000_0000_0000;
array[9421] <= 16'b0000_0000_0000_0000;
array[9422] <= 16'b0000_0000_0000_0000;
array[9423] <= 16'b0000_0000_0000_0000;
array[9424] <= 16'b0000_0000_0000_0000;
array[9425] <= 16'b0000_0000_0000_0000;
array[9426] <= 16'b0000_0000_0000_0000;
array[9427] <= 16'b0000_0000_0000_0000;
array[9428] <= 16'b0000_0000_0000_0000;
array[9429] <= 16'b0000_0000_0000_0000;
array[9430] <= 16'b0000_0000_0000_0000;
array[9431] <= 16'b0000_0000_0000_0000;
array[9432] <= 16'b0000_0000_0000_0000;
array[9433] <= 16'b0000_0000_0000_0000;
array[9434] <= 16'b0000_0000_0000_0000;
array[9435] <= 16'b0000_0000_0000_0000;
array[9436] <= 16'b0000_0000_0000_0000;
array[9437] <= 16'b0000_0000_0000_0000;
array[9438] <= 16'b0000_0000_0000_0000;
array[9439] <= 16'b0000_0000_0000_0000;
array[9440] <= 16'b0000_0000_0000_0000;
array[9441] <= 16'b0000_0000_0000_0000;
array[9442] <= 16'b0000_0000_0000_0000;
array[9443] <= 16'b0000_0000_0000_0000;
array[9444] <= 16'b0000_0000_0000_0000;
array[9445] <= 16'b0000_0000_0000_0000;
array[9446] <= 16'b0000_0000_0000_0000;
array[9447] <= 16'b0000_0000_0000_0000;
array[9448] <= 16'b0000_0000_0000_0000;
array[9449] <= 16'b0000_0000_0000_0000;
array[9450] <= 16'b0000_0000_0000_0000;
array[9451] <= 16'b0000_0000_0000_0000;
array[9452] <= 16'b0000_0000_0000_0000;
array[9453] <= 16'b0000_0000_0000_0000;
array[9454] <= 16'b0000_0000_0000_0000;
array[9455] <= 16'b0000_0000_0000_0000;
array[9456] <= 16'b0000_0000_0000_0000;
array[9457] <= 16'b0000_0000_0000_0000;
array[9458] <= 16'b0000_0000_0000_0000;
array[9459] <= 16'b0000_0000_0000_0000;
array[9460] <= 16'b0000_0000_0000_0000;
array[9461] <= 16'b0000_0000_0000_0000;
array[9462] <= 16'b0000_0000_0000_0000;
array[9463] <= 16'b0000_0000_0000_0000;
array[9464] <= 16'b0000_0000_0000_0000;
array[9465] <= 16'b0000_0000_0000_0000;
array[9466] <= 16'b0000_0000_0000_0000;
array[9467] <= 16'b0000_0000_0000_0000;
array[9468] <= 16'b0000_0000_0000_0000;
array[9469] <= 16'b0000_0000_0000_0000;
array[9470] <= 16'b0000_0000_0000_0000;
array[9471] <= 16'b0000_0000_0000_0000;
array[9472] <= 16'b0000_0000_0000_0000;
array[9473] <= 16'b0000_0000_0000_0000;
array[9474] <= 16'b0000_0000_0000_0000;
array[9475] <= 16'b0000_0000_0000_0000;
array[9476] <= 16'b0000_0000_0000_0000;
array[9477] <= 16'b0000_0000_0000_0000;
array[9478] <= 16'b0000_0000_0000_0000;
array[9479] <= 16'b0000_0000_0000_0000;
array[9480] <= 16'b0000_0000_0000_0000;
array[9481] <= 16'b0000_0000_0000_0000;
array[9482] <= 16'b0000_0000_0000_0000;
array[9483] <= 16'b0000_0000_0000_0000;
array[9484] <= 16'b0000_0000_0000_0000;
array[9485] <= 16'b0000_0000_0000_0000;
array[9486] <= 16'b0000_0000_0000_0000;
array[9487] <= 16'b0000_0000_0000_0000;
array[9488] <= 16'b0000_0000_0000_0000;
array[9489] <= 16'b0000_0000_0000_0000;
array[9490] <= 16'b0000_0000_0000_0000;
array[9491] <= 16'b0000_0000_0000_0000;
array[9492] <= 16'b0000_0000_0000_0000;
array[9493] <= 16'b0000_0000_0000_0000;
array[9494] <= 16'b0000_0000_0000_0000;
array[9495] <= 16'b0000_0000_0000_0000;
array[9496] <= 16'b0000_0000_0000_0000;
array[9497] <= 16'b0000_0000_0000_0000;
array[9498] <= 16'b0000_0000_0000_0000;
array[9499] <= 16'b0000_0000_0000_0000;
array[9500] <= 16'b0000_0000_0000_0000;
array[9501] <= 16'b0000_0000_0000_0000;
array[9502] <= 16'b0000_0000_0000_0000;
array[9503] <= 16'b0000_0000_0000_0000;
array[9504] <= 16'b0000_0000_0000_0000;
array[9505] <= 16'b0000_0000_0000_0000;
array[9506] <= 16'b0000_0000_0000_0000;
array[9507] <= 16'b0000_0000_0000_0000;
array[9508] <= 16'b0000_0000_0000_0000;
array[9509] <= 16'b0000_0000_0000_0000;
array[9510] <= 16'b0000_0000_0000_0000;
array[9511] <= 16'b0000_0000_0000_0000;
array[9512] <= 16'b0000_0000_0000_0000;
array[9513] <= 16'b0000_0000_0000_0000;
array[9514] <= 16'b0000_0000_0000_0000;
array[9515] <= 16'b0000_0000_0000_0000;
array[9516] <= 16'b0000_0000_0000_0000;
array[9517] <= 16'b0000_0000_0000_0000;
array[9518] <= 16'b0000_0000_0000_0000;
array[9519] <= 16'b0000_0000_0000_0000;
array[9520] <= 16'b0000_0000_0000_0000;
array[9521] <= 16'b0000_0000_0000_0000;
array[9522] <= 16'b0000_0000_0000_0000;
array[9523] <= 16'b0000_0000_0000_0000;
array[9524] <= 16'b0000_0000_0000_0000;
array[9525] <= 16'b0000_0000_0000_0000;
array[9526] <= 16'b0000_0000_0000_0000;
array[9527] <= 16'b0000_0000_0000_0000;
array[9528] <= 16'b0000_0000_0000_0000;
array[9529] <= 16'b0000_0000_0000_0000;
array[9530] <= 16'b0000_0000_0000_0000;
array[9531] <= 16'b0000_0000_0000_0000;
array[9532] <= 16'b0000_0000_0000_0000;
array[9533] <= 16'b0000_0000_0000_0000;
array[9534] <= 16'b0000_0000_0000_0000;
array[9535] <= 16'b0000_0000_0000_0000;
array[9536] <= 16'b0000_0000_0000_0000;
array[9537] <= 16'b0000_0000_0000_0000;
array[9538] <= 16'b0000_0000_0000_0000;
array[9539] <= 16'b0000_0000_0000_0000;
array[9540] <= 16'b0000_0000_0000_0000;
array[9541] <= 16'b0000_0000_0000_0000;
array[9542] <= 16'b0000_0000_0000_0000;
array[9543] <= 16'b0000_0000_0000_0000;
array[9544] <= 16'b0000_0000_0000_0000;
array[9545] <= 16'b0000_0000_0000_0000;
array[9546] <= 16'b0000_0000_0000_0000;
array[9547] <= 16'b0000_0000_0000_0000;
array[9548] <= 16'b0000_0000_0000_0000;
array[9549] <= 16'b0000_0000_0000_0000;
array[9550] <= 16'b0000_0000_0000_0000;
array[9551] <= 16'b0000_0000_0000_0000;
array[9552] <= 16'b0000_0000_0000_0000;
array[9553] <= 16'b0000_0000_0000_0000;
array[9554] <= 16'b0000_0000_0000_0000;
array[9555] <= 16'b0000_0000_0000_0000;
array[9556] <= 16'b0000_0000_0000_0000;
array[9557] <= 16'b0000_0000_0000_0000;
array[9558] <= 16'b0000_0000_0000_0000;
array[9559] <= 16'b0000_0000_0000_0000;
array[9560] <= 16'b0000_0000_0000_0000;
array[9561] <= 16'b0000_0000_0000_0000;
array[9562] <= 16'b0000_0000_0000_0000;
array[9563] <= 16'b0000_0000_0000_0000;
array[9564] <= 16'b0000_0000_0000_0000;
array[9565] <= 16'b0000_0000_0000_0000;
array[9566] <= 16'b0000_0000_0000_0000;
array[9567] <= 16'b0000_0000_0000_0000;
array[9568] <= 16'b0000_0000_0000_0000;
array[9569] <= 16'b0000_0000_0000_0000;
array[9570] <= 16'b0000_0000_0000_0000;
array[9571] <= 16'b0000_0000_0000_0000;
array[9572] <= 16'b0000_0000_0000_0000;
array[9573] <= 16'b0000_0000_0000_0000;
array[9574] <= 16'b0000_0000_0000_0000;
array[9575] <= 16'b0000_0000_0000_0000;
array[9576] <= 16'b0000_0000_0000_0000;
array[9577] <= 16'b0000_0000_0000_0000;
array[9578] <= 16'b0000_0000_0000_0000;
array[9579] <= 16'b0000_0000_0000_0000;
array[9580] <= 16'b0000_0000_0000_0000;
array[9581] <= 16'b0000_0000_0000_0000;
array[9582] <= 16'b0000_0000_0000_0000;
array[9583] <= 16'b0000_0000_0000_0000;
array[9584] <= 16'b0000_0000_0000_0000;
array[9585] <= 16'b0000_0000_0000_0000;
array[9586] <= 16'b0000_0000_0000_0000;
array[9587] <= 16'b0000_0000_0000_0000;
array[9588] <= 16'b0000_0000_0000_0000;
array[9589] <= 16'b0000_0000_0000_0000;
array[9590] <= 16'b0000_0000_0000_0000;
array[9591] <= 16'b0000_0000_0000_0000;
array[9592] <= 16'b0000_0000_0000_0000;
array[9593] <= 16'b0000_0000_0000_0000;
array[9594] <= 16'b0000_0000_0000_0000;
array[9595] <= 16'b0000_0000_0000_0000;
array[9596] <= 16'b0000_0000_0000_0000;
array[9597] <= 16'b0000_0000_0000_0000;
array[9598] <= 16'b0000_0000_0000_0000;
array[9599] <= 16'b0000_0000_0000_0000;
array[9600] <= 16'b0000_0000_0000_0000;
array[9601] <= 16'b0000_0000_0000_0000;
array[9602] <= 16'b0000_0000_0000_0000;
array[9603] <= 16'b0000_0000_0000_0000;
array[9604] <= 16'b0000_0000_0000_0000;
array[9605] <= 16'b0000_0000_0000_0000;
array[9606] <= 16'b0000_0000_0000_0000;
array[9607] <= 16'b0000_0000_0000_0000;
array[9608] <= 16'b0000_0000_0000_0000;
array[9609] <= 16'b0000_0000_0000_0000;
array[9610] <= 16'b0000_0000_0000_0000;
array[9611] <= 16'b0000_0000_0000_0000;
array[9612] <= 16'b0000_0000_0000_0000;
array[9613] <= 16'b0000_0000_0000_0000;
array[9614] <= 16'b0000_0000_0000_0000;
array[9615] <= 16'b0000_0000_0000_0000;
array[9616] <= 16'b0000_0000_0000_0000;
array[9617] <= 16'b0000_0000_0000_0000;
array[9618] <= 16'b0000_0000_0000_0000;
array[9619] <= 16'b0000_0000_0000_0000;
array[9620] <= 16'b0000_0000_0000_0000;
array[9621] <= 16'b0000_0000_0000_0000;
array[9622] <= 16'b0000_0000_0000_0000;
array[9623] <= 16'b0000_0000_0000_0000;
array[9624] <= 16'b0000_0000_0000_0000;
array[9625] <= 16'b0000_0000_0000_0000;
array[9626] <= 16'b0000_0000_0000_0000;
array[9627] <= 16'b0000_0000_0000_0000;
array[9628] <= 16'b0000_0000_0000_0000;
array[9629] <= 16'b0000_0000_0000_0000;
array[9630] <= 16'b0000_0000_0000_0000;
array[9631] <= 16'b0000_0000_0000_0000;
array[9632] <= 16'b0000_0000_0000_0000;
array[9633] <= 16'b0000_0000_0000_0000;
array[9634] <= 16'b0000_0000_0000_0000;
array[9635] <= 16'b0000_0000_0000_0000;
array[9636] <= 16'b0000_0000_0000_0000;
array[9637] <= 16'b0000_0000_0000_0000;
array[9638] <= 16'b0000_0000_0000_0000;
array[9639] <= 16'b0000_0000_0000_0000;
array[9640] <= 16'b0000_0000_0000_0000;
array[9641] <= 16'b0000_0000_0000_0000;
array[9642] <= 16'b0000_0000_0000_0000;
array[9643] <= 16'b0000_0000_0000_0000;
array[9644] <= 16'b0000_0000_0000_0000;
array[9645] <= 16'b0000_0000_0000_0000;
array[9646] <= 16'b0000_0000_0000_0000;
array[9647] <= 16'b0000_0000_0000_0000;
array[9648] <= 16'b0000_0000_0000_0000;
array[9649] <= 16'b0000_0000_0000_0000;
array[9650] <= 16'b0000_0000_0000_0000;
array[9651] <= 16'b0000_0000_0000_0000;
array[9652] <= 16'b0000_0000_0000_0000;
array[9653] <= 16'b0000_0000_0000_0000;
array[9654] <= 16'b0000_0000_0000_0000;
array[9655] <= 16'b0000_0000_0000_0000;
array[9656] <= 16'b0000_0000_0000_0000;
array[9657] <= 16'b0000_0000_0000_0000;
array[9658] <= 16'b0000_0000_0000_0000;
array[9659] <= 16'b0000_0000_0000_0000;
array[9660] <= 16'b0000_0000_0000_0000;
array[9661] <= 16'b0000_0000_0000_0000;
array[9662] <= 16'b0000_0000_0000_0000;
array[9663] <= 16'b0000_0000_0000_0000;
array[9664] <= 16'b0000_0000_0000_0000;
array[9665] <= 16'b0000_0000_0000_0000;
array[9666] <= 16'b0000_0000_0000_0000;
array[9667] <= 16'b0000_0000_0000_0000;
array[9668] <= 16'b0000_0000_0000_0000;
array[9669] <= 16'b0000_0000_0000_0000;
array[9670] <= 16'b0000_0000_0000_0000;
array[9671] <= 16'b0000_0000_0000_0000;
array[9672] <= 16'b0000_0000_0000_0000;
array[9673] <= 16'b0000_0000_0000_0000;
array[9674] <= 16'b0000_0000_0000_0000;
array[9675] <= 16'b0000_0000_0000_0000;
array[9676] <= 16'b0000_0000_0000_0000;
array[9677] <= 16'b0000_0000_0000_0000;
array[9678] <= 16'b0000_0000_0000_0000;
array[9679] <= 16'b0000_0000_0000_0000;
array[9680] <= 16'b0000_0000_0000_0000;
array[9681] <= 16'b0000_0000_0000_0000;
array[9682] <= 16'b0000_0000_0000_0000;
array[9683] <= 16'b0000_0000_0000_0000;
array[9684] <= 16'b0000_0000_0000_0000;
array[9685] <= 16'b0000_0000_0000_0000;
array[9686] <= 16'b0000_0000_0000_0000;
array[9687] <= 16'b0000_0000_0000_0000;
array[9688] <= 16'b0000_0000_0000_0000;
array[9689] <= 16'b0000_0000_0000_0000;
array[9690] <= 16'b0000_0000_0000_0000;
array[9691] <= 16'b0000_0000_0000_0000;
array[9692] <= 16'b0000_0000_0000_0000;
array[9693] <= 16'b0000_0000_0000_0000;
array[9694] <= 16'b0000_0000_0000_0000;
array[9695] <= 16'b0000_0000_0000_0000;
array[9696] <= 16'b0000_0000_0000_0000;
array[9697] <= 16'b0000_0000_0000_0000;
array[9698] <= 16'b0000_0000_0000_0000;
array[9699] <= 16'b0000_0000_0000_0000;
array[9700] <= 16'b0000_0000_0000_0000;
array[9701] <= 16'b0000_0000_0000_0000;
array[9702] <= 16'b0000_0000_0000_0000;
array[9703] <= 16'b0000_0000_0000_0000;
array[9704] <= 16'b0000_0000_0000_0000;
array[9705] <= 16'b0000_0000_0000_0000;
array[9706] <= 16'b0000_0000_0000_0000;
array[9707] <= 16'b0000_0000_0000_0000;
array[9708] <= 16'b0000_0000_0000_0000;
array[9709] <= 16'b0000_0000_0000_0000;
array[9710] <= 16'b0000_0000_0000_0000;
array[9711] <= 16'b0000_0000_0000_0000;
array[9712] <= 16'b0000_0000_0000_0000;
array[9713] <= 16'b0000_0000_0000_0000;
array[9714] <= 16'b0000_0000_0000_0000;
array[9715] <= 16'b0000_0000_0000_0000;
array[9716] <= 16'b0000_0000_0000_0000;
array[9717] <= 16'b0000_0000_0000_0000;
array[9718] <= 16'b0000_0000_0000_0000;
array[9719] <= 16'b0000_0000_0000_0000;
array[9720] <= 16'b0000_0000_0000_0000;
array[9721] <= 16'b0000_0000_0000_0000;
array[9722] <= 16'b0000_0000_0000_0000;
array[9723] <= 16'b0000_0000_0000_0000;
array[9724] <= 16'b0000_0000_0000_0000;
array[9725] <= 16'b0000_0000_0000_0000;
array[9726] <= 16'b0000_0000_0000_0000;
array[9727] <= 16'b0000_0000_0000_0000;
array[9728] <= 16'b0000_0000_0000_0000;
array[9729] <= 16'b0000_0000_0000_0000;
array[9730] <= 16'b0000_0000_0000_0000;
array[9731] <= 16'b0000_0000_0000_0000;
array[9732] <= 16'b0000_0000_0000_0000;
array[9733] <= 16'b0000_0000_0000_0000;
array[9734] <= 16'b0000_0000_0000_0000;
array[9735] <= 16'b0000_0000_0000_0000;
array[9736] <= 16'b0000_0000_0000_0000;
array[9737] <= 16'b0000_0000_0000_0000;
array[9738] <= 16'b0000_0000_0000_0000;
array[9739] <= 16'b0000_0000_0000_0000;
array[9740] <= 16'b0000_0000_0000_0000;
array[9741] <= 16'b0000_0000_0000_0000;
array[9742] <= 16'b0000_0000_0000_0000;
array[9743] <= 16'b0000_0000_0000_0000;
array[9744] <= 16'b0000_0000_0000_0000;
array[9745] <= 16'b0000_0000_0000_0000;
array[9746] <= 16'b0000_0000_0000_0000;
array[9747] <= 16'b0000_0000_0000_0000;
array[9748] <= 16'b0000_0000_0000_0000;
array[9749] <= 16'b0000_0000_0000_0000;
array[9750] <= 16'b0000_0000_0000_0000;
array[9751] <= 16'b0000_0000_0000_0000;
array[9752] <= 16'b0000_0000_0000_0000;
array[9753] <= 16'b0000_0000_0000_0000;
array[9754] <= 16'b0000_0000_0000_0000;
array[9755] <= 16'b0000_0000_0000_0000;
array[9756] <= 16'b0000_0000_0000_0000;
array[9757] <= 16'b0000_0000_0000_0000;
array[9758] <= 16'b0000_0000_0000_0000;
array[9759] <= 16'b0000_0000_0000_0000;
array[9760] <= 16'b0000_0000_0000_0000;
array[9761] <= 16'b0000_0000_0000_0000;
array[9762] <= 16'b0000_0000_0000_0000;
array[9763] <= 16'b0000_0000_0000_0000;
array[9764] <= 16'b0000_0000_0000_0000;
array[9765] <= 16'b0000_0000_0000_0000;
array[9766] <= 16'b0000_0000_0000_0000;
array[9767] <= 16'b0000_0000_0000_0000;
array[9768] <= 16'b0000_0000_0000_0000;
array[9769] <= 16'b0000_0000_0000_0000;
array[9770] <= 16'b0000_0000_0000_0000;
array[9771] <= 16'b0000_0000_0000_0000;
array[9772] <= 16'b0000_0000_0000_0000;
array[9773] <= 16'b0000_0000_0000_0000;
array[9774] <= 16'b0000_0000_0000_0000;
array[9775] <= 16'b0000_0000_0000_0000;
array[9776] <= 16'b0000_0000_0000_0000;
array[9777] <= 16'b0000_0000_0000_0000;
array[9778] <= 16'b0000_0000_0000_0000;
array[9779] <= 16'b0000_0000_0000_0000;
array[9780] <= 16'b0000_0000_0000_0000;
array[9781] <= 16'b0000_0000_0000_0000;
array[9782] <= 16'b0000_0000_0000_0000;
array[9783] <= 16'b0000_0000_0000_0000;
array[9784] <= 16'b0000_0000_0000_0000;
array[9785] <= 16'b0000_0000_0000_0000;
array[9786] <= 16'b0000_0000_0000_0000;
array[9787] <= 16'b0000_0000_0000_0000;
array[9788] <= 16'b0000_0000_0000_0000;
array[9789] <= 16'b0000_0000_0000_0000;
array[9790] <= 16'b0000_0000_0000_0000;
array[9791] <= 16'b0000_0000_0000_0000;
array[9792] <= 16'b0000_0000_0000_0000;
array[9793] <= 16'b0000_0000_0000_0000;
array[9794] <= 16'b0000_0000_0000_0000;
array[9795] <= 16'b0000_0000_0000_0000;
array[9796] <= 16'b0000_0000_0000_0000;
array[9797] <= 16'b0000_0000_0000_0000;
array[9798] <= 16'b0000_0000_0000_0000;
array[9799] <= 16'b0000_0000_0000_0000;
array[9800] <= 16'b0000_0000_0000_0000;
array[9801] <= 16'b0000_0000_0000_0000;
array[9802] <= 16'b0000_0000_0000_0000;
array[9803] <= 16'b0000_0000_0000_0000;
array[9804] <= 16'b0000_0000_0000_0000;
array[9805] <= 16'b0000_0000_0000_0000;
array[9806] <= 16'b0000_0000_0000_0000;
array[9807] <= 16'b0000_0000_0000_0000;
array[9808] <= 16'b0000_0000_0000_0000;
array[9809] <= 16'b0000_0000_0000_0000;
array[9810] <= 16'b0000_0000_0000_0000;
array[9811] <= 16'b0000_0000_0000_0000;
array[9812] <= 16'b0000_0000_0000_0000;
array[9813] <= 16'b0000_0000_0000_0000;
array[9814] <= 16'b0000_0000_0000_0000;
array[9815] <= 16'b0000_0000_0000_0000;
array[9816] <= 16'b0000_0000_0000_0000;
array[9817] <= 16'b0000_0000_0000_0000;
array[9818] <= 16'b0000_0000_0000_0000;
array[9819] <= 16'b0000_0000_0000_0000;
array[9820] <= 16'b0000_0000_0000_0000;
array[9821] <= 16'b0000_0000_0000_0000;
array[9822] <= 16'b0000_0000_0000_0000;
array[9823] <= 16'b0000_0000_0000_0000;
array[9824] <= 16'b0000_0000_0000_0000;
array[9825] <= 16'b0000_0000_0000_0000;
array[9826] <= 16'b0000_0000_0000_0000;
array[9827] <= 16'b0000_0000_0000_0000;
array[9828] <= 16'b0000_0000_0000_0000;
array[9829] <= 16'b0000_0000_0000_0000;
array[9830] <= 16'b0000_0000_0000_0000;
array[9831] <= 16'b0000_0000_0000_0000;
array[9832] <= 16'b0000_0000_0000_0000;
array[9833] <= 16'b0000_0000_0000_0000;
array[9834] <= 16'b0000_0000_0000_0000;
array[9835] <= 16'b0000_0000_0000_0000;
array[9836] <= 16'b0000_0000_0000_0000;
array[9837] <= 16'b0000_0000_0000_0000;
array[9838] <= 16'b0000_0000_0000_0000;
array[9839] <= 16'b0000_0000_0000_0000;
array[9840] <= 16'b0000_0000_0000_0000;
array[9841] <= 16'b0000_0000_0000_0000;
array[9842] <= 16'b0000_0000_0000_0000;
array[9843] <= 16'b0000_0000_0000_0000;
array[9844] <= 16'b0000_0000_0000_0000;
array[9845] <= 16'b0000_0000_0000_0000;
array[9846] <= 16'b0000_0000_0000_0000;
array[9847] <= 16'b0000_0000_0000_0000;
array[9848] <= 16'b0000_0000_0000_0000;
array[9849] <= 16'b0000_0000_0000_0000;
array[9850] <= 16'b0000_0000_0000_0000;
array[9851] <= 16'b0000_0000_0000_0000;
array[9852] <= 16'b0000_0000_0000_0000;
array[9853] <= 16'b0000_0000_0000_0000;
array[9854] <= 16'b0000_0000_0000_0000;
array[9855] <= 16'b0000_0000_0000_0000;
array[9856] <= 16'b0000_0000_0000_0000;
array[9857] <= 16'b0000_0000_0000_0000;
array[9858] <= 16'b0000_0000_0000_0000;
array[9859] <= 16'b0000_0000_0000_0000;
array[9860] <= 16'b0000_0000_0000_0000;
array[9861] <= 16'b0000_0000_0000_0000;
array[9862] <= 16'b0000_0000_0000_0000;
array[9863] <= 16'b0000_0000_0000_0000;
array[9864] <= 16'b0000_0000_0000_0000;
array[9865] <= 16'b0000_0000_0000_0000;
array[9866] <= 16'b0000_0000_0000_0000;
array[9867] <= 16'b0000_0000_0000_0000;
array[9868] <= 16'b0000_0000_0000_0000;
array[9869] <= 16'b0000_0000_0000_0000;
array[9870] <= 16'b0000_0000_0000_0000;
array[9871] <= 16'b0000_0000_0000_0000;
array[9872] <= 16'b0000_0000_0000_0000;
array[9873] <= 16'b0000_0000_0000_0000;
array[9874] <= 16'b0000_0000_0000_0000;
array[9875] <= 16'b0000_0000_0000_0000;
array[9876] <= 16'b0000_0000_0000_0000;
array[9877] <= 16'b0000_0000_0000_0000;
array[9878] <= 16'b0000_0000_0000_0000;
array[9879] <= 16'b0000_0000_0000_0000;
array[9880] <= 16'b0000_0000_0000_0000;
array[9881] <= 16'b0000_0000_0000_0000;
array[9882] <= 16'b0000_0000_0000_0000;
array[9883] <= 16'b0000_0000_0000_0000;
array[9884] <= 16'b0000_0000_0000_0000;
array[9885] <= 16'b0000_0000_0000_0000;
array[9886] <= 16'b0000_0000_0000_0000;
array[9887] <= 16'b0000_0000_0000_0000;
array[9888] <= 16'b0000_0000_0000_0000;
array[9889] <= 16'b0000_0000_0000_0000;
array[9890] <= 16'b0000_0000_0000_0000;
array[9891] <= 16'b0000_0000_0000_0000;
array[9892] <= 16'b0000_0000_0000_0000;
array[9893] <= 16'b0000_0000_0000_0000;
array[9894] <= 16'b0000_0000_0000_0000;
array[9895] <= 16'b0000_0000_0000_0000;
array[9896] <= 16'b0000_0000_0000_0000;
array[9897] <= 16'b0000_0000_0000_0000;
array[9898] <= 16'b0000_0000_0000_0000;
array[9899] <= 16'b0000_0000_0000_0000;
array[9900] <= 16'b0000_0000_0000_0000;
array[9901] <= 16'b0000_0000_0000_0000;
array[9902] <= 16'b0000_0000_0000_0000;
array[9903] <= 16'b0000_0000_0000_0000;
array[9904] <= 16'b0000_0000_0000_0000;
array[9905] <= 16'b0000_0000_0000_0000;
array[9906] <= 16'b0000_0000_0000_0000;
array[9907] <= 16'b0000_0000_0000_0000;
array[9908] <= 16'b0000_0000_0000_0000;
array[9909] <= 16'b0000_0000_0000_0000;
array[9910] <= 16'b0000_0000_0000_0000;
array[9911] <= 16'b0000_0000_0000_0000;
array[9912] <= 16'b0000_0000_0000_0000;
array[9913] <= 16'b0000_0000_0000_0000;
array[9914] <= 16'b0000_0000_0000_0000;
array[9915] <= 16'b0000_0000_0000_0000;
array[9916] <= 16'b0000_0000_0000_0000;
array[9917] <= 16'b0000_0000_0000_0000;
array[9918] <= 16'b0000_0000_0000_0000;
array[9919] <= 16'b0000_0000_0000_0000;
array[9920] <= 16'b0000_0000_0000_0000;
array[9921] <= 16'b0000_0000_0000_0000;
array[9922] <= 16'b0000_0000_0000_0000;
array[9923] <= 16'b0000_0000_0000_0000;
array[9924] <= 16'b0000_0000_0000_0000;
array[9925] <= 16'b0000_0000_0000_0000;
array[9926] <= 16'b0000_0000_0000_0000;
array[9927] <= 16'b0000_0000_0000_0000;
array[9928] <= 16'b0000_0000_0000_0000;
array[9929] <= 16'b0000_0000_0000_0000;
array[9930] <= 16'b0000_0000_0000_0000;
array[9931] <= 16'b0000_0000_0000_0000;
array[9932] <= 16'b0000_0000_0000_0000;
array[9933] <= 16'b0000_0000_0000_0000;
array[9934] <= 16'b0000_0000_0000_0000;
array[9935] <= 16'b0000_0000_0000_0000;
array[9936] <= 16'b0000_0000_0000_0000;
array[9937] <= 16'b0000_0000_0000_0000;
array[9938] <= 16'b0000_0000_0000_0000;
array[9939] <= 16'b0000_0000_0000_0000;
array[9940] <= 16'b0000_0000_0000_0000;
array[9941] <= 16'b0000_0000_0000_0000;
array[9942] <= 16'b0000_0000_0000_0000;
array[9943] <= 16'b0000_0000_0000_0000;
array[9944] <= 16'b0000_0000_0000_0000;
array[9945] <= 16'b0000_0000_0000_0000;
array[9946] <= 16'b0000_0000_0000_0000;
array[9947] <= 16'b0000_0000_0000_0000;
array[9948] <= 16'b0000_0000_0000_0000;
array[9949] <= 16'b0000_0000_0000_0000;
array[9950] <= 16'b0000_0000_0000_0000;
array[9951] <= 16'b0000_0000_0000_0000;
array[9952] <= 16'b0000_0000_0000_0000;
array[9953] <= 16'b0000_0000_0000_0000;
array[9954] <= 16'b0000_0000_0000_0000;
array[9955] <= 16'b0000_0000_0000_0000;
array[9956] <= 16'b0000_0000_0000_0000;
array[9957] <= 16'b0000_0000_0000_0000;
array[9958] <= 16'b0000_0000_0000_0000;
array[9959] <= 16'b0000_0000_0000_0000;
array[9960] <= 16'b0000_0000_0000_0000;
array[9961] <= 16'b0000_0000_0000_0000;
array[9962] <= 16'b0000_0000_0000_0000;
array[9963] <= 16'b0000_0000_0000_0000;
array[9964] <= 16'b0000_0000_0000_0000;
array[9965] <= 16'b0000_0000_0000_0000;
array[9966] <= 16'b0000_0000_0000_0000;
array[9967] <= 16'b0000_0000_0000_0000;
array[9968] <= 16'b0000_0000_0000_0000;
array[9969] <= 16'b0000_0000_0000_0000;
array[9970] <= 16'b0000_0000_0000_0000;
array[9971] <= 16'b0000_0000_0000_0000;
array[9972] <= 16'b0000_0000_0000_0000;
array[9973] <= 16'b0000_0000_0000_0000;
array[9974] <= 16'b0000_0000_0000_0000;
array[9975] <= 16'b0000_0000_0000_0000;
array[9976] <= 16'b0000_0000_0000_0000;
array[9977] <= 16'b0000_0000_0000_0000;
array[9978] <= 16'b0000_0000_0000_0000;
array[9979] <= 16'b0000_0000_0000_0000;
array[9980] <= 16'b0000_0000_0000_0000;
array[9981] <= 16'b0000_0000_0000_0000;
array[9982] <= 16'b0000_0000_0000_0000;
array[9983] <= 16'b0000_0000_0000_0000;
array[9984] <= 16'b0000_0000_0000_0000;
array[9985] <= 16'b0000_0000_0000_0000;
array[9986] <= 16'b0000_0000_0000_0000;
array[9987] <= 16'b0000_0000_0000_0000;
array[9988] <= 16'b0000_0000_0000_0000;
array[9989] <= 16'b0000_0000_0000_0000;
array[9990] <= 16'b0000_0000_0000_0000;
array[9991] <= 16'b0000_0000_0000_0000;
array[9992] <= 16'b0000_0000_0000_0000;
array[9993] <= 16'b0000_0000_0000_0000;
array[9994] <= 16'b0000_0000_0000_0000;
array[9995] <= 16'b0000_0000_0000_0000;
array[9996] <= 16'b0000_0000_0000_0000;
array[9997] <= 16'b0000_0000_0000_0000;
array[9998] <= 16'b0000_0000_0000_0000;
array[9999] <= 16'b0000_0000_0000_0000;
array[10000] <= 16'b0000_0000_0000_0000;
array[10001] <= 16'b0000_0000_0000_0000;
array[10002] <= 16'b0000_0000_0000_0000;
array[10003] <= 16'b0000_0000_0000_0000;
array[10004] <= 16'b0000_0000_0000_0000;
array[10005] <= 16'b0000_0000_0000_0000;
array[10006] <= 16'b0000_0000_0000_0000;
array[10007] <= 16'b0000_0000_0000_0000;
array[10008] <= 16'b0000_0000_0000_0000;
array[10009] <= 16'b0000_0000_0000_0000;
array[10010] <= 16'b0000_0000_0000_0000;
array[10011] <= 16'b0000_0000_0000_0000;
array[10012] <= 16'b0000_0000_0000_0000;
array[10013] <= 16'b0000_0000_0000_0000;
array[10014] <= 16'b0000_0000_0000_0000;
array[10015] <= 16'b0000_0000_0000_0000;
array[10016] <= 16'b0000_0000_0000_0000;
array[10017] <= 16'b0000_0000_0000_0000;
array[10018] <= 16'b0000_0000_0000_0000;
array[10019] <= 16'b0000_0000_0000_0000;
array[10020] <= 16'b0000_0000_0000_0000;
array[10021] <= 16'b0000_0000_0000_0000;
array[10022] <= 16'b0000_0000_0000_0000;
array[10023] <= 16'b0000_0000_0000_0000;
array[10024] <= 16'b0000_0000_0000_0000;
array[10025] <= 16'b0000_0000_0000_0000;
array[10026] <= 16'b0000_0000_0000_0000;
array[10027] <= 16'b0000_0000_0000_0000;
array[10028] <= 16'b0000_0000_0000_0000;
array[10029] <= 16'b0000_0000_0000_0000;
array[10030] <= 16'b0000_0000_0000_0000;
array[10031] <= 16'b0000_0000_0000_0000;
array[10032] <= 16'b0000_0000_0000_0000;
array[10033] <= 16'b0000_0000_0000_0000;
array[10034] <= 16'b0000_0000_0000_0000;
array[10035] <= 16'b0000_0000_0000_0000;
array[10036] <= 16'b0000_0000_0000_0000;
array[10037] <= 16'b0000_0000_0000_0000;
array[10038] <= 16'b0000_0000_0000_0000;
array[10039] <= 16'b0000_0000_0000_0000;
array[10040] <= 16'b0000_0000_0000_0000;
array[10041] <= 16'b0000_0000_0000_0000;
array[10042] <= 16'b0000_0000_0000_0000;
array[10043] <= 16'b0000_0000_0000_0000;
array[10044] <= 16'b0000_0000_0000_0000;
array[10045] <= 16'b0000_0000_0000_0000;
array[10046] <= 16'b0000_0000_0000_0000;
array[10047] <= 16'b0000_0000_0000_0000;
array[10048] <= 16'b0000_0000_0000_0000;
array[10049] <= 16'b0000_0000_0000_0000;
array[10050] <= 16'b0000_0000_0000_0000;
array[10051] <= 16'b0000_0000_0000_0000;
array[10052] <= 16'b0000_0000_0000_0000;
array[10053] <= 16'b0000_0000_0000_0000;
array[10054] <= 16'b0000_0000_0000_0000;
array[10055] <= 16'b0000_0000_0000_0000;
array[10056] <= 16'b0000_0000_0000_0000;
array[10057] <= 16'b0000_0000_0000_0000;
array[10058] <= 16'b0000_0000_0000_0000;
array[10059] <= 16'b0000_0000_0000_0000;
array[10060] <= 16'b0000_0000_0000_0000;
array[10061] <= 16'b0000_0000_0000_0000;
array[10062] <= 16'b0000_0000_0000_0000;
array[10063] <= 16'b0000_0000_0000_0000;
array[10064] <= 16'b0000_0000_0000_0000;
array[10065] <= 16'b0000_0000_0000_0000;
array[10066] <= 16'b0000_0000_0000_0000;
array[10067] <= 16'b0000_0000_0000_0000;
array[10068] <= 16'b0000_0000_0000_0000;
array[10069] <= 16'b0000_0000_0000_0000;
array[10070] <= 16'b0000_0000_0000_0000;
array[10071] <= 16'b0000_0000_0000_0000;
array[10072] <= 16'b0000_0000_0000_0000;
array[10073] <= 16'b0000_0000_0000_0000;
array[10074] <= 16'b0000_0000_0000_0000;
array[10075] <= 16'b0000_0000_0000_0000;
array[10076] <= 16'b0000_0000_0000_0000;
array[10077] <= 16'b0000_0000_0000_0000;
array[10078] <= 16'b0000_0000_0000_0000;
array[10079] <= 16'b0000_0000_0000_0000;
array[10080] <= 16'b0000_0000_0000_0000;
array[10081] <= 16'b0000_0000_0000_0000;
array[10082] <= 16'b0000_0000_0000_0000;
array[10083] <= 16'b0000_0000_0000_0000;
array[10084] <= 16'b0000_0000_0000_0000;
array[10085] <= 16'b0000_0000_0000_0000;
array[10086] <= 16'b0000_0000_0000_0000;
array[10087] <= 16'b0000_0000_0000_0000;
array[10088] <= 16'b0000_0000_0000_0000;
array[10089] <= 16'b0000_0000_0000_0000;
array[10090] <= 16'b0000_0000_0000_0000;
array[10091] <= 16'b0000_0000_0000_0000;
array[10092] <= 16'b0000_0000_0000_0000;
array[10093] <= 16'b0000_0000_0000_0000;
array[10094] <= 16'b0000_0000_0000_0000;
array[10095] <= 16'b0000_0000_0000_0000;
array[10096] <= 16'b0000_0000_0000_0000;
array[10097] <= 16'b0000_0000_0000_0000;
array[10098] <= 16'b0000_0000_0000_0000;
array[10099] <= 16'b0000_0000_0000_0000;
array[10100] <= 16'b0000_0000_0000_0000;
array[10101] <= 16'b0000_0000_0000_0000;
array[10102] <= 16'b0000_0000_0000_0000;
array[10103] <= 16'b0000_0000_0000_0000;
array[10104] <= 16'b0000_0000_0000_0000;
array[10105] <= 16'b0000_0000_0000_0000;
array[10106] <= 16'b0000_0000_0000_0000;
array[10107] <= 16'b0000_0000_0000_0000;
array[10108] <= 16'b0000_0000_0000_0000;
array[10109] <= 16'b0000_0000_0000_0000;
array[10110] <= 16'b0000_0000_0000_0000;
array[10111] <= 16'b0000_0000_0000_0000;
array[10112] <= 16'b0000_0000_0000_0000;
array[10113] <= 16'b0000_0000_0000_0000;
array[10114] <= 16'b0000_0000_0000_0000;
array[10115] <= 16'b0000_0000_0000_0000;
array[10116] <= 16'b0000_0000_0000_0000;
array[10117] <= 16'b0000_0000_0000_0000;
array[10118] <= 16'b0000_0000_0000_0000;
array[10119] <= 16'b0000_0000_0000_0000;
array[10120] <= 16'b0000_0000_0000_0000;
array[10121] <= 16'b0000_0000_0000_0000;
array[10122] <= 16'b0000_0000_0000_0000;
array[10123] <= 16'b0000_0000_0000_0000;
array[10124] <= 16'b0000_0000_0000_0000;
array[10125] <= 16'b0000_0000_0000_0000;
array[10126] <= 16'b0000_0000_0000_0000;
array[10127] <= 16'b0000_0000_0000_0000;
array[10128] <= 16'b0000_0000_0000_0000;
array[10129] <= 16'b0000_0000_0000_0000;
array[10130] <= 16'b0000_0000_0000_0000;
array[10131] <= 16'b0000_0000_0000_0000;
array[10132] <= 16'b0000_0000_0000_0000;
array[10133] <= 16'b0000_0000_0000_0000;
array[10134] <= 16'b0000_0000_0000_0000;
array[10135] <= 16'b0000_0000_0000_0000;
array[10136] <= 16'b0000_0000_0000_0000;
array[10137] <= 16'b0000_0000_0000_0000;
array[10138] <= 16'b0000_0000_0000_0000;
array[10139] <= 16'b0000_0000_0000_0000;
array[10140] <= 16'b0000_0000_0000_0000;
array[10141] <= 16'b0000_0000_0000_0000;
array[10142] <= 16'b0000_0000_0000_0000;
array[10143] <= 16'b0000_0000_0000_0000;
array[10144] <= 16'b0000_0000_0000_0000;
array[10145] <= 16'b0000_0000_0000_0000;
array[10146] <= 16'b0000_0000_0000_0000;
array[10147] <= 16'b0000_0000_0000_0000;
array[10148] <= 16'b0000_0000_0000_0000;
array[10149] <= 16'b0000_0000_0000_0000;
array[10150] <= 16'b0000_0000_0000_0000;
array[10151] <= 16'b0000_0000_0000_0000;
array[10152] <= 16'b0000_0000_0000_0000;
array[10153] <= 16'b0000_0000_0000_0000;
array[10154] <= 16'b0000_0000_0000_0000;
array[10155] <= 16'b0000_0000_0000_0000;
array[10156] <= 16'b0000_0000_0000_0000;
array[10157] <= 16'b0000_0000_0000_0000;
array[10158] <= 16'b0000_0000_0000_0000;
array[10159] <= 16'b0000_0000_0000_0000;
array[10160] <= 16'b0000_0000_0000_0000;
array[10161] <= 16'b0000_0000_0000_0000;
array[10162] <= 16'b0000_0000_0000_0000;
array[10163] <= 16'b0000_0000_0000_0000;
array[10164] <= 16'b0000_0000_0000_0000;
array[10165] <= 16'b0000_0000_0000_0000;
array[10166] <= 16'b0000_0000_0000_0000;
array[10167] <= 16'b0000_0000_0000_0000;
array[10168] <= 16'b0000_0000_0000_0000;
array[10169] <= 16'b0000_0000_0000_0000;
array[10170] <= 16'b0000_0000_0000_0000;
array[10171] <= 16'b0000_0000_0000_0000;
array[10172] <= 16'b0000_0000_0000_0000;
array[10173] <= 16'b0000_0000_0000_0000;
array[10174] <= 16'b0000_0000_0000_0000;
array[10175] <= 16'b0000_0000_0000_0000;
array[10176] <= 16'b0000_0000_0000_0000;
array[10177] <= 16'b0000_0000_0000_0000;
array[10178] <= 16'b0000_0000_0000_0000;
array[10179] <= 16'b0000_0000_0000_0000;
array[10180] <= 16'b0000_0000_0000_0000;
array[10181] <= 16'b0000_0000_0000_0000;
array[10182] <= 16'b0000_0000_0000_0000;
array[10183] <= 16'b0000_0000_0000_0000;
array[10184] <= 16'b0000_0000_0000_0000;
array[10185] <= 16'b0000_0000_0000_0000;
array[10186] <= 16'b0000_0000_0000_0000;
array[10187] <= 16'b0000_0000_0000_0000;
array[10188] <= 16'b0000_0000_0000_0000;
array[10189] <= 16'b0000_0000_0000_0000;
array[10190] <= 16'b0000_0000_0000_0000;
array[10191] <= 16'b0000_0000_0000_0000;
array[10192] <= 16'b0000_0000_0000_0000;
array[10193] <= 16'b0000_0000_0000_0000;
array[10194] <= 16'b0000_0000_0000_0000;
array[10195] <= 16'b0000_0000_0000_0000;
array[10196] <= 16'b0000_0000_0000_0000;
array[10197] <= 16'b0000_0000_0000_0000;
array[10198] <= 16'b0000_0000_0000_0000;
array[10199] <= 16'b0000_0000_0000_0000;
array[10200] <= 16'b0000_0000_0000_0000;
array[10201] <= 16'b0000_0000_0000_0000;
array[10202] <= 16'b0000_0000_0000_0000;
array[10203] <= 16'b0000_0000_0000_0000;
array[10204] <= 16'b0000_0000_0000_0000;
array[10205] <= 16'b0000_0000_0000_0000;
array[10206] <= 16'b0000_0000_0000_0000;
array[10207] <= 16'b0000_0000_0000_0000;
array[10208] <= 16'b0000_0000_0000_0000;
array[10209] <= 16'b0000_0000_0000_0000;
array[10210] <= 16'b0000_0000_0000_0000;
array[10211] <= 16'b0000_0000_0000_0000;
array[10212] <= 16'b0000_0000_0000_0000;
array[10213] <= 16'b0000_0000_0000_0000;
array[10214] <= 16'b0000_0000_0000_0000;
array[10215] <= 16'b0000_0000_0000_0000;
array[10216] <= 16'b0000_0000_0000_0000;
array[10217] <= 16'b0000_0000_0000_0000;
array[10218] <= 16'b0000_0000_0000_0000;
array[10219] <= 16'b0000_0000_0000_0000;
array[10220] <= 16'b0000_0000_0000_0000;
array[10221] <= 16'b0000_0000_0000_0000;
array[10222] <= 16'b0000_0000_0000_0000;
array[10223] <= 16'b0000_0000_0000_0000;
array[10224] <= 16'b0000_0000_0000_0000;
array[10225] <= 16'b0000_0000_0000_0000;
array[10226] <= 16'b0000_0000_0000_0000;
array[10227] <= 16'b0000_0000_0000_0000;
array[10228] <= 16'b0000_0000_0000_0000;
array[10229] <= 16'b0000_0000_0000_0000;
array[10230] <= 16'b0000_0000_0000_0000;
array[10231] <= 16'b0000_0000_0000_0000;
array[10232] <= 16'b0000_0000_0000_0000;
array[10233] <= 16'b0000_0000_0000_0000;
array[10234] <= 16'b0000_0000_0000_0000;
array[10235] <= 16'b0000_0000_0000_0000;
array[10236] <= 16'b0000_0000_0000_0000;
array[10237] <= 16'b0000_0000_0000_0000;
array[10238] <= 16'b0000_0000_0000_0000;
array[10239] <= 16'b0000_0000_0000_0000;
array[10240] <= 16'b0000_0000_0000_0000;
array[10241] <= 16'b0000_0000_0000_0000;
array[10242] <= 16'b0000_0000_0000_0000;
array[10243] <= 16'b0000_0000_0000_0000;
array[10244] <= 16'b0000_0000_0000_0000;
array[10245] <= 16'b0000_0000_0000_0000;
array[10246] <= 16'b0000_0000_0000_0000;
array[10247] <= 16'b0000_0000_0000_0000;
array[10248] <= 16'b0000_0000_0000_0000;
array[10249] <= 16'b0000_0000_0000_0000;
array[10250] <= 16'b0000_0000_0000_0000;
array[10251] <= 16'b0000_0000_0000_0000;
array[10252] <= 16'b0000_0000_0000_0000;
array[10253] <= 16'b0000_0000_0000_0000;
array[10254] <= 16'b0000_0000_0000_0000;
array[10255] <= 16'b0000_0000_0000_0000;
array[10256] <= 16'b0000_0000_0000_0000;
array[10257] <= 16'b0000_0000_0000_0000;
array[10258] <= 16'b0000_0000_0000_0000;
array[10259] <= 16'b0000_0000_0000_0000;
array[10260] <= 16'b0000_0000_0000_0000;
array[10261] <= 16'b0000_0000_0000_0000;
array[10262] <= 16'b0000_0000_0000_0000;
array[10263] <= 16'b0000_0000_0000_0000;
array[10264] <= 16'b0000_0000_0000_0000;
array[10265] <= 16'b0000_0000_0000_0000;
array[10266] <= 16'b0000_0000_0000_0000;
array[10267] <= 16'b0000_0000_0000_0000;
array[10268] <= 16'b0000_0000_0000_0000;
array[10269] <= 16'b0000_0000_0000_0000;
array[10270] <= 16'b0000_0000_0000_0000;
array[10271] <= 16'b0000_0000_0000_0000;
array[10272] <= 16'b0000_0000_0000_0000;
array[10273] <= 16'b0000_0000_0000_0000;
array[10274] <= 16'b0000_0000_0000_0000;
array[10275] <= 16'b0000_0000_0000_0000;
array[10276] <= 16'b0000_0000_0000_0000;
array[10277] <= 16'b0000_0000_0000_0000;
array[10278] <= 16'b0000_0000_0000_0000;
array[10279] <= 16'b0000_0000_0000_0000;
array[10280] <= 16'b0000_0000_0000_0000;
array[10281] <= 16'b0000_0000_0000_0000;
array[10282] <= 16'b0000_0000_0000_0000;
array[10283] <= 16'b0000_0000_0000_0000;
array[10284] <= 16'b0000_0000_0000_0000;
array[10285] <= 16'b0000_0000_0000_0000;
array[10286] <= 16'b0000_0000_0000_0000;
array[10287] <= 16'b0000_0000_0000_0000;
array[10288] <= 16'b0000_0000_0000_0000;
array[10289] <= 16'b0000_0000_0000_0000;
array[10290] <= 16'b0000_0000_0000_0000;
array[10291] <= 16'b0000_0000_0000_0000;
array[10292] <= 16'b0000_0000_0000_0000;
array[10293] <= 16'b0000_0000_0000_0000;
array[10294] <= 16'b0000_0000_0000_0000;
array[10295] <= 16'b0000_0000_0000_0000;
array[10296] <= 16'b0000_0000_0000_0000;
array[10297] <= 16'b0000_0000_0000_0000;
array[10298] <= 16'b0000_0000_0000_0000;
array[10299] <= 16'b0000_0000_0000_0000;
array[10300] <= 16'b0000_0000_0000_0000;
array[10301] <= 16'b0000_0000_0000_0000;
array[10302] <= 16'b0000_0000_0000_0000;
array[10303] <= 16'b0000_0000_0000_0000;
array[10304] <= 16'b0000_0000_0000_0000;
array[10305] <= 16'b0000_0000_0000_0000;
array[10306] <= 16'b0000_0000_0000_0000;
array[10307] <= 16'b0000_0000_0000_0000;
array[10308] <= 16'b0000_0000_0000_0000;
array[10309] <= 16'b0000_0000_0000_0000;
array[10310] <= 16'b0000_0000_0000_0000;
array[10311] <= 16'b0000_0000_0000_0000;
array[10312] <= 16'b0000_0000_0000_0000;
array[10313] <= 16'b0000_0000_0000_0000;
array[10314] <= 16'b0000_0000_0000_0000;
array[10315] <= 16'b0000_0000_0000_0000;
array[10316] <= 16'b0000_0000_0000_0000;
array[10317] <= 16'b0000_0000_0000_0000;
array[10318] <= 16'b0000_0000_0000_0000;
array[10319] <= 16'b0000_0000_0000_0000;
array[10320] <= 16'b0000_0000_0000_0000;
array[10321] <= 16'b0000_0000_0000_0000;
array[10322] <= 16'b0000_0000_0000_0000;
array[10323] <= 16'b0000_0000_0000_0000;
array[10324] <= 16'b0000_0000_0000_0000;
array[10325] <= 16'b0000_0000_0000_0000;
array[10326] <= 16'b0000_0000_0000_0000;
array[10327] <= 16'b0000_0000_0000_0000;
array[10328] <= 16'b0000_0000_0000_0000;
array[10329] <= 16'b0000_0000_0000_0000;
array[10330] <= 16'b0000_0000_0000_0000;
array[10331] <= 16'b0000_0000_0000_0000;
array[10332] <= 16'b0000_0000_0000_0000;
array[10333] <= 16'b0000_0000_0000_0000;
array[10334] <= 16'b0000_0000_0000_0000;
array[10335] <= 16'b0000_0000_0000_0000;
array[10336] <= 16'b0000_0000_0000_0000;
array[10337] <= 16'b0000_0000_0000_0000;
array[10338] <= 16'b0000_0000_0000_0000;
array[10339] <= 16'b0000_0000_0000_0000;
array[10340] <= 16'b0000_0000_0000_0000;
array[10341] <= 16'b0000_0000_0000_0000;
array[10342] <= 16'b0000_0000_0000_0000;
array[10343] <= 16'b0000_0000_0000_0000;
array[10344] <= 16'b0000_0000_0000_0000;
array[10345] <= 16'b0000_0000_0000_0000;
array[10346] <= 16'b0000_0000_0000_0000;
array[10347] <= 16'b0000_0000_0000_0000;
array[10348] <= 16'b0000_0000_0000_0000;
array[10349] <= 16'b0000_0000_0000_0000;
array[10350] <= 16'b0000_0000_0000_0000;
array[10351] <= 16'b0000_0000_0000_0000;
array[10352] <= 16'b0000_0000_0000_0000;
array[10353] <= 16'b0000_0000_0000_0000;
array[10354] <= 16'b0000_0000_0000_0000;
array[10355] <= 16'b0000_0000_0000_0000;
array[10356] <= 16'b0000_0000_0000_0000;
array[10357] <= 16'b0000_0000_0000_0000;
array[10358] <= 16'b0000_0000_0000_0000;
array[10359] <= 16'b0000_0000_0000_0000;
array[10360] <= 16'b0000_0000_0000_0000;
array[10361] <= 16'b0000_0000_0000_0000;
array[10362] <= 16'b0000_0000_0000_0000;
array[10363] <= 16'b0000_0000_0000_0000;
array[10364] <= 16'b0000_0000_0000_0000;
array[10365] <= 16'b0000_0000_0000_0000;
array[10366] <= 16'b0000_0000_0000_0000;
array[10367] <= 16'b0000_0000_0000_0000;
array[10368] <= 16'b0000_0000_0000_0000;
array[10369] <= 16'b0000_0000_0000_0000;
array[10370] <= 16'b0000_0000_0000_0000;
array[10371] <= 16'b0000_0000_0000_0000;
array[10372] <= 16'b0000_0000_0000_0000;
array[10373] <= 16'b0000_0000_0000_0000;
array[10374] <= 16'b0000_0000_0000_0000;
array[10375] <= 16'b0000_0000_0000_0000;
array[10376] <= 16'b0000_0000_0000_0000;
array[10377] <= 16'b0000_0000_0000_0000;
array[10378] <= 16'b0000_0000_0000_0000;
array[10379] <= 16'b0000_0000_0000_0000;
array[10380] <= 16'b0000_0000_0000_0000;
array[10381] <= 16'b0000_0000_0000_0000;
array[10382] <= 16'b0000_0000_0000_0000;
array[10383] <= 16'b0000_0000_0000_0000;
array[10384] <= 16'b0000_0000_0000_0000;
array[10385] <= 16'b0000_0000_0000_0000;
array[10386] <= 16'b0000_0000_0000_0000;
array[10387] <= 16'b0000_0000_0000_0000;
array[10388] <= 16'b0000_0000_0000_0000;
array[10389] <= 16'b0000_0000_0000_0000;
array[10390] <= 16'b0000_0000_0000_0000;
array[10391] <= 16'b0000_0000_0000_0000;
array[10392] <= 16'b0000_0000_0000_0000;
array[10393] <= 16'b0000_0000_0000_0000;
array[10394] <= 16'b0000_0000_0000_0000;
array[10395] <= 16'b0000_0000_0000_0000;
array[10396] <= 16'b0000_0000_0000_0000;
array[10397] <= 16'b0000_0000_0000_0000;
array[10398] <= 16'b0000_0000_0000_0000;
array[10399] <= 16'b0000_0000_0000_0000;
array[10400] <= 16'b0000_0000_0000_0000;
array[10401] <= 16'b0000_0000_0000_0000;
array[10402] <= 16'b0000_0000_0000_0000;
array[10403] <= 16'b0000_0000_0000_0000;
array[10404] <= 16'b0000_0000_0000_0000;
array[10405] <= 16'b0000_0000_0000_0000;
array[10406] <= 16'b0000_0000_0000_0000;
array[10407] <= 16'b0000_0000_0000_0000;
array[10408] <= 16'b0000_0000_0000_0000;
array[10409] <= 16'b0000_0000_0000_0000;
array[10410] <= 16'b0000_0000_0000_0000;
array[10411] <= 16'b0000_0000_0000_0000;
array[10412] <= 16'b0000_0000_0000_0000;
array[10413] <= 16'b0000_0000_0000_0000;
array[10414] <= 16'b0000_0000_0000_0000;
array[10415] <= 16'b0000_0000_0000_0000;
array[10416] <= 16'b0000_0000_0000_0000;
array[10417] <= 16'b0000_0000_0000_0000;
array[10418] <= 16'b0000_0000_0000_0000;
array[10419] <= 16'b0000_0000_0000_0000;
array[10420] <= 16'b0000_0000_0000_0000;
array[10421] <= 16'b0000_0000_0000_0000;
array[10422] <= 16'b0000_0000_0000_0000;
array[10423] <= 16'b0000_0000_0000_0000;
array[10424] <= 16'b0000_0000_0000_0000;
array[10425] <= 16'b0000_0000_0000_0000;
array[10426] <= 16'b0000_0000_0000_0000;
array[10427] <= 16'b0000_0000_0000_0000;
array[10428] <= 16'b0000_0000_0000_0000;
array[10429] <= 16'b0000_0000_0000_0000;
array[10430] <= 16'b0000_0000_0000_0000;
array[10431] <= 16'b0000_0000_0000_0000;
array[10432] <= 16'b0000_0000_0000_0000;
array[10433] <= 16'b0000_0000_0000_0000;
array[10434] <= 16'b0000_0000_0000_0000;
array[10435] <= 16'b0000_0000_0000_0000;
array[10436] <= 16'b0000_0000_0000_0000;
array[10437] <= 16'b0000_0000_0000_0000;
array[10438] <= 16'b0000_0000_0000_0000;
array[10439] <= 16'b0000_0000_0000_0000;
array[10440] <= 16'b0000_0000_0000_0000;
array[10441] <= 16'b0000_0000_0000_0000;
array[10442] <= 16'b0000_0000_0000_0000;
array[10443] <= 16'b0000_0000_0000_0000;
array[10444] <= 16'b0000_0000_0000_0000;
array[10445] <= 16'b0000_0000_0000_0000;
array[10446] <= 16'b0000_0000_0000_0000;
array[10447] <= 16'b0000_0000_0000_0000;
array[10448] <= 16'b0000_0000_0000_0000;
array[10449] <= 16'b0000_0000_0000_0000;
array[10450] <= 16'b0000_0000_0000_0000;
array[10451] <= 16'b0000_0000_0000_0000;
array[10452] <= 16'b0000_0000_0000_0000;
array[10453] <= 16'b0000_0000_0000_0000;
array[10454] <= 16'b0000_0000_0000_0000;
array[10455] <= 16'b0000_0000_0000_0000;
array[10456] <= 16'b0000_0000_0000_0000;
array[10457] <= 16'b0000_0000_0000_0000;
array[10458] <= 16'b0000_0000_0000_0000;
array[10459] <= 16'b0000_0000_0000_0000;
array[10460] <= 16'b0000_0000_0000_0000;
array[10461] <= 16'b0000_0000_0000_0000;
array[10462] <= 16'b0000_0000_0000_0000;
array[10463] <= 16'b0000_0000_0000_0000;
array[10464] <= 16'b0000_0000_0000_0000;
array[10465] <= 16'b0000_0000_0000_0000;
array[10466] <= 16'b0000_0000_0000_0000;
array[10467] <= 16'b0000_0000_0000_0000;
array[10468] <= 16'b0000_0000_0000_0000;
array[10469] <= 16'b0000_0000_0000_0000;
array[10470] <= 16'b0000_0000_0000_0000;
array[10471] <= 16'b0000_0000_0000_0000;
array[10472] <= 16'b0000_0000_0000_0000;
array[10473] <= 16'b0000_0000_0000_0000;
array[10474] <= 16'b0000_0000_0000_0000;
array[10475] <= 16'b0000_0000_0000_0000;
array[10476] <= 16'b0000_0000_0000_0000;
array[10477] <= 16'b0000_0000_0000_0000;
array[10478] <= 16'b0000_0000_0000_0000;
array[10479] <= 16'b0000_0000_0000_0000;
array[10480] <= 16'b0000_0000_0000_0000;
array[10481] <= 16'b0000_0000_0000_0000;
array[10482] <= 16'b0000_0000_0000_0000;
array[10483] <= 16'b0000_0000_0000_0000;
array[10484] <= 16'b0000_0000_0000_0000;
array[10485] <= 16'b0000_0000_0000_0000;
array[10486] <= 16'b0000_0000_0000_0000;
array[10487] <= 16'b0000_0000_0000_0000;
array[10488] <= 16'b0000_0000_0000_0000;
array[10489] <= 16'b0000_0000_0000_0000;
array[10490] <= 16'b0000_0000_0000_0000;
array[10491] <= 16'b0000_0000_0000_0000;
array[10492] <= 16'b0000_0000_0000_0000;
array[10493] <= 16'b0000_0000_0000_0000;
array[10494] <= 16'b0000_0000_0000_0000;
array[10495] <= 16'b0000_0000_0000_0000;
array[10496] <= 16'b0000_0000_0000_0000;
array[10497] <= 16'b0000_0000_0000_0000;
array[10498] <= 16'b0000_0000_0000_0000;
array[10499] <= 16'b0000_0000_0000_0000;
array[10500] <= 16'b0000_0000_0000_0000;
array[10501] <= 16'b0000_0000_0000_0000;
array[10502] <= 16'b0000_0000_0000_0000;
array[10503] <= 16'b0000_0000_0000_0000;
array[10504] <= 16'b0000_0000_0000_0000;
array[10505] <= 16'b0000_0000_0000_0000;
array[10506] <= 16'b0000_0000_0000_0000;
array[10507] <= 16'b0000_0000_0000_0000;
array[10508] <= 16'b0000_0000_0000_0000;
array[10509] <= 16'b0000_0000_0000_0000;
array[10510] <= 16'b0000_0000_0000_0000;
array[10511] <= 16'b0000_0000_0000_0000;
array[10512] <= 16'b0000_0000_0000_0000;
array[10513] <= 16'b0000_0000_0000_0000;
array[10514] <= 16'b0000_0000_0000_0000;
array[10515] <= 16'b0000_0000_0000_0000;
array[10516] <= 16'b0000_0000_0000_0000;
array[10517] <= 16'b0000_0000_0000_0000;
array[10518] <= 16'b0000_0000_0000_0000;
array[10519] <= 16'b0000_0000_0000_0000;
array[10520] <= 16'b0000_0000_0000_0000;
array[10521] <= 16'b0000_0000_0000_0000;
array[10522] <= 16'b0000_0000_0000_0000;
array[10523] <= 16'b0000_0000_0000_0000;
array[10524] <= 16'b0000_0000_0000_0000;
array[10525] <= 16'b0000_0000_0000_0000;
array[10526] <= 16'b0000_0000_0000_0000;
array[10527] <= 16'b0000_0000_0000_0000;
array[10528] <= 16'b0000_0000_0000_0000;
array[10529] <= 16'b0000_0000_0000_0000;
array[10530] <= 16'b0000_0000_0000_0000;
array[10531] <= 16'b0000_0000_0000_0000;
array[10532] <= 16'b0000_0000_0000_0000;
array[10533] <= 16'b0000_0000_0000_0000;
array[10534] <= 16'b0000_0000_0000_0000;
array[10535] <= 16'b0000_0000_0000_0000;
array[10536] <= 16'b0000_0000_0000_0000;
array[10537] <= 16'b0000_0000_0000_0000;
array[10538] <= 16'b0000_0000_0000_0000;
array[10539] <= 16'b0000_0000_0000_0000;
array[10540] <= 16'b0000_0000_0000_0000;
array[10541] <= 16'b0000_0000_0000_0000;
array[10542] <= 16'b0000_0000_0000_0000;
array[10543] <= 16'b0000_0000_0000_0000;
array[10544] <= 16'b0000_0000_0000_0000;
array[10545] <= 16'b0000_0000_0000_0000;
array[10546] <= 16'b0000_0000_0000_0000;
array[10547] <= 16'b0000_0000_0000_0000;
array[10548] <= 16'b0000_0000_0000_0000;
array[10549] <= 16'b0000_0000_0000_0000;
array[10550] <= 16'b0000_0000_0000_0000;
array[10551] <= 16'b0000_0000_0000_0000;
array[10552] <= 16'b0000_0000_0000_0000;
array[10553] <= 16'b0000_0000_0000_0000;
array[10554] <= 16'b0000_0000_0000_0000;
array[10555] <= 16'b0000_0000_0000_0000;
array[10556] <= 16'b0000_0000_0000_0000;
array[10557] <= 16'b0000_0000_0000_0000;
array[10558] <= 16'b0000_0000_0000_0000;
array[10559] <= 16'b0000_0000_0000_0000;
array[10560] <= 16'b0000_0000_0000_0000;
array[10561] <= 16'b0000_0000_0000_0000;
array[10562] <= 16'b0000_0000_0000_0000;
array[10563] <= 16'b0000_0000_0000_0000;
array[10564] <= 16'b0000_0000_0000_0000;
array[10565] <= 16'b0000_0000_0000_0000;
array[10566] <= 16'b0000_0000_0000_0000;
array[10567] <= 16'b0000_0000_0000_0000;
array[10568] <= 16'b0000_0000_0000_0000;
array[10569] <= 16'b0000_0000_0000_0000;
array[10570] <= 16'b0000_0000_0000_0000;
array[10571] <= 16'b0000_0000_0000_0000;
array[10572] <= 16'b0000_0000_0000_0000;
array[10573] <= 16'b0000_0000_0000_0000;
array[10574] <= 16'b0000_0000_0000_0000;
array[10575] <= 16'b0000_0000_0000_0000;
array[10576] <= 16'b0000_0000_0000_0000;
array[10577] <= 16'b0000_0000_0000_0000;
array[10578] <= 16'b0000_0000_0000_0000;
array[10579] <= 16'b0000_0000_0000_0000;
array[10580] <= 16'b0000_0000_0000_0000;
array[10581] <= 16'b0000_0000_0000_0000;
array[10582] <= 16'b0000_0000_0000_0000;
array[10583] <= 16'b0000_0000_0000_0000;
array[10584] <= 16'b0000_0000_0000_0000;
array[10585] <= 16'b0000_0000_0000_0000;
array[10586] <= 16'b0000_0000_0000_0000;
array[10587] <= 16'b0000_0000_0000_0000;
array[10588] <= 16'b0000_0000_0000_0000;
array[10589] <= 16'b0000_0000_0000_0000;
array[10590] <= 16'b0000_0000_0000_0000;
array[10591] <= 16'b0000_0000_0000_0000;
array[10592] <= 16'b0000_0000_0000_0000;
array[10593] <= 16'b0000_0000_0000_0000;
array[10594] <= 16'b0000_0000_0000_0000;
array[10595] <= 16'b0000_0000_0000_0000;
array[10596] <= 16'b0000_0000_0000_0000;
array[10597] <= 16'b0000_0000_0000_0000;
array[10598] <= 16'b0000_0000_0000_0000;
array[10599] <= 16'b0000_0000_0000_0000;
array[10600] <= 16'b0000_0000_0000_0000;
array[10601] <= 16'b0000_0000_0000_0000;
array[10602] <= 16'b0000_0000_0000_0000;
array[10603] <= 16'b0000_0000_0000_0000;
array[10604] <= 16'b0000_0000_0000_0000;
array[10605] <= 16'b0000_0000_0000_0000;
array[10606] <= 16'b0000_0000_0000_0000;
array[10607] <= 16'b0000_0000_0000_0000;
array[10608] <= 16'b0000_0000_0000_0000;
array[10609] <= 16'b0000_0000_0000_0000;
array[10610] <= 16'b0000_0000_0000_0000;
array[10611] <= 16'b0000_0000_0000_0000;
array[10612] <= 16'b0000_0000_0000_0000;
array[10613] <= 16'b0000_0000_0000_0000;
array[10614] <= 16'b0000_0000_0000_0000;
array[10615] <= 16'b0000_0000_0000_0000;
array[10616] <= 16'b0000_0000_0000_0000;
array[10617] <= 16'b0000_0000_0000_0000;
array[10618] <= 16'b0000_0000_0000_0000;
array[10619] <= 16'b0000_0000_0000_0000;
array[10620] <= 16'b0000_0000_0000_0000;
array[10621] <= 16'b0000_0000_0000_0000;
array[10622] <= 16'b0000_0000_0000_0000;
array[10623] <= 16'b0000_0000_0000_0000;
array[10624] <= 16'b0000_0000_0000_0000;
array[10625] <= 16'b0000_0000_0000_0000;
array[10626] <= 16'b0000_0000_0000_0000;
array[10627] <= 16'b0000_0000_0000_0000;
array[10628] <= 16'b0000_0000_0000_0000;
array[10629] <= 16'b0000_0000_0000_0000;
array[10630] <= 16'b0000_0000_0000_0000;
array[10631] <= 16'b0000_0000_0000_0000;
array[10632] <= 16'b0000_0000_0000_0000;
array[10633] <= 16'b0000_0000_0000_0000;
array[10634] <= 16'b0000_0000_0000_0000;
array[10635] <= 16'b0000_0000_0000_0000;
array[10636] <= 16'b0000_0000_0000_0000;
array[10637] <= 16'b0000_0000_0000_0000;
array[10638] <= 16'b0000_0000_0000_0000;
array[10639] <= 16'b0000_0000_0000_0000;
array[10640] <= 16'b0000_0000_0000_0000;
array[10641] <= 16'b0000_0000_0000_0000;
array[10642] <= 16'b0000_0000_0000_0000;
array[10643] <= 16'b0000_0000_0000_0000;
array[10644] <= 16'b0000_0000_0000_0000;
array[10645] <= 16'b0000_0000_0000_0000;
array[10646] <= 16'b0000_0000_0000_0000;
array[10647] <= 16'b0000_0000_0000_0000;
array[10648] <= 16'b0000_0000_0000_0000;
array[10649] <= 16'b0000_0000_0000_0000;
array[10650] <= 16'b0000_0000_0000_0000;
array[10651] <= 16'b0000_0000_0000_0000;
array[10652] <= 16'b0000_0000_0000_0000;
array[10653] <= 16'b0000_0000_0000_0000;
array[10654] <= 16'b0000_0000_0000_0000;
array[10655] <= 16'b0000_0000_0000_0000;
array[10656] <= 16'b0000_0000_0000_0000;
array[10657] <= 16'b0000_0000_0000_0000;
array[10658] <= 16'b0000_0000_0000_0000;
array[10659] <= 16'b0000_0000_0000_0000;
array[10660] <= 16'b0000_0000_0000_0000;
array[10661] <= 16'b0000_0000_0000_0000;
array[10662] <= 16'b0000_0000_0000_0000;
array[10663] <= 16'b0000_0000_0000_0000;
array[10664] <= 16'b0000_0000_0000_0000;
array[10665] <= 16'b0000_0000_0000_0000;
array[10666] <= 16'b0000_0000_0000_0000;
array[10667] <= 16'b0000_0000_0000_0000;
array[10668] <= 16'b0000_0000_0000_0000;
array[10669] <= 16'b0000_0000_0000_0000;
array[10670] <= 16'b0000_0000_0000_0000;
array[10671] <= 16'b0000_0000_0000_0000;
array[10672] <= 16'b0000_0000_0000_0000;
array[10673] <= 16'b0000_0000_0000_0000;
array[10674] <= 16'b0000_0000_0000_0000;
array[10675] <= 16'b0000_0000_0000_0000;
array[10676] <= 16'b0000_0000_0000_0000;
array[10677] <= 16'b0000_0000_0000_0000;
array[10678] <= 16'b0000_0000_0000_0000;
array[10679] <= 16'b0000_0000_0000_0000;
array[10680] <= 16'b0000_0000_0000_0000;
array[10681] <= 16'b0000_0000_0000_0000;
array[10682] <= 16'b0000_0000_0000_0000;
array[10683] <= 16'b0000_0000_0000_0000;
array[10684] <= 16'b0000_0000_0000_0000;
array[10685] <= 16'b0000_0000_0000_0000;
array[10686] <= 16'b0000_0000_0000_0000;
array[10687] <= 16'b0000_0000_0000_0000;
array[10688] <= 16'b0000_0000_0000_0000;
array[10689] <= 16'b0000_0000_0000_0000;
array[10690] <= 16'b0000_0000_0000_0000;
array[10691] <= 16'b0000_0000_0000_0000;
array[10692] <= 16'b0000_0000_0000_0000;
array[10693] <= 16'b0000_0000_0000_0000;
array[10694] <= 16'b0000_0000_0000_0000;
array[10695] <= 16'b0000_0000_0000_0000;
array[10696] <= 16'b0000_0000_0000_0000;
array[10697] <= 16'b0000_0000_0000_0000;
array[10698] <= 16'b0000_0000_0000_0000;
array[10699] <= 16'b0000_0000_0000_0000;
array[10700] <= 16'b0000_0000_0000_0000;
array[10701] <= 16'b0000_0000_0000_0000;
array[10702] <= 16'b0000_0000_0000_0000;
array[10703] <= 16'b0000_0000_0000_0000;
array[10704] <= 16'b0000_0000_0000_0000;
array[10705] <= 16'b0000_0000_0000_0000;
array[10706] <= 16'b0000_0000_0000_0000;
array[10707] <= 16'b0000_0000_0000_0000;
array[10708] <= 16'b0000_0000_0000_0000;
array[10709] <= 16'b0000_0000_0000_0000;
array[10710] <= 16'b0000_0000_0000_0000;
array[10711] <= 16'b0000_0000_0000_0000;
array[10712] <= 16'b0000_0000_0000_0000;
array[10713] <= 16'b0000_0000_0000_0000;
array[10714] <= 16'b0000_0000_0000_0000;
array[10715] <= 16'b0000_0000_0000_0000;
array[10716] <= 16'b0000_0000_0000_0000;
array[10717] <= 16'b0000_0000_0000_0000;
array[10718] <= 16'b0000_0000_0000_0000;
array[10719] <= 16'b0000_0000_0000_0000;
array[10720] <= 16'b0000_0000_0000_0000;
array[10721] <= 16'b0000_0000_0000_0000;
array[10722] <= 16'b0000_0000_0000_0000;
array[10723] <= 16'b0000_0000_0000_0000;
array[10724] <= 16'b0000_0000_0000_0000;
array[10725] <= 16'b0000_0000_0000_0000;
array[10726] <= 16'b0000_0000_0000_0000;
array[10727] <= 16'b0000_0000_0000_0000;
array[10728] <= 16'b0000_0000_0000_0000;
array[10729] <= 16'b0000_0000_0000_0000;
array[10730] <= 16'b0000_0000_0000_0000;
array[10731] <= 16'b0000_0000_0000_0000;
array[10732] <= 16'b0000_0000_0000_0000;
array[10733] <= 16'b0000_0000_0000_0000;
array[10734] <= 16'b0000_0000_0000_0000;
array[10735] <= 16'b0000_0000_0000_0000;
array[10736] <= 16'b0000_0000_0000_0000;
array[10737] <= 16'b0000_0000_0000_0000;
array[10738] <= 16'b0000_0000_0000_0000;
array[10739] <= 16'b0000_0000_0000_0000;
array[10740] <= 16'b0000_0000_0000_0000;
array[10741] <= 16'b0000_0000_0000_0000;
array[10742] <= 16'b0000_0000_0000_0000;
array[10743] <= 16'b0000_0000_0000_0000;
array[10744] <= 16'b0000_0000_0000_0000;
array[10745] <= 16'b0000_0000_0000_0000;
array[10746] <= 16'b0000_0000_0000_0000;
array[10747] <= 16'b0000_0000_0000_0000;
array[10748] <= 16'b0000_0000_0000_0000;
array[10749] <= 16'b0000_0000_0000_0000;
array[10750] <= 16'b0000_0000_0000_0000;
array[10751] <= 16'b0000_0000_0000_0000;
array[10752] <= 16'b0000_0000_0000_0000;
array[10753] <= 16'b0000_0000_0000_0000;
array[10754] <= 16'b0000_0000_0000_0000;
array[10755] <= 16'b0000_0000_0000_0000;
array[10756] <= 16'b0000_0000_0000_0000;
array[10757] <= 16'b0000_0000_0000_0000;
array[10758] <= 16'b0000_0000_0000_0000;
array[10759] <= 16'b0000_0000_0000_0000;
array[10760] <= 16'b0000_0000_0000_0000;
array[10761] <= 16'b0000_0000_0000_0000;
array[10762] <= 16'b0000_0000_0000_0000;
array[10763] <= 16'b0000_0000_0000_0000;
array[10764] <= 16'b0000_0000_0000_0000;
array[10765] <= 16'b0000_0000_0000_0000;
array[10766] <= 16'b0000_0000_0000_0000;
array[10767] <= 16'b0000_0000_0000_0000;
array[10768] <= 16'b0000_0000_0000_0000;
array[10769] <= 16'b0000_0000_0000_0000;
array[10770] <= 16'b0000_0000_0000_0000;
array[10771] <= 16'b0000_0000_0000_0000;
array[10772] <= 16'b0000_0000_0000_0000;
array[10773] <= 16'b0000_0000_0000_0000;
array[10774] <= 16'b0000_0000_0000_0000;
array[10775] <= 16'b0000_0000_0000_0000;
array[10776] <= 16'b0000_0000_0000_0000;
array[10777] <= 16'b0000_0000_0000_0000;
array[10778] <= 16'b0000_0000_0000_0000;
array[10779] <= 16'b0000_0000_0000_0000;
array[10780] <= 16'b0000_0000_0000_0000;
array[10781] <= 16'b0000_0000_0000_0000;
array[10782] <= 16'b0000_0000_0000_0000;
array[10783] <= 16'b0000_0000_0000_0000;
array[10784] <= 16'b0000_0000_0000_0000;
array[10785] <= 16'b0000_0000_0000_0000;
array[10786] <= 16'b0000_0000_0000_0000;
array[10787] <= 16'b0000_0000_0000_0000;
array[10788] <= 16'b0000_0000_0000_0000;
array[10789] <= 16'b0000_0000_0000_0000;
array[10790] <= 16'b0000_0000_0000_0000;
array[10791] <= 16'b0000_0000_0000_0000;
array[10792] <= 16'b0000_0000_0000_0000;
array[10793] <= 16'b0000_0000_0000_0000;
array[10794] <= 16'b0000_0000_0000_0000;
array[10795] <= 16'b0000_0000_0000_0000;
array[10796] <= 16'b0000_0000_0000_0000;
array[10797] <= 16'b0000_0000_0000_0000;
array[10798] <= 16'b0000_0000_0000_0000;
array[10799] <= 16'b0000_0000_0000_0000;
array[10800] <= 16'b0000_0000_0000_0000;
array[10801] <= 16'b0000_0000_0000_0000;
array[10802] <= 16'b0000_0000_0000_0000;
array[10803] <= 16'b0000_0000_0000_0000;
array[10804] <= 16'b0000_0000_0000_0000;
array[10805] <= 16'b0000_0000_0000_0000;
array[10806] <= 16'b0000_0000_0000_0000;
array[10807] <= 16'b0000_0000_0000_0000;
array[10808] <= 16'b0000_0000_0000_0000;
array[10809] <= 16'b0000_0000_0000_0000;
array[10810] <= 16'b0000_0000_0000_0000;
array[10811] <= 16'b0000_0000_0000_0000;
array[10812] <= 16'b0000_0000_0000_0000;
array[10813] <= 16'b0000_0000_0000_0000;
array[10814] <= 16'b0000_0000_0000_0000;
array[10815] <= 16'b0000_0000_0000_0000;
array[10816] <= 16'b0000_0000_0000_0000;
array[10817] <= 16'b0000_0000_0000_0000;
array[10818] <= 16'b0000_0000_0000_0000;
array[10819] <= 16'b0000_0000_0000_0000;
array[10820] <= 16'b0000_0000_0000_0000;
array[10821] <= 16'b0000_0000_0000_0000;
array[10822] <= 16'b0000_0000_0000_0000;
array[10823] <= 16'b0000_0000_0000_0000;
array[10824] <= 16'b0000_0000_0000_0000;
array[10825] <= 16'b0000_0000_0000_0000;
array[10826] <= 16'b0000_0000_0000_0000;
array[10827] <= 16'b0000_0000_0000_0000;
array[10828] <= 16'b0000_0000_0000_0000;
array[10829] <= 16'b0000_0000_0000_0000;
array[10830] <= 16'b0000_0000_0000_0000;
array[10831] <= 16'b0000_0000_0000_0000;
array[10832] <= 16'b0000_0000_0000_0000;
array[10833] <= 16'b0000_0000_0000_0000;
array[10834] <= 16'b0000_0000_0000_0000;
array[10835] <= 16'b0000_0000_0000_0000;
array[10836] <= 16'b0000_0000_0000_0000;
array[10837] <= 16'b0000_0000_0000_0000;
array[10838] <= 16'b0000_0000_0000_0000;
array[10839] <= 16'b0000_0000_0000_0000;
array[10840] <= 16'b0000_0000_0000_0000;
array[10841] <= 16'b0000_0000_0000_0000;
array[10842] <= 16'b0000_0000_0000_0000;
array[10843] <= 16'b0000_0000_0000_0000;
array[10844] <= 16'b0000_0000_0000_0000;
array[10845] <= 16'b0000_0000_0000_0000;
array[10846] <= 16'b0000_0000_0000_0000;
array[10847] <= 16'b0000_0000_0000_0000;
array[10848] <= 16'b0000_0000_0000_0000;
array[10849] <= 16'b0000_0000_0000_0000;
array[10850] <= 16'b0000_0000_0000_0000;
array[10851] <= 16'b0000_0000_0000_0000;
array[10852] <= 16'b0000_0000_0000_0000;
array[10853] <= 16'b0000_0000_0000_0000;
array[10854] <= 16'b0000_0000_0000_0000;
array[10855] <= 16'b0000_0000_0000_0000;
array[10856] <= 16'b0000_0000_0000_0000;
array[10857] <= 16'b0000_0000_0000_0000;
array[10858] <= 16'b0000_0000_0000_0000;
array[10859] <= 16'b0000_0000_0000_0000;
array[10860] <= 16'b0000_0000_0000_0000;
array[10861] <= 16'b0000_0000_0000_0000;
array[10862] <= 16'b0000_0000_0000_0000;
array[10863] <= 16'b0000_0000_0000_0000;
array[10864] <= 16'b0000_0000_0000_0000;
array[10865] <= 16'b0000_0000_0000_0000;
array[10866] <= 16'b0000_0000_0000_0000;
array[10867] <= 16'b0000_0000_0000_0000;
array[10868] <= 16'b0000_0000_0000_0000;
array[10869] <= 16'b0000_0000_0000_0000;
array[10870] <= 16'b0000_0000_0000_0000;
array[10871] <= 16'b0000_0000_0000_0000;
array[10872] <= 16'b0000_0000_0000_0000;
array[10873] <= 16'b0000_0000_0000_0000;
array[10874] <= 16'b0000_0000_0000_0000;
array[10875] <= 16'b0000_0000_0000_0000;
array[10876] <= 16'b0000_0000_0000_0000;
array[10877] <= 16'b0000_0000_0000_0000;
array[10878] <= 16'b0000_0000_0000_0000;
array[10879] <= 16'b0000_0000_0000_0000;
array[10880] <= 16'b0000_0000_0000_0000;
array[10881] <= 16'b0000_0000_0000_0000;
array[10882] <= 16'b0000_0000_0000_0000;
array[10883] <= 16'b0000_0000_0000_0000;
array[10884] <= 16'b0000_0000_0000_0000;
array[10885] <= 16'b0000_0000_0000_0000;
array[10886] <= 16'b0000_0000_0000_0000;
array[10887] <= 16'b0000_0000_0000_0000;
array[10888] <= 16'b0000_0000_0000_0000;
array[10889] <= 16'b0000_0000_0000_0000;
array[10890] <= 16'b0000_0000_0000_0000;
array[10891] <= 16'b0000_0000_0000_0000;
array[10892] <= 16'b0000_0000_0000_0000;
array[10893] <= 16'b0000_0000_0000_0000;
array[10894] <= 16'b0000_0000_0000_0000;
array[10895] <= 16'b0000_0000_0000_0000;
array[10896] <= 16'b0000_0000_0000_0000;
array[10897] <= 16'b0000_0000_0000_0000;
array[10898] <= 16'b0000_0000_0000_0000;
array[10899] <= 16'b0000_0000_0000_0000;
array[10900] <= 16'b0000_0000_0000_0000;
array[10901] <= 16'b0000_0000_0000_0000;
array[10902] <= 16'b0000_0000_0000_0000;
array[10903] <= 16'b0000_0000_0000_0000;
array[10904] <= 16'b0000_0000_0000_0000;
array[10905] <= 16'b0000_0000_0000_0000;
array[10906] <= 16'b0000_0000_0000_0000;
array[10907] <= 16'b0000_0000_0000_0000;
array[10908] <= 16'b0000_0000_0000_0000;
array[10909] <= 16'b0000_0000_0000_0000;
array[10910] <= 16'b0000_0000_0000_0000;
array[10911] <= 16'b0000_0000_0000_0000;
array[10912] <= 16'b0000_0000_0000_0000;
array[10913] <= 16'b0000_0000_0000_0000;
array[10914] <= 16'b0000_0000_0000_0000;
array[10915] <= 16'b0000_0000_0000_0000;
array[10916] <= 16'b0000_0000_0000_0000;
array[10917] <= 16'b0000_0000_0000_0000;
array[10918] <= 16'b0000_0000_0000_0000;
array[10919] <= 16'b0000_0000_0000_0000;
array[10920] <= 16'b0000_0000_0000_0000;
array[10921] <= 16'b0000_0000_0000_0000;
array[10922] <= 16'b0000_0000_0000_0000;
array[10923] <= 16'b0000_0000_0000_0000;
array[10924] <= 16'b0000_0000_0000_0000;
array[10925] <= 16'b0000_0000_0000_0000;
array[10926] <= 16'b0000_0000_0000_0000;
array[10927] <= 16'b0000_0000_0000_0000;
array[10928] <= 16'b0000_0000_0000_0000;
array[10929] <= 16'b0000_0000_0000_0000;
array[10930] <= 16'b0000_0000_0000_0000;
array[10931] <= 16'b0000_0000_0000_0000;
array[10932] <= 16'b0000_0000_0000_0000;
array[10933] <= 16'b0000_0000_0000_0000;
array[10934] <= 16'b0000_0000_0000_0000;
array[10935] <= 16'b0000_0000_0000_0000;
array[10936] <= 16'b0000_0000_0000_0000;
array[10937] <= 16'b0000_0000_0000_0000;
array[10938] <= 16'b0000_0000_0000_0000;
array[10939] <= 16'b0000_0000_0000_0000;
array[10940] <= 16'b0000_0000_0000_0000;
array[10941] <= 16'b0000_0000_0000_0000;
array[10942] <= 16'b0000_0000_0000_0000;
array[10943] <= 16'b0000_0000_0000_0000;
array[10944] <= 16'b0000_0000_0000_0000;
array[10945] <= 16'b0000_0000_0000_0000;
array[10946] <= 16'b0000_0000_0000_0000;
array[10947] <= 16'b0000_0000_0000_0000;
array[10948] <= 16'b0000_0000_0000_0000;
array[10949] <= 16'b0000_0000_0000_0000;
array[10950] <= 16'b0000_0000_0000_0000;
array[10951] <= 16'b0000_0000_0000_0000;
array[10952] <= 16'b0000_0000_0000_0000;
array[10953] <= 16'b0000_0000_0000_0000;
array[10954] <= 16'b0000_0000_0000_0000;
array[10955] <= 16'b0000_0000_0000_0000;
array[10956] <= 16'b0000_0000_0000_0000;
array[10957] <= 16'b0000_0000_0000_0000;
array[10958] <= 16'b0000_0000_0000_0000;
array[10959] <= 16'b0000_0000_0000_0000;
array[10960] <= 16'b0000_0000_0000_0000;
array[10961] <= 16'b0000_0000_0000_0000;
array[10962] <= 16'b0000_0000_0000_0000;
array[10963] <= 16'b0000_0000_0000_0000;
array[10964] <= 16'b0000_0000_0000_0000;
array[10965] <= 16'b0000_0000_0000_0000;
array[10966] <= 16'b0000_0000_0000_0000;
array[10967] <= 16'b0000_0000_0000_0000;
array[10968] <= 16'b0000_0000_0000_0000;
array[10969] <= 16'b0000_0000_0000_0000;
array[10970] <= 16'b0000_0000_0000_0000;
array[10971] <= 16'b0000_0000_0000_0000;
array[10972] <= 16'b0000_0000_0000_0000;
array[10973] <= 16'b0000_0000_0000_0000;
array[10974] <= 16'b0000_0000_0000_0000;
array[10975] <= 16'b0000_0000_0000_0000;
array[10976] <= 16'b0000_0000_0000_0000;
array[10977] <= 16'b0000_0000_0000_0000;
array[10978] <= 16'b0000_0000_0000_0000;
array[10979] <= 16'b0000_0000_0000_0000;
array[10980] <= 16'b0000_0000_0000_0000;
array[10981] <= 16'b0000_0000_0000_0000;
array[10982] <= 16'b0000_0000_0000_0000;
array[10983] <= 16'b0000_0000_0000_0000;
array[10984] <= 16'b0000_0000_0000_0000;
array[10985] <= 16'b0000_0000_0000_0000;
array[10986] <= 16'b0000_0000_0000_0000;
array[10987] <= 16'b0000_0000_0000_0000;
array[10988] <= 16'b0000_0000_0000_0000;
array[10989] <= 16'b0000_0000_0000_0000;
array[10990] <= 16'b0000_0000_0000_0000;
array[10991] <= 16'b0000_0000_0000_0000;
array[10992] <= 16'b0000_0000_0000_0000;
array[10993] <= 16'b0000_0000_0000_0000;
array[10994] <= 16'b0000_0000_0000_0000;
array[10995] <= 16'b0000_0000_0000_0000;
array[10996] <= 16'b0000_0000_0000_0000;
array[10997] <= 16'b0000_0000_0000_0000;
array[10998] <= 16'b0000_0000_0000_0000;
array[10999] <= 16'b0000_0000_0000_0000;
array[11000] <= 16'b0000_0000_0000_0000;
array[11001] <= 16'b0000_0000_0000_0000;
array[11002] <= 16'b0000_0000_0000_0000;
array[11003] <= 16'b0000_0000_0000_0000;
array[11004] <= 16'b0000_0000_0000_0000;
array[11005] <= 16'b0000_0000_0000_0000;
array[11006] <= 16'b0000_0000_0000_0000;
array[11007] <= 16'b0000_0000_0000_0000;
array[11008] <= 16'b0000_0000_0000_0000;
array[11009] <= 16'b0000_0000_0000_0000;
array[11010] <= 16'b0000_0000_0000_0000;
array[11011] <= 16'b0000_0000_0000_0000;
array[11012] <= 16'b0000_0000_0000_0000;
array[11013] <= 16'b0000_0000_0000_0000;
array[11014] <= 16'b0000_0000_0000_0000;
array[11015] <= 16'b0000_0000_0000_0000;
array[11016] <= 16'b0000_0000_0000_0000;
array[11017] <= 16'b0000_0000_0000_0000;
array[11018] <= 16'b0000_0000_0000_0000;
array[11019] <= 16'b0000_0000_0000_0000;
array[11020] <= 16'b0000_0000_0000_0000;
array[11021] <= 16'b0000_0000_0000_0000;
array[11022] <= 16'b0000_0000_0000_0000;
array[11023] <= 16'b0000_0000_0000_0000;
array[11024] <= 16'b0000_0000_0000_0000;
array[11025] <= 16'b0000_0000_0000_0000;
array[11026] <= 16'b0000_0000_0000_0000;
array[11027] <= 16'b0000_0000_0000_0000;
array[11028] <= 16'b0000_0000_0000_0000;
array[11029] <= 16'b0000_0000_0000_0000;
array[11030] <= 16'b0000_0000_0000_0000;
array[11031] <= 16'b0000_0000_0000_0000;
array[11032] <= 16'b0000_0000_0000_0000;
array[11033] <= 16'b0000_0000_0000_0000;
array[11034] <= 16'b0000_0000_0000_0000;
array[11035] <= 16'b0000_0000_0000_0000;
array[11036] <= 16'b0000_0000_0000_0000;
array[11037] <= 16'b0000_0000_0000_0000;
array[11038] <= 16'b0000_0000_0000_0000;
array[11039] <= 16'b0000_0000_0000_0000;
array[11040] <= 16'b0000_0000_0000_0000;
array[11041] <= 16'b0000_0000_0000_0000;
array[11042] <= 16'b0000_0000_0000_0000;
array[11043] <= 16'b0000_0000_0000_0000;
array[11044] <= 16'b0000_0000_0000_0000;
array[11045] <= 16'b0000_0000_0000_0000;
array[11046] <= 16'b0000_0000_0000_0000;
array[11047] <= 16'b0000_0000_0000_0000;
array[11048] <= 16'b0000_0000_0000_0000;
array[11049] <= 16'b0000_0000_0000_0000;
array[11050] <= 16'b0000_0000_0000_0000;
array[11051] <= 16'b0000_0000_0000_0000;
array[11052] <= 16'b0000_0000_0000_0000;
array[11053] <= 16'b0000_0000_0000_0000;
array[11054] <= 16'b0000_0000_0000_0000;
array[11055] <= 16'b0000_0000_0000_0000;
array[11056] <= 16'b0000_0000_0000_0000;
array[11057] <= 16'b0000_0000_0000_0000;
array[11058] <= 16'b0000_0000_0000_0000;
array[11059] <= 16'b0000_0000_0000_0000;
array[11060] <= 16'b0000_0000_0000_0000;
array[11061] <= 16'b0000_0000_0000_0000;
array[11062] <= 16'b0000_0000_0000_0000;
array[11063] <= 16'b0000_0000_0000_0000;
array[11064] <= 16'b0000_0000_0000_0000;
array[11065] <= 16'b0000_0000_0000_0000;
array[11066] <= 16'b0000_0000_0000_0000;
array[11067] <= 16'b0000_0000_0000_0000;
array[11068] <= 16'b0000_0000_0000_0000;
array[11069] <= 16'b0000_0000_0000_0000;
array[11070] <= 16'b0000_0000_0000_0000;
array[11071] <= 16'b0000_0000_0000_0000;
array[11072] <= 16'b0000_0000_0000_0000;
array[11073] <= 16'b0000_0000_0000_0000;
array[11074] <= 16'b0000_0000_0000_0000;
array[11075] <= 16'b0000_0000_0000_0000;
array[11076] <= 16'b0000_0000_0000_0000;
array[11077] <= 16'b0000_0000_0000_0000;
array[11078] <= 16'b0000_0000_0000_0000;
array[11079] <= 16'b0000_0000_0000_0000;
array[11080] <= 16'b0000_0000_0000_0000;
array[11081] <= 16'b0000_0000_0000_0000;
array[11082] <= 16'b0000_0000_0000_0000;
array[11083] <= 16'b0000_0000_0000_0000;
array[11084] <= 16'b0000_0000_0000_0000;
array[11085] <= 16'b0000_0000_0000_0000;
array[11086] <= 16'b0000_0000_0000_0000;
array[11087] <= 16'b0000_0000_0000_0000;
array[11088] <= 16'b0000_0000_0000_0000;
array[11089] <= 16'b0000_0000_0000_0000;
array[11090] <= 16'b0000_0000_0000_0000;
array[11091] <= 16'b0000_0000_0000_0000;
array[11092] <= 16'b0000_0000_0000_0000;
array[11093] <= 16'b0000_0000_0000_0000;
array[11094] <= 16'b0000_0000_0000_0000;
array[11095] <= 16'b0000_0000_0000_0000;
array[11096] <= 16'b0000_0000_0000_0000;
array[11097] <= 16'b0000_0000_0000_0000;
array[11098] <= 16'b0000_0000_0000_0000;
array[11099] <= 16'b0000_0000_0000_0000;
array[11100] <= 16'b0000_0000_0000_0000;
array[11101] <= 16'b0000_0000_0000_0000;
array[11102] <= 16'b0000_0000_0000_0000;
array[11103] <= 16'b0000_0000_0000_0000;
array[11104] <= 16'b0000_0000_0000_0000;
array[11105] <= 16'b0000_0000_0000_0000;
array[11106] <= 16'b0000_0000_0000_0000;
array[11107] <= 16'b0000_0000_0000_0000;
array[11108] <= 16'b0000_0000_0000_0000;
array[11109] <= 16'b0000_0000_0000_0000;
array[11110] <= 16'b0000_0000_0000_0000;
array[11111] <= 16'b0000_0000_0000_0000;
array[11112] <= 16'b0000_0000_0000_0000;
array[11113] <= 16'b0000_0000_0000_0000;
array[11114] <= 16'b0000_0000_0000_0000;
array[11115] <= 16'b0000_0000_0000_0000;
array[11116] <= 16'b0000_0000_0000_0000;
array[11117] <= 16'b0000_0000_0000_0000;
array[11118] <= 16'b0000_0000_0000_0000;
array[11119] <= 16'b0000_0000_0000_0000;
array[11120] <= 16'b0000_0000_0000_0000;
array[11121] <= 16'b0000_0000_0000_0000;
array[11122] <= 16'b0000_0000_0000_0000;
array[11123] <= 16'b0000_0000_0000_0000;
array[11124] <= 16'b0000_0000_0000_0000;
array[11125] <= 16'b0000_0000_0000_0000;
array[11126] <= 16'b0000_0000_0000_0000;
array[11127] <= 16'b0000_0000_0000_0000;
array[11128] <= 16'b0000_0000_0000_0000;
array[11129] <= 16'b0000_0000_0000_0000;
array[11130] <= 16'b0000_0000_0000_0000;
array[11131] <= 16'b0000_0000_0000_0000;
array[11132] <= 16'b0000_0000_0000_0000;
array[11133] <= 16'b0000_0000_0000_0000;
array[11134] <= 16'b0000_0000_0000_0000;
array[11135] <= 16'b0000_0000_0000_0000;
array[11136] <= 16'b0000_0000_0000_0000;
array[11137] <= 16'b0000_0000_0000_0000;
array[11138] <= 16'b0000_0000_0000_0000;
array[11139] <= 16'b0000_0000_0000_0000;
array[11140] <= 16'b0000_0000_0000_0000;
array[11141] <= 16'b0000_0000_0000_0000;
array[11142] <= 16'b0000_0000_0000_0000;
array[11143] <= 16'b0000_0000_0000_0000;
array[11144] <= 16'b0000_0000_0000_0000;
array[11145] <= 16'b0000_0000_0000_0000;
array[11146] <= 16'b0000_0000_0000_0000;
array[11147] <= 16'b0000_0000_0000_0000;
array[11148] <= 16'b0000_0000_0000_0000;
array[11149] <= 16'b0000_0000_0000_0000;
array[11150] <= 16'b0000_0000_0000_0000;
array[11151] <= 16'b0000_0000_0000_0000;
array[11152] <= 16'b0000_0000_0000_0000;
array[11153] <= 16'b0000_0000_0000_0000;
array[11154] <= 16'b0000_0000_0000_0000;
array[11155] <= 16'b0000_0000_0000_0000;
array[11156] <= 16'b0000_0000_0000_0000;
array[11157] <= 16'b0000_0000_0000_0000;
array[11158] <= 16'b0000_0000_0000_0000;
array[11159] <= 16'b0000_0000_0000_0000;
array[11160] <= 16'b0000_0000_0000_0000;
array[11161] <= 16'b0000_0000_0000_0000;
array[11162] <= 16'b0000_0000_0000_0000;
array[11163] <= 16'b0000_0000_0000_0000;
array[11164] <= 16'b0000_0000_0000_0000;
array[11165] <= 16'b0000_0000_0000_0000;
array[11166] <= 16'b0000_0000_0000_0000;
array[11167] <= 16'b0000_0000_0000_0000;
array[11168] <= 16'b0000_0000_0000_0000;
array[11169] <= 16'b0000_0000_0000_0000;
array[11170] <= 16'b0000_0000_0000_0000;
array[11171] <= 16'b0000_0000_0000_0000;
array[11172] <= 16'b0000_0000_0000_0000;
array[11173] <= 16'b0000_0000_0000_0000;
array[11174] <= 16'b0000_0000_0000_0000;
array[11175] <= 16'b0000_0000_0000_0000;
array[11176] <= 16'b0000_0000_0000_0000;
array[11177] <= 16'b0000_0000_0000_0000;
array[11178] <= 16'b0000_0000_0000_0000;
array[11179] <= 16'b0000_0000_0000_0000;
array[11180] <= 16'b0000_0000_0000_0000;
array[11181] <= 16'b0000_0000_0000_0000;
array[11182] <= 16'b0000_0000_0000_0000;
array[11183] <= 16'b0000_0000_0000_0000;
array[11184] <= 16'b0000_0000_0000_0000;
array[11185] <= 16'b0000_0000_0000_0000;
array[11186] <= 16'b0000_0000_0000_0000;
array[11187] <= 16'b0000_0000_0000_0000;
array[11188] <= 16'b0000_0000_0000_0000;
array[11189] <= 16'b0000_0000_0000_0000;
array[11190] <= 16'b0000_0000_0000_0000;
array[11191] <= 16'b0000_0000_0000_0000;
array[11192] <= 16'b0000_0000_0000_0000;
array[11193] <= 16'b0000_0000_0000_0000;
array[11194] <= 16'b0000_0000_0000_0000;
array[11195] <= 16'b0000_0000_0000_0000;
array[11196] <= 16'b0000_0000_0000_0000;
array[11197] <= 16'b0000_0000_0000_0000;
array[11198] <= 16'b0000_0000_0000_0000;
array[11199] <= 16'b0000_0000_0000_0000;
array[11200] <= 16'b0000_0000_0000_0000;
array[11201] <= 16'b0000_0000_0000_0000;
array[11202] <= 16'b0000_0000_0000_0000;
array[11203] <= 16'b0000_0000_0000_0000;
array[11204] <= 16'b0000_0000_0000_0000;
array[11205] <= 16'b0000_0000_0000_0000;
array[11206] <= 16'b0000_0000_0000_0000;
array[11207] <= 16'b0000_0000_0000_0000;
array[11208] <= 16'b0000_0000_0000_0000;
array[11209] <= 16'b0000_0000_0000_0000;
array[11210] <= 16'b0000_0000_0000_0000;
array[11211] <= 16'b0000_0000_0000_0000;
array[11212] <= 16'b0000_0000_0000_0000;
array[11213] <= 16'b0000_0000_0000_0000;
array[11214] <= 16'b0000_0000_0000_0000;
array[11215] <= 16'b0000_0000_0000_0000;
array[11216] <= 16'b0000_0000_0000_0000;
array[11217] <= 16'b0000_0000_0000_0000;
array[11218] <= 16'b0000_0000_0000_0000;
array[11219] <= 16'b0000_0000_0000_0000;
array[11220] <= 16'b0000_0000_0000_0000;
array[11221] <= 16'b0000_0000_0000_0000;
array[11222] <= 16'b0000_0000_0000_0000;
array[11223] <= 16'b0000_0000_0000_0000;
array[11224] <= 16'b0000_0000_0000_0000;
array[11225] <= 16'b0000_0000_0000_0000;
array[11226] <= 16'b0000_0000_0000_0000;
array[11227] <= 16'b0000_0000_0000_0000;
array[11228] <= 16'b0000_0000_0000_0000;
array[11229] <= 16'b0000_0000_0000_0000;
array[11230] <= 16'b0000_0000_0000_0000;
array[11231] <= 16'b0000_0000_0000_0000;
array[11232] <= 16'b0000_0000_0000_0000;
array[11233] <= 16'b0000_0000_0000_0000;
array[11234] <= 16'b0000_0000_0000_0000;
array[11235] <= 16'b0000_0000_0000_0000;
array[11236] <= 16'b0000_0000_0000_0000;
array[11237] <= 16'b0000_0000_0000_0000;
array[11238] <= 16'b0000_0000_0000_0000;
array[11239] <= 16'b0000_0000_0000_0000;
array[11240] <= 16'b0000_0000_0000_0000;
array[11241] <= 16'b0000_0000_0000_0000;
array[11242] <= 16'b0000_0000_0000_0000;
array[11243] <= 16'b0000_0000_0000_0000;
array[11244] <= 16'b0000_0000_0000_0000;
array[11245] <= 16'b0000_0000_0000_0000;
array[11246] <= 16'b0000_0000_0000_0000;
array[11247] <= 16'b0000_0000_0000_0000;
array[11248] <= 16'b0000_0000_0000_0000;
array[11249] <= 16'b0000_0000_0000_0000;
array[11250] <= 16'b0000_0000_0000_0000;
array[11251] <= 16'b0000_0000_0000_0000;
array[11252] <= 16'b0000_0000_0000_0000;
array[11253] <= 16'b0000_0000_0000_0000;
array[11254] <= 16'b0000_0000_0000_0000;
array[11255] <= 16'b0000_0000_0000_0000;
array[11256] <= 16'b0000_0000_0000_0000;
array[11257] <= 16'b0000_0000_0000_0000;
array[11258] <= 16'b0000_0000_0000_0000;
array[11259] <= 16'b0000_0000_0000_0000;
array[11260] <= 16'b0000_0000_0000_0000;
array[11261] <= 16'b0000_0000_0000_0000;
array[11262] <= 16'b0000_0000_0000_0000;
array[11263] <= 16'b0000_0000_0000_0000;
array[11264] <= 16'b0000_0000_0000_0000;
array[11265] <= 16'b0000_0000_0000_0000;
array[11266] <= 16'b0000_0000_0000_0000;
array[11267] <= 16'b0000_0000_0000_0000;
array[11268] <= 16'b0000_0000_0000_0000;
array[11269] <= 16'b0000_0000_0000_0000;
array[11270] <= 16'b0000_0000_0000_0000;
array[11271] <= 16'b0000_0000_0000_0000;
array[11272] <= 16'b0000_0000_0000_0000;
array[11273] <= 16'b0000_0000_0000_0000;
array[11274] <= 16'b0000_0000_0000_0000;
array[11275] <= 16'b0000_0000_0000_0000;
array[11276] <= 16'b0000_0000_0000_0000;
array[11277] <= 16'b0000_0000_0000_0000;
array[11278] <= 16'b0000_0000_0000_0000;
array[11279] <= 16'b0000_0000_0000_0000;
array[11280] <= 16'b0000_0000_0000_0000;
array[11281] <= 16'b0000_0000_0000_0000;
array[11282] <= 16'b0000_0000_0000_0000;
array[11283] <= 16'b0000_0000_0000_0000;
array[11284] <= 16'b0000_0000_0000_0000;
array[11285] <= 16'b0000_0000_0000_0000;
array[11286] <= 16'b0000_0000_0000_0000;
array[11287] <= 16'b0000_0000_0000_0000;
array[11288] <= 16'b0000_0000_0000_0000;
array[11289] <= 16'b0000_0000_0000_0000;
array[11290] <= 16'b0000_0000_0000_0000;
array[11291] <= 16'b0000_0000_0000_0000;
array[11292] <= 16'b0000_0000_0000_0000;
array[11293] <= 16'b0000_0000_0000_0000;
array[11294] <= 16'b0000_0000_0000_0000;
array[11295] <= 16'b0000_0000_0000_0000;
array[11296] <= 16'b0000_0000_0000_0000;
array[11297] <= 16'b0000_0000_0000_0000;
array[11298] <= 16'b0000_0000_0000_0000;
array[11299] <= 16'b0000_0000_0000_0000;
array[11300] <= 16'b0000_0000_0000_0000;
array[11301] <= 16'b0000_0000_0000_0000;
array[11302] <= 16'b0000_0000_0000_0000;
array[11303] <= 16'b0000_0000_0000_0000;
array[11304] <= 16'b0000_0000_0000_0000;
array[11305] <= 16'b0000_0000_0000_0000;
array[11306] <= 16'b0000_0000_0000_0000;
array[11307] <= 16'b0000_0000_0000_0000;
array[11308] <= 16'b0000_0000_0000_0000;
array[11309] <= 16'b0000_0000_0000_0000;
array[11310] <= 16'b0000_0000_0000_0000;
array[11311] <= 16'b0000_0000_0000_0000;
array[11312] <= 16'b0000_0000_0000_0000;
array[11313] <= 16'b0000_0000_0000_0000;
array[11314] <= 16'b0000_0000_0000_0000;
array[11315] <= 16'b0000_0000_0000_0000;
array[11316] <= 16'b0000_0000_0000_0000;
array[11317] <= 16'b0000_0000_0000_0000;
array[11318] <= 16'b0000_0000_0000_0000;
array[11319] <= 16'b0000_0000_0000_0000;
array[11320] <= 16'b0000_0000_0000_0000;
array[11321] <= 16'b0000_0000_0000_0000;
array[11322] <= 16'b0000_0000_0000_0000;
array[11323] <= 16'b0000_0000_0000_0000;
array[11324] <= 16'b0000_0000_0000_0000;
array[11325] <= 16'b0000_0000_0000_0000;
array[11326] <= 16'b0000_0000_0000_0000;
array[11327] <= 16'b0000_0000_0000_0000;
array[11328] <= 16'b0000_0000_0000_0000;
array[11329] <= 16'b0000_0000_0000_0000;
array[11330] <= 16'b0000_0000_0000_0000;
array[11331] <= 16'b0000_0000_0000_0000;
array[11332] <= 16'b0000_0000_0000_0000;
array[11333] <= 16'b0000_0000_0000_0000;
array[11334] <= 16'b0000_0000_0000_0000;
array[11335] <= 16'b0000_0000_0000_0000;
array[11336] <= 16'b0000_0000_0000_0000;
array[11337] <= 16'b0000_0000_0000_0000;
array[11338] <= 16'b0000_0000_0000_0000;
array[11339] <= 16'b0000_0000_0000_0000;
array[11340] <= 16'b0000_0000_0000_0000;
array[11341] <= 16'b0000_0000_0000_0000;
array[11342] <= 16'b0000_0000_0000_0000;
array[11343] <= 16'b0000_0000_0000_0000;
array[11344] <= 16'b0000_0000_0000_0000;
array[11345] <= 16'b0000_0000_0000_0000;
array[11346] <= 16'b0000_0000_0000_0000;
array[11347] <= 16'b0000_0000_0000_0000;
array[11348] <= 16'b0000_0000_0000_0000;
array[11349] <= 16'b0000_0000_0000_0000;
array[11350] <= 16'b0000_0000_0000_0000;
array[11351] <= 16'b0000_0000_0000_0000;
array[11352] <= 16'b0000_0000_0000_0000;
array[11353] <= 16'b0000_0000_0000_0000;
array[11354] <= 16'b0000_0000_0000_0000;
array[11355] <= 16'b0000_0000_0000_0000;
array[11356] <= 16'b0000_0000_0000_0000;
array[11357] <= 16'b0000_0000_0000_0000;
array[11358] <= 16'b0000_0000_0000_0000;
array[11359] <= 16'b0000_0000_0000_0000;
array[11360] <= 16'b0000_0000_0000_0000;
array[11361] <= 16'b0000_0000_0000_0000;
array[11362] <= 16'b0000_0000_0000_0000;
array[11363] <= 16'b0000_0000_0000_0000;
array[11364] <= 16'b0000_0000_0000_0000;
array[11365] <= 16'b0000_0000_0000_0000;
array[11366] <= 16'b0000_0000_0000_0000;
array[11367] <= 16'b0000_0000_0000_0000;
array[11368] <= 16'b0000_0000_0000_0000;
array[11369] <= 16'b0000_0000_0000_0000;
array[11370] <= 16'b0000_0000_0000_0000;
array[11371] <= 16'b0000_0000_0000_0000;
array[11372] <= 16'b0000_0000_0000_0000;
array[11373] <= 16'b0000_0000_0000_0000;
array[11374] <= 16'b0000_0000_0000_0000;
array[11375] <= 16'b0000_0000_0000_0000;
array[11376] <= 16'b0000_0000_0000_0000;
array[11377] <= 16'b0000_0000_0000_0000;
array[11378] <= 16'b0000_0000_0000_0000;
array[11379] <= 16'b0000_0000_0000_0000;
array[11380] <= 16'b0000_0000_0000_0000;
array[11381] <= 16'b0000_0000_0000_0000;
array[11382] <= 16'b0000_0000_0000_0000;
array[11383] <= 16'b0000_0000_0000_0000;
array[11384] <= 16'b0000_0000_0000_0000;
array[11385] <= 16'b0000_0000_0000_0000;
array[11386] <= 16'b0000_0000_0000_0000;
array[11387] <= 16'b0000_0000_0000_0000;
array[11388] <= 16'b0000_0000_0000_0000;
array[11389] <= 16'b0000_0000_0000_0000;
array[11390] <= 16'b0000_0000_0000_0000;
array[11391] <= 16'b0000_0000_0000_0000;
array[11392] <= 16'b0000_0000_0000_0000;
array[11393] <= 16'b0000_0000_0000_0000;
array[11394] <= 16'b0000_0000_0000_0000;
array[11395] <= 16'b0000_0000_0000_0000;
array[11396] <= 16'b0000_0000_0000_0000;
array[11397] <= 16'b0000_0000_0000_0000;
array[11398] <= 16'b0000_0000_0000_0000;
array[11399] <= 16'b0000_0000_0000_0000;
array[11400] <= 16'b0000_0000_0000_0000;
array[11401] <= 16'b0000_0000_0000_0000;
array[11402] <= 16'b0000_0000_0000_0000;
array[11403] <= 16'b0000_0000_0000_0000;
array[11404] <= 16'b0000_0000_0000_0000;
array[11405] <= 16'b0000_0000_0000_0000;
array[11406] <= 16'b0000_0000_0000_0000;
array[11407] <= 16'b0000_0000_0000_0000;
array[11408] <= 16'b0000_0000_0000_0000;
array[11409] <= 16'b0000_0000_0000_0000;
array[11410] <= 16'b0000_0000_0000_0000;
array[11411] <= 16'b0000_0000_0000_0000;
array[11412] <= 16'b0000_0000_0000_0000;
array[11413] <= 16'b0000_0000_0000_0000;
array[11414] <= 16'b0000_0000_0000_0000;
array[11415] <= 16'b0000_0000_0000_0000;
array[11416] <= 16'b0000_0000_0000_0000;
array[11417] <= 16'b0000_0000_0000_0000;
array[11418] <= 16'b0000_0000_0000_0000;
array[11419] <= 16'b0000_0000_0000_0000;
array[11420] <= 16'b0000_0000_0000_0000;
array[11421] <= 16'b0000_0000_0000_0000;
array[11422] <= 16'b0000_0000_0000_0000;
array[11423] <= 16'b0000_0000_0000_0000;
array[11424] <= 16'b0000_0000_0000_0000;
array[11425] <= 16'b0000_0000_0000_0000;
array[11426] <= 16'b0000_0000_0000_0000;
array[11427] <= 16'b0000_0000_0000_0000;
array[11428] <= 16'b0000_0000_0000_0000;
array[11429] <= 16'b0000_0000_0000_0000;
array[11430] <= 16'b0000_0000_0000_0000;
array[11431] <= 16'b0000_0000_0000_0000;
array[11432] <= 16'b0000_0000_0000_0000;
array[11433] <= 16'b0000_0000_0000_0000;
array[11434] <= 16'b0000_0000_0000_0000;
array[11435] <= 16'b0000_0000_0000_0000;
array[11436] <= 16'b0000_0000_0000_0000;
array[11437] <= 16'b0000_0000_0000_0000;
array[11438] <= 16'b0000_0000_0000_0000;
array[11439] <= 16'b0000_0000_0000_0000;
array[11440] <= 16'b0000_0000_0000_0000;
array[11441] <= 16'b0000_0000_0000_0000;
array[11442] <= 16'b0000_0000_0000_0000;
array[11443] <= 16'b0000_0000_0000_0000;
array[11444] <= 16'b0000_0000_0000_0000;
array[11445] <= 16'b0000_0000_0000_0000;
array[11446] <= 16'b0000_0000_0000_0000;
array[11447] <= 16'b0000_0000_0000_0000;
array[11448] <= 16'b0000_0000_0000_0000;
array[11449] <= 16'b0000_0000_0000_0000;
array[11450] <= 16'b0000_0000_0000_0000;
array[11451] <= 16'b0000_0000_0000_0000;
array[11452] <= 16'b0000_0000_0000_0000;
array[11453] <= 16'b0000_0000_0000_0000;
array[11454] <= 16'b0000_0000_0000_0000;
array[11455] <= 16'b0000_0000_0000_0000;
array[11456] <= 16'b0000_0000_0000_0000;
array[11457] <= 16'b0000_0000_0000_0000;
array[11458] <= 16'b0000_0000_0000_0000;
array[11459] <= 16'b0000_0000_0000_0000;
array[11460] <= 16'b0000_0000_0000_0000;
array[11461] <= 16'b0000_0000_0000_0000;
array[11462] <= 16'b0000_0000_0000_0000;
array[11463] <= 16'b0000_0000_0000_0000;
array[11464] <= 16'b0000_0000_0000_0000;
array[11465] <= 16'b0000_0000_0000_0000;
array[11466] <= 16'b0000_0000_0000_0000;
array[11467] <= 16'b0000_0000_0000_0000;
array[11468] <= 16'b0000_0000_0000_0000;
array[11469] <= 16'b0000_0000_0000_0000;
array[11470] <= 16'b0000_0000_0000_0000;
array[11471] <= 16'b0000_0000_0000_0000;
array[11472] <= 16'b0000_0000_0000_0000;
array[11473] <= 16'b0000_0000_0000_0000;
array[11474] <= 16'b0000_0000_0000_0000;
array[11475] <= 16'b0000_0000_0000_0000;
array[11476] <= 16'b0000_0000_0000_0000;
array[11477] <= 16'b0000_0000_0000_0000;
array[11478] <= 16'b0000_0000_0000_0000;
array[11479] <= 16'b0000_0000_0000_0000;
array[11480] <= 16'b0000_0000_0000_0000;
array[11481] <= 16'b0000_0000_0000_0000;
array[11482] <= 16'b0000_0000_0000_0000;
array[11483] <= 16'b0000_0000_0000_0000;
array[11484] <= 16'b0000_0000_0000_0000;
array[11485] <= 16'b0000_0000_0000_0000;
array[11486] <= 16'b0000_0000_0000_0000;
array[11487] <= 16'b0000_0000_0000_0000;
array[11488] <= 16'b0000_0000_0000_0000;
array[11489] <= 16'b0000_0000_0000_0000;
array[11490] <= 16'b0000_0000_0000_0000;
array[11491] <= 16'b0000_0000_0000_0000;
array[11492] <= 16'b0000_0000_0000_0000;
array[11493] <= 16'b0000_0000_0000_0000;
array[11494] <= 16'b0000_0000_0000_0000;
array[11495] <= 16'b0000_0000_0000_0000;
array[11496] <= 16'b0000_0000_0000_0000;
array[11497] <= 16'b0000_0000_0000_0000;
array[11498] <= 16'b0000_0000_0000_0000;
array[11499] <= 16'b0000_0000_0000_0000;
array[11500] <= 16'b0000_0000_0000_0000;
array[11501] <= 16'b0000_0000_0000_0000;
array[11502] <= 16'b0000_0000_0000_0000;
array[11503] <= 16'b0000_0000_0000_0000;
array[11504] <= 16'b0000_0000_0000_0000;
array[11505] <= 16'b0000_0000_0000_0000;
array[11506] <= 16'b0000_0000_0000_0000;
array[11507] <= 16'b0000_0000_0000_0000;
array[11508] <= 16'b0000_0000_0000_0000;
array[11509] <= 16'b0000_0000_0000_0000;
array[11510] <= 16'b0000_0000_0000_0000;
array[11511] <= 16'b0000_0000_0000_0000;
array[11512] <= 16'b0000_0000_0000_0000;
array[11513] <= 16'b0000_0000_0000_0000;
array[11514] <= 16'b0000_0000_0000_0000;
array[11515] <= 16'b0000_0000_0000_0000;
array[11516] <= 16'b0000_0000_0000_0000;
array[11517] <= 16'b0000_0000_0000_0000;
array[11518] <= 16'b0000_0000_0000_0000;
array[11519] <= 16'b0000_0000_0000_0000;
array[11520] <= 16'b0000_0000_0000_0000;
array[11521] <= 16'b0000_0000_0000_0000;
array[11522] <= 16'b0000_0000_0000_0000;
array[11523] <= 16'b0000_0000_0000_0000;
array[11524] <= 16'b0000_0000_0000_0000;
array[11525] <= 16'b0000_0000_0000_0000;
array[11526] <= 16'b0000_0000_0000_0000;
array[11527] <= 16'b0000_0000_0000_0000;
array[11528] <= 16'b0000_0000_0000_0000;
array[11529] <= 16'b0000_0000_0000_0000;
array[11530] <= 16'b0000_0000_0000_0000;
array[11531] <= 16'b0000_0000_0000_0000;
array[11532] <= 16'b0000_0000_0000_0000;
array[11533] <= 16'b0000_0000_0000_0000;
array[11534] <= 16'b0000_0000_0000_0000;
array[11535] <= 16'b0000_0000_0000_0000;
array[11536] <= 16'b0000_0000_0000_0000;
array[11537] <= 16'b0000_0000_0000_0000;
array[11538] <= 16'b0000_0000_0000_0000;
array[11539] <= 16'b0000_0000_0000_0000;
array[11540] <= 16'b0000_0000_0000_0000;
array[11541] <= 16'b0000_0000_0000_0000;
array[11542] <= 16'b0000_0000_0000_0000;
array[11543] <= 16'b0000_0000_0000_0000;
array[11544] <= 16'b0000_0000_0000_0000;
array[11545] <= 16'b0000_0000_0000_0000;
array[11546] <= 16'b0000_0000_0000_0000;
array[11547] <= 16'b0000_0000_0000_0000;
array[11548] <= 16'b0000_0000_0000_0000;
array[11549] <= 16'b0000_0000_0000_0000;
array[11550] <= 16'b0000_0000_0000_0000;
array[11551] <= 16'b0000_0000_0000_0000;
array[11552] <= 16'b0000_0000_0000_0000;
array[11553] <= 16'b0000_0000_0000_0000;
array[11554] <= 16'b0000_0000_0000_0000;
array[11555] <= 16'b0000_0000_0000_0000;
array[11556] <= 16'b0000_0000_0000_0000;
array[11557] <= 16'b0000_0000_0000_0000;
array[11558] <= 16'b0000_0000_0000_0000;
array[11559] <= 16'b0000_0000_0000_0000;
array[11560] <= 16'b0000_0000_0000_0000;
array[11561] <= 16'b0000_0000_0000_0000;
array[11562] <= 16'b0000_0000_0000_0000;
array[11563] <= 16'b0000_0000_0000_0000;
array[11564] <= 16'b0000_0000_0000_0000;
array[11565] <= 16'b0000_0000_0000_0000;
array[11566] <= 16'b0000_0000_0000_0000;
array[11567] <= 16'b0000_0000_0000_0000;
array[11568] <= 16'b0000_0000_0000_0000;
array[11569] <= 16'b0000_0000_0000_0000;
array[11570] <= 16'b0000_0000_0000_0000;
array[11571] <= 16'b0000_0000_0000_0000;
array[11572] <= 16'b0000_0000_0000_0000;
array[11573] <= 16'b0000_0000_0000_0000;
array[11574] <= 16'b0000_0000_0000_0000;
array[11575] <= 16'b0000_0000_0000_0000;
array[11576] <= 16'b0000_0000_0000_0000;
array[11577] <= 16'b0000_0000_0000_0000;
array[11578] <= 16'b0000_0000_0000_0000;
array[11579] <= 16'b0000_0000_0000_0000;
array[11580] <= 16'b0000_0000_0000_0000;
array[11581] <= 16'b0000_0000_0000_0000;
array[11582] <= 16'b0000_0000_0000_0000;
array[11583] <= 16'b0000_0000_0000_0000;
array[11584] <= 16'b0000_0000_0000_0000;
array[11585] <= 16'b0000_0000_0000_0000;
array[11586] <= 16'b0000_0000_0000_0000;
array[11587] <= 16'b0000_0000_0000_0000;
array[11588] <= 16'b0000_0000_0000_0000;
array[11589] <= 16'b0000_0000_0000_0000;
array[11590] <= 16'b0000_0000_0000_0000;
array[11591] <= 16'b0000_0000_0000_0000;
array[11592] <= 16'b0000_0000_0000_0000;
array[11593] <= 16'b0000_0000_0000_0000;
array[11594] <= 16'b0000_0000_0000_0000;
array[11595] <= 16'b0000_0000_0000_0000;
array[11596] <= 16'b0000_0000_0000_0000;
array[11597] <= 16'b0000_0000_0000_0000;
array[11598] <= 16'b0000_0000_0000_0000;
array[11599] <= 16'b0000_0000_0000_0000;
array[11600] <= 16'b0000_0000_0000_0000;
array[11601] <= 16'b0000_0000_0000_0000;
array[11602] <= 16'b0000_0000_0000_0000;
array[11603] <= 16'b0000_0000_0000_0000;
array[11604] <= 16'b0000_0000_0000_0000;
array[11605] <= 16'b0000_0000_0000_0000;
array[11606] <= 16'b0000_0000_0000_0000;
array[11607] <= 16'b0000_0000_0000_0000;
array[11608] <= 16'b0000_0000_0000_0000;
array[11609] <= 16'b0000_0000_0000_0000;
array[11610] <= 16'b0000_0000_0000_0000;
array[11611] <= 16'b0000_0000_0000_0000;
array[11612] <= 16'b0000_0000_0000_0000;
array[11613] <= 16'b0000_0000_0000_0000;
array[11614] <= 16'b0000_0000_0000_0000;
array[11615] <= 16'b0000_0000_0000_0000;
array[11616] <= 16'b0000_0000_0000_0000;
array[11617] <= 16'b0000_0000_0000_0000;
array[11618] <= 16'b0000_0000_0000_0000;
array[11619] <= 16'b0000_0000_0000_0000;
array[11620] <= 16'b0000_0000_0000_0000;
array[11621] <= 16'b0000_0000_0000_0000;
array[11622] <= 16'b0000_0000_0000_0000;
array[11623] <= 16'b0000_0000_0000_0000;
array[11624] <= 16'b0000_0000_0000_0000;
array[11625] <= 16'b0000_0000_0000_0000;
array[11626] <= 16'b0000_0000_0000_0000;
array[11627] <= 16'b0000_0000_0000_0000;
array[11628] <= 16'b0000_0000_0000_0000;
array[11629] <= 16'b0000_0000_0000_0000;
array[11630] <= 16'b0000_0000_0000_0000;
array[11631] <= 16'b0000_0000_0000_0000;
array[11632] <= 16'b0000_0000_0000_0000;
array[11633] <= 16'b0000_0000_0000_0000;
array[11634] <= 16'b0000_0000_0000_0000;
array[11635] <= 16'b0000_0000_0000_0000;
array[11636] <= 16'b0000_0000_0000_0000;
array[11637] <= 16'b0000_0000_0000_0000;
array[11638] <= 16'b0000_0000_0000_0000;
array[11639] <= 16'b0000_0000_0000_0000;
array[11640] <= 16'b0000_0000_0000_0000;
array[11641] <= 16'b0000_0000_0000_0000;
array[11642] <= 16'b0000_0000_0000_0000;
array[11643] <= 16'b0000_0000_0000_0000;
array[11644] <= 16'b0000_0000_0000_0000;
array[11645] <= 16'b0000_0000_0000_0000;
array[11646] <= 16'b0000_0000_0000_0000;
array[11647] <= 16'b0000_0000_0000_0000;
array[11648] <= 16'b0000_0000_0000_0000;
array[11649] <= 16'b0000_0000_0000_0000;
array[11650] <= 16'b0000_0000_0000_0000;
array[11651] <= 16'b0000_0000_0000_0000;
array[11652] <= 16'b0000_0000_0000_0000;
array[11653] <= 16'b0000_0000_0000_0000;
array[11654] <= 16'b0000_0000_0000_0000;
array[11655] <= 16'b0000_0000_0000_0000;
array[11656] <= 16'b0000_0000_0000_0000;
array[11657] <= 16'b0000_0000_0000_0000;
array[11658] <= 16'b0000_0000_0000_0000;
array[11659] <= 16'b0000_0000_0000_0000;
array[11660] <= 16'b0000_0000_0000_0000;
array[11661] <= 16'b0000_0000_0000_0000;
array[11662] <= 16'b0000_0000_0000_0000;
array[11663] <= 16'b0000_0000_0000_0000;
array[11664] <= 16'b0000_0000_0000_0000;
array[11665] <= 16'b0000_0000_0000_0000;
array[11666] <= 16'b0000_0000_0000_0000;
array[11667] <= 16'b0000_0000_0000_0000;
array[11668] <= 16'b0000_0000_0000_0000;
array[11669] <= 16'b0000_0000_0000_0000;
array[11670] <= 16'b0000_0000_0000_0000;
array[11671] <= 16'b0000_0000_0000_0000;
array[11672] <= 16'b0000_0000_0000_0000;
array[11673] <= 16'b0000_0000_0000_0000;
array[11674] <= 16'b0000_0000_0000_0000;
array[11675] <= 16'b0000_0000_0000_0000;
array[11676] <= 16'b0000_0000_0000_0000;
array[11677] <= 16'b0000_0000_0000_0000;
array[11678] <= 16'b0000_0000_0000_0000;
array[11679] <= 16'b0000_0000_0000_0000;
array[11680] <= 16'b0000_0000_0000_0000;
array[11681] <= 16'b0000_0000_0000_0000;
array[11682] <= 16'b0000_0000_0000_0000;
array[11683] <= 16'b0000_0000_0000_0000;
array[11684] <= 16'b0000_0000_0000_0000;
array[11685] <= 16'b0000_0000_0000_0000;
array[11686] <= 16'b0000_0000_0000_0000;
array[11687] <= 16'b0000_0000_0000_0000;
array[11688] <= 16'b0000_0000_0000_0000;
array[11689] <= 16'b0000_0000_0000_0000;
array[11690] <= 16'b0000_0000_0000_0000;
array[11691] <= 16'b0000_0000_0000_0000;
array[11692] <= 16'b0000_0000_0000_0000;
array[11693] <= 16'b0000_0000_0000_0000;
array[11694] <= 16'b0000_0000_0000_0000;
array[11695] <= 16'b0000_0000_0000_0000;
array[11696] <= 16'b0000_0000_0000_0000;
array[11697] <= 16'b0000_0000_0000_0000;
array[11698] <= 16'b0000_0000_0000_0000;
array[11699] <= 16'b0000_0000_0000_0000;
array[11700] <= 16'b0000_0000_0000_0000;
array[11701] <= 16'b0000_0000_0000_0000;
array[11702] <= 16'b0000_0000_0000_0000;
array[11703] <= 16'b0000_0000_0000_0000;
array[11704] <= 16'b0000_0000_0000_0000;
array[11705] <= 16'b0000_0000_0000_0000;
array[11706] <= 16'b0000_0000_0000_0000;
array[11707] <= 16'b0000_0000_0000_0000;
array[11708] <= 16'b0000_0000_0000_0000;
array[11709] <= 16'b0000_0000_0000_0000;
array[11710] <= 16'b0000_0000_0000_0000;
array[11711] <= 16'b0000_0000_0000_0000;
array[11712] <= 16'b0000_0000_0000_0000;
array[11713] <= 16'b0000_0000_0000_0000;
array[11714] <= 16'b0000_0000_0000_0000;
array[11715] <= 16'b0000_0000_0000_0000;
array[11716] <= 16'b0000_0000_0000_0000;
array[11717] <= 16'b0000_0000_0000_0000;
array[11718] <= 16'b0000_0000_0000_0000;
array[11719] <= 16'b0000_0000_0000_0000;
array[11720] <= 16'b0000_0000_0000_0000;
array[11721] <= 16'b0000_0000_0000_0000;
array[11722] <= 16'b0000_0000_0000_0000;
array[11723] <= 16'b0000_0000_0000_0000;
array[11724] <= 16'b0000_0000_0000_0000;
array[11725] <= 16'b0000_0000_0000_0000;
array[11726] <= 16'b0000_0000_0000_0000;
array[11727] <= 16'b0000_0000_0000_0000;
array[11728] <= 16'b0000_0000_0000_0000;
array[11729] <= 16'b0000_0000_0000_0000;
array[11730] <= 16'b0000_0000_0000_0000;
array[11731] <= 16'b0000_0000_0000_0000;
array[11732] <= 16'b0000_0000_0000_0000;
array[11733] <= 16'b0000_0000_0000_0000;
array[11734] <= 16'b0000_0000_0000_0000;
array[11735] <= 16'b0000_0000_0000_0000;
array[11736] <= 16'b0000_0000_0000_0000;
array[11737] <= 16'b0000_0000_0000_0000;
array[11738] <= 16'b0000_0000_0000_0000;
array[11739] <= 16'b0000_0000_0000_0000;
array[11740] <= 16'b0000_0000_0000_0000;
array[11741] <= 16'b0000_0000_0000_0000;
array[11742] <= 16'b0000_0000_0000_0000;
array[11743] <= 16'b0000_0000_0000_0000;
array[11744] <= 16'b0000_0000_0000_0000;
array[11745] <= 16'b0000_0000_0000_0000;
array[11746] <= 16'b0000_0000_0000_0000;
array[11747] <= 16'b0000_0000_0000_0000;
array[11748] <= 16'b0000_0000_0000_0000;
array[11749] <= 16'b0000_0000_0000_0000;
array[11750] <= 16'b0000_0000_0000_0000;
array[11751] <= 16'b0000_0000_0000_0000;
array[11752] <= 16'b0000_0000_0000_0000;
array[11753] <= 16'b0000_0000_0000_0000;
array[11754] <= 16'b0000_0000_0000_0000;
array[11755] <= 16'b0000_0000_0000_0000;
array[11756] <= 16'b0000_0000_0000_0000;
array[11757] <= 16'b0000_0000_0000_0000;
array[11758] <= 16'b0000_0000_0000_0000;
array[11759] <= 16'b0000_0000_0000_0000;
array[11760] <= 16'b0000_0000_0000_0000;
array[11761] <= 16'b0000_0000_0000_0000;
array[11762] <= 16'b0000_0000_0000_0000;
array[11763] <= 16'b0000_0000_0000_0000;
array[11764] <= 16'b0000_0000_0000_0000;
array[11765] <= 16'b0000_0000_0000_0000;
array[11766] <= 16'b0000_0000_0000_0000;
array[11767] <= 16'b0000_0000_0000_0000;
array[11768] <= 16'b0000_0000_0000_0000;
array[11769] <= 16'b0000_0000_0000_0000;
array[11770] <= 16'b0000_0000_0000_0000;
array[11771] <= 16'b0000_0000_0000_0000;
array[11772] <= 16'b0000_0000_0000_0000;
array[11773] <= 16'b0000_0000_0000_0000;
array[11774] <= 16'b0000_0000_0000_0000;
array[11775] <= 16'b0000_0000_0000_0000;
array[11776] <= 16'b0000_0000_0000_0000;
array[11777] <= 16'b0000_0000_0000_0000;
array[11778] <= 16'b0000_0000_0000_0000;
array[11779] <= 16'b0000_0000_0000_0000;
array[11780] <= 16'b0000_0000_0000_0000;
array[11781] <= 16'b0000_0000_0000_0000;
array[11782] <= 16'b0000_0000_0000_0000;
array[11783] <= 16'b0000_0000_0000_0000;
array[11784] <= 16'b0000_0000_0000_0000;
array[11785] <= 16'b0000_0000_0000_0000;
array[11786] <= 16'b0000_0000_0000_0000;
array[11787] <= 16'b0000_0000_0000_0000;
array[11788] <= 16'b0000_0000_0000_0000;
array[11789] <= 16'b0000_0000_0000_0000;
array[11790] <= 16'b0000_0000_0000_0000;
array[11791] <= 16'b0000_0000_0000_0000;
array[11792] <= 16'b0000_0000_0000_0000;
array[11793] <= 16'b0000_0000_0000_0000;
array[11794] <= 16'b0000_0000_0000_0000;
array[11795] <= 16'b0000_0000_0000_0000;
array[11796] <= 16'b0000_0000_0000_0000;
array[11797] <= 16'b0000_0000_0000_0000;
array[11798] <= 16'b0000_0000_0000_0000;
array[11799] <= 16'b0000_0000_0000_0000;
array[11800] <= 16'b0000_0000_0000_0000;
array[11801] <= 16'b0000_0000_0000_0000;
array[11802] <= 16'b0000_0000_0000_0000;
array[11803] <= 16'b0000_0000_0000_0000;
array[11804] <= 16'b0000_0000_0000_0000;
array[11805] <= 16'b0000_0000_0000_0000;
array[11806] <= 16'b0000_0000_0000_0000;
array[11807] <= 16'b0000_0000_0000_0000;
array[11808] <= 16'b0000_0000_0000_0000;
array[11809] <= 16'b0000_0000_0000_0000;
array[11810] <= 16'b0000_0000_0000_0000;
array[11811] <= 16'b0000_0000_0000_0000;
array[11812] <= 16'b0000_0000_0000_0000;
array[11813] <= 16'b0000_0000_0000_0000;
array[11814] <= 16'b0000_0000_0000_0000;
array[11815] <= 16'b0000_0000_0000_0000;
array[11816] <= 16'b0000_0000_0000_0000;
array[11817] <= 16'b0000_0000_0000_0000;
array[11818] <= 16'b0000_0000_0000_0000;
array[11819] <= 16'b0000_0000_0000_0000;
array[11820] <= 16'b0000_0000_0000_0000;
array[11821] <= 16'b0000_0000_0000_0000;
array[11822] <= 16'b0000_0000_0000_0000;
array[11823] <= 16'b0000_0000_0000_0000;
array[11824] <= 16'b0000_0000_0000_0000;
array[11825] <= 16'b0000_0000_0000_0000;
array[11826] <= 16'b0000_0000_0000_0000;
array[11827] <= 16'b0000_0000_0000_0000;
array[11828] <= 16'b0000_0000_0000_0000;
array[11829] <= 16'b0000_0000_0000_0000;
array[11830] <= 16'b0000_0000_0000_0000;
array[11831] <= 16'b0000_0000_0000_0000;
array[11832] <= 16'b0000_0000_0000_0000;
array[11833] <= 16'b0000_0000_0000_0000;
array[11834] <= 16'b0000_0000_0000_0000;
array[11835] <= 16'b0000_0000_0000_0000;
array[11836] <= 16'b0000_0000_0000_0000;
array[11837] <= 16'b0000_0000_0000_0000;
array[11838] <= 16'b0000_0000_0000_0000;
array[11839] <= 16'b0000_0000_0000_0000;
array[11840] <= 16'b0000_0000_0000_0000;
array[11841] <= 16'b0000_0000_0000_0000;
array[11842] <= 16'b0000_0000_0000_0000;
array[11843] <= 16'b0000_0000_0000_0000;
array[11844] <= 16'b0000_0000_0000_0000;
array[11845] <= 16'b0000_0000_0000_0000;
array[11846] <= 16'b0000_0000_0000_0000;
array[11847] <= 16'b0000_0000_0000_0000;
array[11848] <= 16'b0000_0000_0000_0000;
array[11849] <= 16'b0000_0000_0000_0000;
array[11850] <= 16'b0000_0000_0000_0000;
array[11851] <= 16'b0000_0000_0000_0000;
array[11852] <= 16'b0000_0000_0000_0000;
array[11853] <= 16'b0000_0000_0000_0000;
array[11854] <= 16'b0000_0000_0000_0000;
array[11855] <= 16'b0000_0000_0000_0000;
array[11856] <= 16'b0000_0000_0000_0000;
array[11857] <= 16'b0000_0000_0000_0000;
array[11858] <= 16'b0000_0000_0000_0000;
array[11859] <= 16'b0000_0000_0000_0000;
array[11860] <= 16'b0000_0000_0000_0000;
array[11861] <= 16'b0000_0000_0000_0000;
array[11862] <= 16'b0000_0000_0000_0000;
array[11863] <= 16'b0000_0000_0000_0000;
array[11864] <= 16'b0000_0000_0000_0000;
array[11865] <= 16'b0000_0000_0000_0000;
array[11866] <= 16'b0000_0000_0000_0000;
array[11867] <= 16'b0000_0000_0000_0000;
array[11868] <= 16'b0000_0000_0000_0000;
array[11869] <= 16'b0000_0000_0000_0000;
array[11870] <= 16'b0000_0000_0000_0000;
array[11871] <= 16'b0000_0000_0000_0000;
array[11872] <= 16'b0000_0000_0000_0000;
array[11873] <= 16'b0000_0000_0000_0000;
array[11874] <= 16'b0000_0000_0000_0000;
array[11875] <= 16'b0000_0000_0000_0000;
array[11876] <= 16'b0000_0000_0000_0000;
array[11877] <= 16'b0000_0000_0000_0000;
array[11878] <= 16'b0000_0000_0000_0000;
array[11879] <= 16'b0000_0000_0000_0000;
array[11880] <= 16'b0000_0000_0000_0000;
array[11881] <= 16'b0000_0000_0000_0000;
array[11882] <= 16'b0000_0000_0000_0000;
array[11883] <= 16'b0000_0000_0000_0000;
array[11884] <= 16'b0000_0000_0000_0000;
array[11885] <= 16'b0000_0000_0000_0000;
array[11886] <= 16'b0000_0000_0000_0000;
array[11887] <= 16'b0000_0000_0000_0000;
array[11888] <= 16'b0000_0000_0000_0000;
array[11889] <= 16'b0000_0000_0000_0000;
array[11890] <= 16'b0000_0000_0000_0000;
array[11891] <= 16'b0000_0000_0000_0000;
array[11892] <= 16'b0000_0000_0000_0000;
array[11893] <= 16'b0000_0000_0000_0000;
array[11894] <= 16'b0000_0000_0000_0000;
array[11895] <= 16'b0000_0000_0000_0000;
array[11896] <= 16'b0000_0000_0000_0000;
array[11897] <= 16'b0000_0000_0000_0000;
array[11898] <= 16'b0000_0000_0000_0000;
array[11899] <= 16'b0000_0000_0000_0000;
array[11900] <= 16'b0000_0000_0000_0000;
array[11901] <= 16'b0000_0000_0000_0000;
array[11902] <= 16'b0000_0000_0000_0000;
array[11903] <= 16'b0000_0000_0000_0000;
array[11904] <= 16'b0000_0000_0000_0000;
array[11905] <= 16'b0000_0000_0000_0000;
array[11906] <= 16'b0000_0000_0000_0000;
array[11907] <= 16'b0000_0000_0000_0000;
array[11908] <= 16'b0000_0000_0000_0000;
array[11909] <= 16'b0000_0000_0000_0000;
array[11910] <= 16'b0000_0000_0000_0000;
array[11911] <= 16'b0000_0000_0000_0000;
array[11912] <= 16'b0000_0000_0000_0000;
array[11913] <= 16'b0000_0000_0000_0000;
array[11914] <= 16'b0000_0000_0000_0000;
array[11915] <= 16'b0000_0000_0000_0000;
array[11916] <= 16'b0000_0000_0000_0000;
array[11917] <= 16'b0000_0000_0000_0000;
array[11918] <= 16'b0000_0000_0000_0000;
array[11919] <= 16'b0000_0000_0000_0000;
array[11920] <= 16'b0000_0000_0000_0000;
array[11921] <= 16'b0000_0000_0000_0000;
array[11922] <= 16'b0000_0000_0000_0000;
array[11923] <= 16'b0000_0000_0000_0000;
array[11924] <= 16'b0000_0000_0000_0000;
array[11925] <= 16'b0000_0000_0000_0000;
array[11926] <= 16'b0000_0000_0000_0000;
array[11927] <= 16'b0000_0000_0000_0000;
array[11928] <= 16'b0000_0000_0000_0000;
array[11929] <= 16'b0000_0000_0000_0000;
array[11930] <= 16'b0000_0000_0000_0000;
array[11931] <= 16'b0000_0000_0000_0000;
array[11932] <= 16'b0000_0000_0000_0000;
array[11933] <= 16'b0000_0000_0000_0000;
array[11934] <= 16'b0000_0000_0000_0000;
array[11935] <= 16'b0000_0000_0000_0000;
array[11936] <= 16'b0000_0000_0000_0000;
array[11937] <= 16'b0000_0000_0000_0000;
array[11938] <= 16'b0000_0000_0000_0000;
array[11939] <= 16'b0000_0000_0000_0000;
array[11940] <= 16'b0000_0000_0000_0000;
array[11941] <= 16'b0000_0000_0000_0000;
array[11942] <= 16'b0000_0000_0000_0000;
array[11943] <= 16'b0000_0000_0000_0000;
array[11944] <= 16'b0000_0000_0000_0000;
array[11945] <= 16'b0000_0000_0000_0000;
array[11946] <= 16'b0000_0000_0000_0000;
array[11947] <= 16'b0000_0000_0000_0000;
array[11948] <= 16'b0000_0000_0000_0000;
array[11949] <= 16'b0000_0000_0000_0000;
array[11950] <= 16'b0000_0000_0000_0000;
array[11951] <= 16'b0000_0000_0000_0000;
array[11952] <= 16'b0000_0000_0000_0000;
array[11953] <= 16'b0000_0000_0000_0000;
array[11954] <= 16'b0000_0000_0000_0000;
array[11955] <= 16'b0000_0000_0000_0000;
array[11956] <= 16'b0000_0000_0000_0000;
array[11957] <= 16'b0000_0000_0000_0000;
array[11958] <= 16'b0000_0000_0000_0000;
array[11959] <= 16'b0000_0000_0000_0000;
array[11960] <= 16'b0000_0000_0000_0000;
array[11961] <= 16'b0000_0000_0000_0000;
array[11962] <= 16'b0000_0000_0000_0000;
array[11963] <= 16'b0000_0000_0000_0000;
array[11964] <= 16'b0000_0000_0000_0000;
array[11965] <= 16'b0000_0000_0000_0000;
array[11966] <= 16'b0000_0000_0000_0000;
array[11967] <= 16'b0000_0000_0000_0000;
array[11968] <= 16'b0000_0000_0000_0000;
array[11969] <= 16'b0000_0000_0000_0000;
array[11970] <= 16'b0000_0000_0000_0000;
array[11971] <= 16'b0000_0000_0000_0000;
array[11972] <= 16'b0000_0000_0000_0000;
array[11973] <= 16'b0000_0000_0000_0000;
array[11974] <= 16'b0000_0000_0000_0000;
array[11975] <= 16'b0000_0000_0000_0000;
array[11976] <= 16'b0000_0000_0000_0000;
array[11977] <= 16'b0000_0000_0000_0000;
array[11978] <= 16'b0000_0000_0000_0000;
array[11979] <= 16'b0000_0000_0000_0000;
array[11980] <= 16'b0000_0000_0000_0000;
array[11981] <= 16'b0000_0000_0000_0000;
array[11982] <= 16'b0000_0000_0000_0000;
array[11983] <= 16'b0000_0000_0000_0000;
array[11984] <= 16'b0000_0000_0000_0000;
array[11985] <= 16'b0000_0000_0000_0000;
array[11986] <= 16'b0000_0000_0000_0000;
array[11987] <= 16'b0000_0000_0000_0000;
array[11988] <= 16'b0000_0000_0000_0000;
array[11989] <= 16'b0000_0000_0000_0000;
array[11990] <= 16'b0000_0000_0000_0000;
array[11991] <= 16'b0000_0000_0000_0000;
array[11992] <= 16'b0000_0000_0000_0000;
array[11993] <= 16'b0000_0000_0000_0000;
array[11994] <= 16'b0000_0000_0000_0000;
array[11995] <= 16'b0000_0000_0000_0000;
array[11996] <= 16'b0000_0000_0000_0000;
array[11997] <= 16'b0000_0000_0000_0000;
array[11998] <= 16'b0000_0000_0000_0000;
array[11999] <= 16'b0000_0000_0000_0000;
array[12000] <= 16'b0000_0000_0000_0000;
array[12001] <= 16'b0000_0000_0000_0000;
array[12002] <= 16'b0000_0000_0000_0000;
array[12003] <= 16'b0000_0000_0000_0000;
array[12004] <= 16'b0000_0000_0000_0000;
array[12005] <= 16'b0000_0000_0000_0000;
array[12006] <= 16'b0000_0000_0000_0000;
array[12007] <= 16'b0000_0000_0000_0000;
array[12008] <= 16'b0000_0000_0000_0000;
array[12009] <= 16'b0000_0000_0000_0000;
array[12010] <= 16'b0000_0000_0000_0000;
array[12011] <= 16'b0000_0000_0000_0000;
array[12012] <= 16'b0000_0000_0000_0000;
array[12013] <= 16'b0000_0000_0000_0000;
array[12014] <= 16'b0000_0000_0000_0000;
array[12015] <= 16'b0000_0000_0000_0000;
array[12016] <= 16'b0000_0000_0000_0000;
array[12017] <= 16'b0000_0000_0000_0000;
array[12018] <= 16'b0000_0000_0000_0000;
array[12019] <= 16'b0000_0000_0000_0000;
array[12020] <= 16'b0000_0000_0000_0000;
array[12021] <= 16'b0000_0000_0000_0000;
array[12022] <= 16'b0000_0000_0000_0000;
array[12023] <= 16'b0000_0000_0000_0000;
array[12024] <= 16'b0000_0000_0000_0000;
array[12025] <= 16'b0000_0000_0000_0000;
array[12026] <= 16'b0000_0000_0000_0000;
array[12027] <= 16'b0000_0000_0000_0000;
array[12028] <= 16'b0000_0000_0000_0000;
array[12029] <= 16'b0000_0000_0000_0000;
array[12030] <= 16'b0000_0000_0000_0000;
array[12031] <= 16'b0000_0000_0000_0000;
array[12032] <= 16'b0000_0000_0000_0000;
array[12033] <= 16'b0000_0000_0000_0000;
array[12034] <= 16'b0000_0000_0000_0000;
array[12035] <= 16'b0000_0000_0000_0000;
array[12036] <= 16'b0000_0000_0000_0000;
array[12037] <= 16'b0000_0000_0000_0000;
array[12038] <= 16'b0000_0000_0000_0000;
array[12039] <= 16'b0000_0000_0000_0000;
array[12040] <= 16'b0000_0000_0000_0000;
array[12041] <= 16'b0000_0000_0000_0000;
array[12042] <= 16'b0000_0000_0000_0000;
array[12043] <= 16'b0000_0000_0000_0000;
array[12044] <= 16'b0000_0000_0000_0000;
array[12045] <= 16'b0000_0000_0000_0000;
array[12046] <= 16'b0000_0000_0000_0000;
array[12047] <= 16'b0000_0000_0000_0000;
array[12048] <= 16'b0000_0000_0000_0000;
array[12049] <= 16'b0000_0000_0000_0000;
array[12050] <= 16'b0000_0000_0000_0000;
array[12051] <= 16'b0000_0000_0000_0000;
array[12052] <= 16'b0000_0000_0000_0000;
array[12053] <= 16'b0000_0000_0000_0000;
array[12054] <= 16'b0000_0000_0000_0000;
array[12055] <= 16'b0000_0000_0000_0000;
array[12056] <= 16'b0000_0000_0000_0000;
array[12057] <= 16'b0000_0000_0000_0000;
array[12058] <= 16'b0000_0000_0000_0000;
array[12059] <= 16'b0000_0000_0000_0000;
array[12060] <= 16'b0000_0000_0000_0000;
array[12061] <= 16'b0000_0000_0000_0000;
array[12062] <= 16'b0000_0000_0000_0000;
array[12063] <= 16'b0000_0000_0000_0000;
array[12064] <= 16'b0000_0000_0000_0000;
array[12065] <= 16'b0000_0000_0000_0000;
array[12066] <= 16'b0000_0000_0000_0000;
array[12067] <= 16'b0000_0000_0000_0000;
array[12068] <= 16'b0000_0000_0000_0000;
array[12069] <= 16'b0000_0000_0000_0000;
array[12070] <= 16'b0000_0000_0000_0000;
array[12071] <= 16'b0000_0000_0000_0000;
array[12072] <= 16'b0000_0000_0000_0000;
array[12073] <= 16'b0000_0000_0000_0000;
array[12074] <= 16'b0000_0000_0000_0000;
array[12075] <= 16'b0000_0000_0000_0000;
array[12076] <= 16'b0000_0000_0000_0000;
array[12077] <= 16'b0000_0000_0000_0000;
array[12078] <= 16'b0000_0000_0000_0000;
array[12079] <= 16'b0000_0000_0000_0000;
array[12080] <= 16'b0000_0000_0000_0000;
array[12081] <= 16'b0000_0000_0000_0000;
array[12082] <= 16'b0000_0000_0000_0000;
array[12083] <= 16'b0000_0000_0000_0000;
array[12084] <= 16'b0000_0000_0000_0000;
array[12085] <= 16'b0000_0000_0000_0000;
array[12086] <= 16'b0000_0000_0000_0000;
array[12087] <= 16'b0000_0000_0000_0000;
array[12088] <= 16'b0000_0000_0000_0000;
array[12089] <= 16'b0000_0000_0000_0000;
array[12090] <= 16'b0000_0000_0000_0000;
array[12091] <= 16'b0000_0000_0000_0000;
array[12092] <= 16'b0000_0000_0000_0000;
array[12093] <= 16'b0000_0000_0000_0000;
array[12094] <= 16'b0000_0000_0000_0000;
array[12095] <= 16'b0000_0000_0000_0000;
array[12096] <= 16'b0000_0000_0000_0000;
array[12097] <= 16'b0000_0000_0000_0000;
array[12098] <= 16'b0000_0000_0000_0000;
array[12099] <= 16'b0000_0000_0000_0000;
array[12100] <= 16'b0000_0000_0000_0000;
array[12101] <= 16'b0000_0000_0000_0000;
array[12102] <= 16'b0000_0000_0000_0000;
array[12103] <= 16'b0000_0000_0000_0000;
array[12104] <= 16'b0000_0000_0000_0000;
array[12105] <= 16'b0000_0000_0000_0000;
array[12106] <= 16'b0000_0000_0000_0000;
array[12107] <= 16'b0000_0000_0000_0000;
array[12108] <= 16'b0000_0000_0000_0000;
array[12109] <= 16'b0000_0000_0000_0000;
array[12110] <= 16'b0000_0000_0000_0000;
array[12111] <= 16'b0000_0000_0000_0000;
array[12112] <= 16'b0000_0000_0000_0000;
array[12113] <= 16'b0000_0000_0000_0000;
array[12114] <= 16'b0000_0000_0000_0000;
array[12115] <= 16'b0000_0000_0000_0000;
array[12116] <= 16'b0000_0000_0000_0000;
array[12117] <= 16'b0000_0000_0000_0000;
array[12118] <= 16'b0000_0000_0000_0000;
array[12119] <= 16'b0000_0000_0000_0000;
array[12120] <= 16'b0000_0000_0000_0000;
array[12121] <= 16'b0000_0000_0000_0000;
array[12122] <= 16'b0000_0000_0000_0000;
array[12123] <= 16'b0000_0000_0000_0000;
array[12124] <= 16'b0000_0000_0000_0000;
array[12125] <= 16'b0000_0000_0000_0000;
array[12126] <= 16'b0000_0000_0000_0000;
array[12127] <= 16'b0000_0000_0000_0000;
array[12128] <= 16'b0000_0000_0000_0000;
array[12129] <= 16'b0000_0000_0000_0000;
array[12130] <= 16'b0000_0000_0000_0000;
array[12131] <= 16'b0000_0000_0000_0000;
array[12132] <= 16'b0000_0000_0000_0000;
array[12133] <= 16'b0000_0000_0000_0000;
array[12134] <= 16'b0000_0000_0000_0000;
array[12135] <= 16'b0000_0000_0000_0000;
array[12136] <= 16'b0000_0000_0000_0000;
array[12137] <= 16'b0000_0000_0000_0000;
array[12138] <= 16'b0000_0000_0000_0000;
array[12139] <= 16'b0000_0000_0000_0000;
array[12140] <= 16'b0000_0000_0000_0000;
array[12141] <= 16'b0000_0000_0000_0000;
array[12142] <= 16'b0000_0000_0000_0000;
array[12143] <= 16'b0000_0000_0000_0000;
array[12144] <= 16'b0000_0000_0000_0000;
array[12145] <= 16'b0000_0000_0000_0000;
array[12146] <= 16'b0000_0000_0000_0000;
array[12147] <= 16'b0000_0000_0000_0000;
array[12148] <= 16'b0000_0000_0000_0000;
array[12149] <= 16'b0000_0000_0000_0000;
array[12150] <= 16'b0000_0000_0000_0000;
array[12151] <= 16'b0000_0000_0000_0000;
array[12152] <= 16'b0000_0000_0000_0000;
array[12153] <= 16'b0000_0000_0000_0000;
array[12154] <= 16'b0000_0000_0000_0000;
array[12155] <= 16'b0000_0000_0000_0000;
array[12156] <= 16'b0000_0000_0000_0000;
array[12157] <= 16'b0000_0000_0000_0000;
array[12158] <= 16'b0000_0000_0000_0000;
array[12159] <= 16'b0000_0000_0000_0000;
array[12160] <= 16'b0000_0000_0000_0000;
array[12161] <= 16'b0000_0000_0000_0000;
array[12162] <= 16'b0000_0000_0000_0000;
array[12163] <= 16'b0000_0000_0000_0000;
array[12164] <= 16'b0000_0000_0000_0000;
array[12165] <= 16'b0000_0000_0000_0000;
array[12166] <= 16'b0000_0000_0000_0000;
array[12167] <= 16'b0000_0000_0000_0000;
array[12168] <= 16'b0000_0000_0000_0000;
array[12169] <= 16'b0000_0000_0000_0000;
array[12170] <= 16'b0000_0000_0000_0000;
array[12171] <= 16'b0000_0000_0000_0000;
array[12172] <= 16'b0000_0000_0000_0000;
array[12173] <= 16'b0000_0000_0000_0000;
array[12174] <= 16'b0000_0000_0000_0000;
array[12175] <= 16'b0000_0000_0000_0000;
array[12176] <= 16'b0000_0000_0000_0000;
array[12177] <= 16'b0000_0000_0000_0000;
array[12178] <= 16'b0000_0000_0000_0000;
array[12179] <= 16'b0000_0000_0000_0000;
array[12180] <= 16'b0000_0000_0000_0000;
array[12181] <= 16'b0000_0000_0000_0000;
array[12182] <= 16'b0000_0000_0000_0000;
array[12183] <= 16'b0000_0000_0000_0000;
array[12184] <= 16'b0000_0000_0000_0000;
array[12185] <= 16'b0000_0000_0000_0000;
array[12186] <= 16'b0000_0000_0000_0000;
array[12187] <= 16'b0000_0000_0000_0000;
array[12188] <= 16'b0000_0000_0000_0000;
array[12189] <= 16'b0000_0000_0000_0000;
array[12190] <= 16'b0000_0000_0000_0000;
array[12191] <= 16'b0000_0000_0000_0000;
array[12192] <= 16'b0000_0000_0000_0000;
array[12193] <= 16'b0000_0000_0000_0000;
array[12194] <= 16'b0000_0000_0000_0000;
array[12195] <= 16'b0000_0000_0000_0000;
array[12196] <= 16'b0000_0000_0000_0000;
array[12197] <= 16'b0000_0000_0000_0000;
array[12198] <= 16'b0000_0000_0000_0000;
array[12199] <= 16'b0000_0000_0000_0000;
array[12200] <= 16'b0000_0000_0000_0000;
array[12201] <= 16'b0000_0000_0000_0000;
array[12202] <= 16'b0000_0000_0000_0000;
array[12203] <= 16'b0000_0000_0000_0000;
array[12204] <= 16'b0000_0000_0000_0000;
array[12205] <= 16'b0000_0000_0000_0000;
array[12206] <= 16'b0000_0000_0000_0000;
array[12207] <= 16'b0000_0000_0000_0000;
array[12208] <= 16'b0000_0000_0000_0000;
array[12209] <= 16'b0000_0000_0000_0000;
array[12210] <= 16'b0000_0000_0000_0000;
array[12211] <= 16'b0000_0000_0000_0000;
array[12212] <= 16'b0000_0000_0000_0000;
array[12213] <= 16'b0000_0000_0000_0000;
array[12214] <= 16'b0000_0000_0000_0000;
array[12215] <= 16'b0000_0000_0000_0000;
array[12216] <= 16'b0000_0000_0000_0000;
array[12217] <= 16'b0000_0000_0000_0000;
array[12218] <= 16'b0000_0000_0000_0000;
array[12219] <= 16'b0000_0000_0000_0000;
array[12220] <= 16'b0000_0000_0000_0000;
array[12221] <= 16'b0000_0000_0000_0000;
array[12222] <= 16'b0000_0000_0000_0000;
array[12223] <= 16'b0000_0000_0000_0000;
array[12224] <= 16'b0000_0000_0000_0000;
array[12225] <= 16'b0000_0000_0000_0000;
array[12226] <= 16'b0000_0000_0000_0000;
array[12227] <= 16'b0000_0000_0000_0000;
array[12228] <= 16'b0000_0000_0000_0000;
array[12229] <= 16'b0000_0000_0000_0000;
array[12230] <= 16'b0000_0000_0000_0000;
array[12231] <= 16'b0000_0000_0000_0000;
array[12232] <= 16'b0000_0000_0000_0000;
array[12233] <= 16'b0000_0000_0000_0000;
array[12234] <= 16'b0000_0000_0000_0000;
array[12235] <= 16'b0000_0000_0000_0000;
array[12236] <= 16'b0000_0000_0000_0000;
array[12237] <= 16'b0000_0000_0000_0000;
array[12238] <= 16'b0000_0000_0000_0000;
array[12239] <= 16'b0000_0000_0000_0000;
array[12240] <= 16'b0000_0000_0000_0000;
array[12241] <= 16'b0000_0000_0000_0000;
array[12242] <= 16'b0000_0000_0000_0000;
array[12243] <= 16'b0000_0000_0000_0000;
array[12244] <= 16'b0000_0000_0000_0000;
array[12245] <= 16'b0000_0000_0000_0000;
array[12246] <= 16'b0000_0000_0000_0000;
array[12247] <= 16'b0000_0000_0000_0000;
array[12248] <= 16'b0000_0000_0000_0000;
array[12249] <= 16'b0000_0000_0000_0000;
array[12250] <= 16'b0000_0000_0000_0000;
array[12251] <= 16'b0000_0000_0000_0000;
array[12252] <= 16'b0000_0000_0000_0000;
array[12253] <= 16'b0000_0000_0000_0000;
array[12254] <= 16'b0000_0000_0000_0000;
array[12255] <= 16'b0000_0000_0000_0000;
array[12256] <= 16'b0000_0000_0000_0000;
array[12257] <= 16'b0000_0000_0000_0000;
array[12258] <= 16'b0000_0000_0000_0000;
array[12259] <= 16'b0000_0000_0000_0000;
array[12260] <= 16'b0000_0000_0000_0000;
array[12261] <= 16'b0000_0000_0000_0000;
array[12262] <= 16'b0000_0000_0000_0000;
array[12263] <= 16'b0000_0000_0000_0000;
array[12264] <= 16'b0000_0000_0000_0000;
array[12265] <= 16'b0000_0000_0000_0000;
array[12266] <= 16'b0000_0000_0000_0000;
array[12267] <= 16'b0000_0000_0000_0000;
array[12268] <= 16'b0000_0000_0000_0000;
array[12269] <= 16'b0000_0000_0000_0000;
array[12270] <= 16'b0000_0000_0000_0000;
array[12271] <= 16'b0000_0000_0000_0000;
array[12272] <= 16'b0000_0000_0000_0000;
array[12273] <= 16'b0000_0000_0000_0000;
array[12274] <= 16'b0000_0000_0000_0000;
array[12275] <= 16'b0000_0000_0000_0000;
array[12276] <= 16'b0000_0000_0000_0000;
array[12277] <= 16'b0000_0000_0000_0000;
array[12278] <= 16'b0000_0000_0000_0000;
array[12279] <= 16'b0000_0000_0000_0000;
array[12280] <= 16'b0000_0000_0000_0000;
array[12281] <= 16'b0000_0000_0000_0000;
array[12282] <= 16'b0000_0000_0000_0000;
array[12283] <= 16'b0000_0000_0000_0000;
array[12284] <= 16'b0000_0000_0000_0000;
array[12285] <= 16'b0000_0000_0000_0000;
array[12286] <= 16'b0000_0000_0000_0000;
array[12287] <= 16'b0000_0000_0000_0000;
array[12288] <= 16'b0000_0000_0000_0000;
array[12289] <= 16'b0000_0000_0000_0000;
array[12290] <= 16'b0000_0000_0000_0000;
array[12291] <= 16'b0000_0000_0000_0000;
array[12292] <= 16'b0000_0000_0000_0000;
array[12293] <= 16'b0000_0000_0000_0000;
array[12294] <= 16'b0000_0000_0000_0000;
array[12295] <= 16'b0000_0000_0000_0000;
array[12296] <= 16'b0000_0000_0000_0000;
array[12297] <= 16'b0000_0000_0000_0000;
array[12298] <= 16'b0000_0000_0000_0000;
array[12299] <= 16'b0000_0000_0000_0000;
array[12300] <= 16'b0000_0000_0000_0000;
array[12301] <= 16'b0000_0000_0000_0000;
array[12302] <= 16'b0000_0000_0000_0000;
array[12303] <= 16'b0000_0000_0000_0000;
array[12304] <= 16'b0000_0000_0000_0000;
array[12305] <= 16'b0000_0000_0000_0000;
array[12306] <= 16'b0000_0000_0000_0000;
array[12307] <= 16'b0000_0000_0000_0000;
array[12308] <= 16'b0000_0000_0000_0000;
array[12309] <= 16'b0000_0000_0000_0000;
array[12310] <= 16'b0000_0000_0000_0000;
array[12311] <= 16'b0000_0000_0000_0000;
array[12312] <= 16'b0000_0000_0000_0000;
array[12313] <= 16'b0000_0000_0000_0000;
array[12314] <= 16'b0000_0000_0000_0000;
array[12315] <= 16'b0000_0000_0000_0000;
array[12316] <= 16'b0000_0000_0000_0000;
array[12317] <= 16'b0000_0000_0000_0000;
array[12318] <= 16'b0000_0000_0000_0000;
array[12319] <= 16'b0000_0000_0000_0000;
array[12320] <= 16'b0000_0000_0000_0000;
array[12321] <= 16'b0000_0000_0000_0000;
array[12322] <= 16'b0000_0000_0000_0000;
array[12323] <= 16'b0000_0000_0000_0000;
array[12324] <= 16'b0000_0000_0000_0000;
array[12325] <= 16'b0000_0000_0000_0000;
array[12326] <= 16'b0000_0000_0000_0000;
array[12327] <= 16'b0000_0000_0000_0000;
array[12328] <= 16'b0000_0000_0000_0000;
array[12329] <= 16'b0000_0000_0000_0000;
array[12330] <= 16'b0000_0000_0000_0000;
array[12331] <= 16'b0000_0000_0000_0000;
array[12332] <= 16'b0000_0000_0000_0000;
array[12333] <= 16'b0000_0000_0000_0000;
array[12334] <= 16'b0000_0000_0000_0000;
array[12335] <= 16'b0000_0000_0000_0000;
array[12336] <= 16'b0000_0000_0000_0000;
array[12337] <= 16'b0000_0000_0000_0000;
array[12338] <= 16'b0000_0000_0000_0000;
array[12339] <= 16'b0000_0000_0000_0000;
array[12340] <= 16'b0000_0000_0000_0000;
array[12341] <= 16'b0000_0000_0000_0000;
array[12342] <= 16'b0000_0000_0000_0000;
array[12343] <= 16'b0000_0000_0000_0000;
array[12344] <= 16'b0000_0000_0000_0000;
array[12345] <= 16'b0000_0000_0000_0000;
array[12346] <= 16'b0000_0000_0000_0000;
array[12347] <= 16'b0000_0000_0000_0000;
array[12348] <= 16'b0000_0000_0000_0000;
array[12349] <= 16'b0000_0000_0000_0000;
array[12350] <= 16'b0000_0000_0000_0000;
array[12351] <= 16'b0000_0000_0000_0000;
array[12352] <= 16'b0000_0000_0000_0000;
array[12353] <= 16'b0000_0000_0000_0000;
array[12354] <= 16'b0000_0000_0000_0000;
array[12355] <= 16'b0000_0000_0000_0000;
array[12356] <= 16'b0000_0000_0000_0000;
array[12357] <= 16'b0000_0000_0000_0000;
array[12358] <= 16'b0000_0000_0000_0000;
array[12359] <= 16'b0000_0000_0000_0000;
array[12360] <= 16'b0000_0000_0000_0000;
array[12361] <= 16'b0000_0000_0000_0000;
array[12362] <= 16'b0000_0000_0000_0000;
array[12363] <= 16'b0000_0000_0000_0000;
array[12364] <= 16'b0000_0000_0000_0000;
array[12365] <= 16'b0000_0000_0000_0000;
array[12366] <= 16'b0000_0000_0000_0000;
array[12367] <= 16'b0000_0000_0000_0000;
array[12368] <= 16'b0000_0000_0000_0000;
array[12369] <= 16'b0000_0000_0000_0000;
array[12370] <= 16'b0000_0000_0000_0000;
array[12371] <= 16'b0000_0000_0000_0000;
array[12372] <= 16'b0000_0000_0000_0000;
array[12373] <= 16'b0000_0000_0000_0000;
array[12374] <= 16'b0000_0000_0000_0000;
array[12375] <= 16'b0000_0000_0000_0000;
array[12376] <= 16'b0000_0000_0000_0000;
array[12377] <= 16'b0000_0000_0000_0000;
array[12378] <= 16'b0000_0000_0000_0000;
array[12379] <= 16'b0000_0000_0000_0000;
array[12380] <= 16'b0000_0000_0000_0000;
array[12381] <= 16'b0000_0000_0000_0000;
array[12382] <= 16'b0000_0000_0000_0000;
array[12383] <= 16'b0000_0000_0000_0000;
array[12384] <= 16'b0000_0000_0000_0000;
array[12385] <= 16'b0000_0000_0000_0000;
array[12386] <= 16'b0000_0000_0000_0000;
array[12387] <= 16'b0000_0000_0000_0000;
array[12388] <= 16'b0000_0000_0000_0000;
array[12389] <= 16'b0000_0000_0000_0000;
array[12390] <= 16'b0000_0000_0000_0000;
array[12391] <= 16'b0000_0000_0000_0000;
array[12392] <= 16'b0000_0000_0000_0000;
array[12393] <= 16'b0000_0000_0000_0000;
array[12394] <= 16'b0000_0000_0000_0000;
array[12395] <= 16'b0000_0000_0000_0000;
array[12396] <= 16'b0000_0000_0000_0000;
array[12397] <= 16'b0000_0000_0000_0000;
array[12398] <= 16'b0000_0000_0000_0000;
array[12399] <= 16'b0000_0000_0000_0000;
array[12400] <= 16'b0000_0000_0000_0000;
array[12401] <= 16'b0000_0000_0000_0000;
array[12402] <= 16'b0000_0000_0000_0000;
array[12403] <= 16'b0000_0000_0000_0000;
array[12404] <= 16'b0000_0000_0000_0000;
array[12405] <= 16'b0000_0000_0000_0000;
array[12406] <= 16'b0000_0000_0000_0000;
array[12407] <= 16'b0000_0000_0000_0000;
array[12408] <= 16'b0000_0000_0000_0000;
array[12409] <= 16'b0000_0000_0000_0000;
array[12410] <= 16'b0000_0000_0000_0000;
array[12411] <= 16'b0000_0000_0000_0000;
array[12412] <= 16'b0000_0000_0000_0000;
array[12413] <= 16'b0000_0000_0000_0000;
array[12414] <= 16'b0000_0000_0000_0000;
array[12415] <= 16'b0000_0000_0000_0000;
array[12416] <= 16'b0000_0000_0000_0000;
array[12417] <= 16'b0000_0000_0000_0000;
array[12418] <= 16'b0000_0000_0000_0000;
array[12419] <= 16'b0000_0000_0000_0000;
array[12420] <= 16'b0000_0000_0000_0000;
array[12421] <= 16'b0000_0000_0000_0000;
array[12422] <= 16'b0000_0000_0000_0000;
array[12423] <= 16'b0000_0000_0000_0000;
array[12424] <= 16'b0000_0000_0000_0000;
array[12425] <= 16'b0000_0000_0000_0000;
array[12426] <= 16'b0000_0000_0000_0000;
array[12427] <= 16'b0000_0000_0000_0000;
array[12428] <= 16'b0000_0000_0000_0000;
array[12429] <= 16'b0000_0000_0000_0000;
array[12430] <= 16'b0000_0000_0000_0000;
array[12431] <= 16'b0000_0000_0000_0000;
array[12432] <= 16'b0000_0000_0000_0000;
array[12433] <= 16'b0000_0000_0000_0000;
array[12434] <= 16'b0000_0000_0000_0000;
array[12435] <= 16'b0000_0000_0000_0000;
array[12436] <= 16'b0000_0000_0000_0000;
array[12437] <= 16'b0000_0000_0000_0000;
array[12438] <= 16'b0000_0000_0000_0000;
array[12439] <= 16'b0000_0000_0000_0000;
array[12440] <= 16'b0000_0000_0000_0000;
array[12441] <= 16'b0000_0000_0000_0000;
array[12442] <= 16'b0000_0000_0000_0000;
array[12443] <= 16'b0000_0000_0000_0000;
array[12444] <= 16'b0000_0000_0000_0000;
array[12445] <= 16'b0000_0000_0000_0000;
array[12446] <= 16'b0000_0000_0000_0000;
array[12447] <= 16'b0000_0000_0000_0000;
array[12448] <= 16'b0000_0000_0000_0000;
array[12449] <= 16'b0000_0000_0000_0000;
array[12450] <= 16'b0000_0000_0000_0000;
array[12451] <= 16'b0000_0000_0000_0000;
array[12452] <= 16'b0000_0000_0000_0000;
array[12453] <= 16'b0000_0000_0000_0000;
array[12454] <= 16'b0000_0000_0000_0000;
array[12455] <= 16'b0000_0000_0000_0000;
array[12456] <= 16'b0000_0000_0000_0000;
array[12457] <= 16'b0000_0000_0000_0000;
array[12458] <= 16'b0000_0000_0000_0000;
array[12459] <= 16'b0000_0000_0000_0000;
array[12460] <= 16'b0000_0000_0000_0000;
array[12461] <= 16'b0000_0000_0000_0000;
array[12462] <= 16'b0000_0000_0000_0000;
array[12463] <= 16'b0000_0000_0000_0000;
array[12464] <= 16'b0000_0000_0000_0000;
array[12465] <= 16'b0000_0000_0000_0000;
array[12466] <= 16'b0000_0000_0000_0000;
array[12467] <= 16'b0000_0000_0000_0000;
array[12468] <= 16'b0000_0000_0000_0000;
array[12469] <= 16'b0000_0000_0000_0000;
array[12470] <= 16'b0000_0000_0000_0000;
array[12471] <= 16'b0000_0000_0000_0000;
array[12472] <= 16'b0000_0000_0000_0000;
array[12473] <= 16'b0000_0000_0000_0000;
array[12474] <= 16'b0000_0000_0000_0000;
array[12475] <= 16'b0000_0000_0000_0000;
array[12476] <= 16'b0000_0000_0000_0000;
array[12477] <= 16'b0000_0000_0000_0000;
array[12478] <= 16'b0000_0000_0000_0000;
array[12479] <= 16'b0000_0000_0000_0000;
array[12480] <= 16'b0000_0000_0000_0000;
array[12481] <= 16'b0000_0000_0000_0000;
array[12482] <= 16'b0000_0000_0000_0000;
array[12483] <= 16'b0000_0000_0000_0000;
array[12484] <= 16'b0000_0000_0000_0000;
array[12485] <= 16'b0000_0000_0000_0000;
array[12486] <= 16'b0000_0000_0000_0000;
array[12487] <= 16'b0000_0000_0000_0000;
array[12488] <= 16'b0000_0000_0000_0000;
array[12489] <= 16'b0000_0000_0000_0000;
array[12490] <= 16'b0000_0000_0000_0000;
array[12491] <= 16'b0000_0000_0000_0000;
array[12492] <= 16'b0000_0000_0000_0000;
array[12493] <= 16'b0000_0000_0000_0000;
array[12494] <= 16'b0000_0000_0000_0000;
array[12495] <= 16'b0000_0000_0000_0000;
array[12496] <= 16'b0000_0000_0000_0000;
array[12497] <= 16'b0000_0000_0000_0000;
array[12498] <= 16'b0000_0000_0000_0000;
array[12499] <= 16'b0000_0000_0000_0000;
array[12500] <= 16'b0000_0000_0000_0000;
array[12501] <= 16'b0000_0000_0000_0000;
array[12502] <= 16'b0000_0000_0000_0000;
array[12503] <= 16'b0000_0000_0000_0000;
array[12504] <= 16'b0000_0000_0000_0000;
array[12505] <= 16'b0000_0000_0000_0000;
array[12506] <= 16'b0000_0000_0000_0000;
array[12507] <= 16'b0000_0000_0000_0000;
array[12508] <= 16'b0000_0000_0000_0000;
array[12509] <= 16'b0000_0000_0000_0000;
array[12510] <= 16'b0000_0000_0000_0000;
array[12511] <= 16'b0000_0000_0000_0000;
array[12512] <= 16'b0000_0000_0000_0000;
array[12513] <= 16'b0000_0000_0000_0000;
array[12514] <= 16'b0000_0000_0000_0000;
array[12515] <= 16'b0000_0000_0000_0000;
array[12516] <= 16'b0000_0000_0000_0000;
array[12517] <= 16'b0000_0000_0000_0000;
array[12518] <= 16'b0000_0000_0000_0000;
array[12519] <= 16'b0000_0000_0000_0000;
array[12520] <= 16'b0000_0000_0000_0000;
array[12521] <= 16'b0000_0000_0000_0000;
array[12522] <= 16'b0000_0000_0000_0000;
array[12523] <= 16'b0000_0000_0000_0000;
array[12524] <= 16'b0000_0000_0000_0000;
array[12525] <= 16'b0000_0000_0000_0000;
array[12526] <= 16'b0000_0000_0000_0000;
array[12527] <= 16'b0000_0000_0000_0000;
array[12528] <= 16'b0000_0000_0000_0000;
array[12529] <= 16'b0000_0000_0000_0000;
array[12530] <= 16'b0000_0000_0000_0000;
array[12531] <= 16'b0000_0000_0000_0000;
array[12532] <= 16'b0000_0000_0000_0000;
array[12533] <= 16'b0000_0000_0000_0000;
array[12534] <= 16'b0000_0000_0000_0000;
array[12535] <= 16'b0000_0000_0000_0000;
array[12536] <= 16'b0000_0000_0000_0000;
array[12537] <= 16'b0000_0000_0000_0000;
array[12538] <= 16'b0000_0000_0000_0000;
array[12539] <= 16'b0000_0000_0000_0000;
array[12540] <= 16'b0000_0000_0000_0000;
array[12541] <= 16'b0000_0000_0000_0000;
array[12542] <= 16'b0000_0000_0000_0000;
array[12543] <= 16'b0000_0000_0000_0000;
array[12544] <= 16'b0000_0000_0000_0000;
array[12545] <= 16'b0000_0000_0000_0000;
array[12546] <= 16'b0000_0000_0000_0000;
array[12547] <= 16'b0000_0000_0000_0000;
array[12548] <= 16'b0000_0000_0000_0000;
array[12549] <= 16'b0000_0000_0000_0000;
array[12550] <= 16'b0000_0000_0000_0000;
array[12551] <= 16'b0000_0000_0000_0000;
array[12552] <= 16'b0000_0000_0000_0000;
array[12553] <= 16'b0000_0000_0000_0000;
array[12554] <= 16'b0000_0000_0000_0000;
array[12555] <= 16'b0000_0000_0000_0000;
array[12556] <= 16'b0000_0000_0000_0000;
array[12557] <= 16'b0000_0000_0000_0000;
array[12558] <= 16'b0000_0000_0000_0000;
array[12559] <= 16'b0000_0000_0000_0000;
array[12560] <= 16'b0000_0000_0000_0000;
array[12561] <= 16'b0000_0000_0000_0000;
array[12562] <= 16'b0000_0000_0000_0000;
array[12563] <= 16'b0000_0000_0000_0000;
array[12564] <= 16'b0000_0000_0000_0000;
array[12565] <= 16'b0000_0000_0000_0000;
array[12566] <= 16'b0000_0000_0000_0000;
array[12567] <= 16'b0000_0000_0000_0000;
array[12568] <= 16'b0000_0000_0000_0000;
array[12569] <= 16'b0000_0000_0000_0000;
array[12570] <= 16'b0000_0000_0000_0000;
array[12571] <= 16'b0000_0000_0000_0000;
array[12572] <= 16'b0000_0000_0000_0000;
array[12573] <= 16'b0000_0000_0000_0000;
array[12574] <= 16'b0000_0000_0000_0000;
array[12575] <= 16'b0000_0000_0000_0000;
array[12576] <= 16'b0000_0000_0000_0000;
array[12577] <= 16'b0000_0000_0000_0000;
array[12578] <= 16'b0000_0000_0000_0000;
array[12579] <= 16'b0000_0000_0000_0000;
array[12580] <= 16'b0000_0000_0000_0000;
array[12581] <= 16'b0000_0000_0000_0000;
array[12582] <= 16'b0000_0000_0000_0000;
array[12583] <= 16'b0000_0000_0000_0000;
array[12584] <= 16'b0000_0000_0000_0000;
array[12585] <= 16'b0000_0000_0000_0000;
array[12586] <= 16'b0000_0000_0000_0000;
array[12587] <= 16'b0000_0000_0000_0000;
array[12588] <= 16'b0000_0000_0000_0000;
array[12589] <= 16'b0000_0000_0000_0000;
array[12590] <= 16'b0000_0000_0000_0000;
array[12591] <= 16'b0000_0000_0000_0000;
array[12592] <= 16'b0000_0000_0000_0000;
array[12593] <= 16'b0000_0000_0000_0000;
array[12594] <= 16'b0000_0000_0000_0000;
array[12595] <= 16'b0000_0000_0000_0000;
array[12596] <= 16'b0000_0000_0000_0000;
array[12597] <= 16'b0000_0000_0000_0000;
array[12598] <= 16'b0000_0000_0000_0000;
array[12599] <= 16'b0000_0000_0000_0000;
array[12600] <= 16'b0000_0000_0000_0000;
array[12601] <= 16'b0000_0000_0000_0000;
array[12602] <= 16'b0000_0000_0000_0000;
array[12603] <= 16'b0000_0000_0000_0000;
array[12604] <= 16'b0000_0000_0000_0000;
array[12605] <= 16'b0000_0000_0000_0000;
array[12606] <= 16'b0000_0000_0000_0000;
array[12607] <= 16'b0000_0000_0000_0000;
array[12608] <= 16'b0000_0000_0000_0000;
array[12609] <= 16'b0000_0000_0000_0000;
array[12610] <= 16'b0000_0000_0000_0000;
array[12611] <= 16'b0000_0000_0000_0000;
array[12612] <= 16'b0000_0000_0000_0000;
array[12613] <= 16'b0000_0000_0000_0000;
array[12614] <= 16'b0000_0000_0000_0000;
array[12615] <= 16'b0000_0000_0000_0000;
array[12616] <= 16'b0000_0000_0000_0000;
array[12617] <= 16'b0000_0000_0000_0000;
array[12618] <= 16'b0000_0000_0000_0000;
array[12619] <= 16'b0000_0000_0000_0000;
array[12620] <= 16'b0000_0000_0000_0000;
array[12621] <= 16'b0000_0000_0000_0000;
array[12622] <= 16'b0000_0000_0000_0000;
array[12623] <= 16'b0000_0000_0000_0000;
array[12624] <= 16'b0000_0000_0000_0000;
array[12625] <= 16'b0000_0000_0000_0000;
array[12626] <= 16'b0000_0000_0000_0000;
array[12627] <= 16'b0000_0000_0000_0000;
array[12628] <= 16'b0000_0000_0000_0000;
array[12629] <= 16'b0000_0000_0000_0000;
array[12630] <= 16'b0000_0000_0000_0000;
array[12631] <= 16'b0000_0000_0000_0000;
array[12632] <= 16'b0000_0000_0000_0000;
array[12633] <= 16'b0000_0000_0000_0000;
array[12634] <= 16'b0000_0000_0000_0000;
array[12635] <= 16'b0000_0000_0000_0000;
array[12636] <= 16'b0000_0000_0000_0000;
array[12637] <= 16'b0000_0000_0000_0000;
array[12638] <= 16'b0000_0000_0000_0000;
array[12639] <= 16'b0000_0000_0000_0000;
array[12640] <= 16'b0000_0000_0000_0000;
array[12641] <= 16'b0000_0000_0000_0000;
array[12642] <= 16'b0000_0000_0000_0000;
array[12643] <= 16'b0000_0000_0000_0000;
array[12644] <= 16'b0000_0000_0000_0000;
array[12645] <= 16'b0000_0000_0000_0000;
array[12646] <= 16'b0000_0000_0000_0000;
array[12647] <= 16'b0000_0000_0000_0000;
array[12648] <= 16'b0000_0000_0000_0000;
array[12649] <= 16'b0000_0000_0000_0000;
array[12650] <= 16'b0000_0000_0000_0000;
array[12651] <= 16'b0000_0000_0000_0000;
array[12652] <= 16'b0000_0000_0000_0000;
array[12653] <= 16'b0000_0000_0000_0000;
array[12654] <= 16'b0000_0000_0000_0000;
array[12655] <= 16'b0000_0000_0000_0000;
array[12656] <= 16'b0000_0000_0000_0000;
array[12657] <= 16'b0000_0000_0000_0000;
array[12658] <= 16'b0000_0000_0000_0000;
array[12659] <= 16'b0000_0000_0000_0000;
array[12660] <= 16'b0000_0000_0000_0000;
array[12661] <= 16'b0000_0000_0000_0000;
array[12662] <= 16'b0000_0000_0000_0000;
array[12663] <= 16'b0000_0000_0000_0000;
array[12664] <= 16'b0000_0000_0000_0000;
array[12665] <= 16'b0000_0000_0000_0000;
array[12666] <= 16'b0000_0000_0000_0000;
array[12667] <= 16'b0000_0000_0000_0000;
array[12668] <= 16'b0000_0000_0000_0000;
array[12669] <= 16'b0000_0000_0000_0000;
array[12670] <= 16'b0000_0000_0000_0000;
array[12671] <= 16'b0000_0000_0000_0000;
array[12672] <= 16'b0000_0000_0000_0000;
array[12673] <= 16'b0000_0000_0000_0000;
array[12674] <= 16'b0000_0000_0000_0000;
array[12675] <= 16'b0000_0000_0000_0000;
array[12676] <= 16'b0000_0000_0000_0000;
array[12677] <= 16'b0000_0000_0000_0000;
array[12678] <= 16'b0000_0000_0000_0000;
array[12679] <= 16'b0000_0000_0000_0000;
array[12680] <= 16'b0000_0000_0000_0000;
array[12681] <= 16'b0000_0000_0000_0000;
array[12682] <= 16'b0000_0000_0000_0000;
array[12683] <= 16'b0000_0000_0000_0000;
array[12684] <= 16'b0000_0000_0000_0000;
array[12685] <= 16'b0000_0000_0000_0000;
array[12686] <= 16'b0000_0000_0000_0000;
array[12687] <= 16'b0000_0000_0000_0000;
array[12688] <= 16'b0000_0000_0000_0000;
array[12689] <= 16'b0000_0000_0000_0000;
array[12690] <= 16'b0000_0000_0000_0000;
array[12691] <= 16'b0000_0000_0000_0000;
array[12692] <= 16'b0000_0000_0000_0000;
array[12693] <= 16'b0000_0000_0000_0000;
array[12694] <= 16'b0000_0000_0000_0000;
array[12695] <= 16'b0000_0000_0000_0000;
array[12696] <= 16'b0000_0000_0000_0000;
array[12697] <= 16'b0000_0000_0000_0000;
array[12698] <= 16'b0000_0000_0000_0000;
array[12699] <= 16'b0000_0000_0000_0000;
array[12700] <= 16'b0000_0000_0000_0000;
array[12701] <= 16'b0000_0000_0000_0000;
array[12702] <= 16'b0000_0000_0000_0000;
array[12703] <= 16'b0000_0000_0000_0000;
array[12704] <= 16'b0000_0000_0000_0000;
array[12705] <= 16'b0000_0000_0000_0000;
array[12706] <= 16'b0000_0000_0000_0000;
array[12707] <= 16'b0000_0000_0000_0000;
array[12708] <= 16'b0000_0000_0000_0000;
array[12709] <= 16'b0000_0000_0000_0000;
array[12710] <= 16'b0000_0000_0000_0000;
array[12711] <= 16'b0000_0000_0000_0000;
array[12712] <= 16'b0000_0000_0000_0000;
array[12713] <= 16'b0000_0000_0000_0000;
array[12714] <= 16'b0000_0000_0000_0000;
array[12715] <= 16'b0000_0000_0000_0000;
array[12716] <= 16'b0000_0000_0000_0000;
array[12717] <= 16'b0000_0000_0000_0000;
array[12718] <= 16'b0000_0000_0000_0000;
array[12719] <= 16'b0000_0000_0000_0000;
array[12720] <= 16'b0000_0000_0000_0000;
array[12721] <= 16'b0000_0000_0000_0000;
array[12722] <= 16'b0000_0000_0000_0000;
array[12723] <= 16'b0000_0000_0000_0000;
array[12724] <= 16'b0000_0000_0000_0000;
array[12725] <= 16'b0000_0000_0000_0000;
array[12726] <= 16'b0000_0000_0000_0000;
array[12727] <= 16'b0000_0000_0000_0000;
array[12728] <= 16'b0000_0000_0000_0000;
array[12729] <= 16'b0000_0000_0000_0000;
array[12730] <= 16'b0000_0000_0000_0000;
array[12731] <= 16'b0000_0000_0000_0000;
array[12732] <= 16'b0000_0000_0000_0000;
array[12733] <= 16'b0000_0000_0000_0000;
array[12734] <= 16'b0000_0000_0000_0000;
array[12735] <= 16'b0000_0000_0000_0000;
array[12736] <= 16'b0000_0000_0000_0000;
array[12737] <= 16'b0000_0000_0000_0000;
array[12738] <= 16'b0000_0000_0000_0000;
array[12739] <= 16'b0000_0000_0000_0000;
array[12740] <= 16'b0000_0000_0000_0000;
array[12741] <= 16'b0000_0000_0000_0000;
array[12742] <= 16'b0000_0000_0000_0000;
array[12743] <= 16'b0000_0000_0000_0000;
array[12744] <= 16'b0000_0000_0000_0000;
array[12745] <= 16'b0000_0000_0000_0000;
array[12746] <= 16'b0000_0000_0000_0000;
array[12747] <= 16'b0000_0000_0000_0000;
array[12748] <= 16'b0000_0000_0000_0000;
array[12749] <= 16'b0000_0000_0000_0000;
array[12750] <= 16'b0000_0000_0000_0000;
array[12751] <= 16'b0000_0000_0000_0000;
array[12752] <= 16'b0000_0000_0000_0000;
array[12753] <= 16'b0000_0000_0000_0000;
array[12754] <= 16'b0000_0000_0000_0000;
array[12755] <= 16'b0000_0000_0000_0000;
array[12756] <= 16'b0000_0000_0000_0000;
array[12757] <= 16'b0000_0000_0000_0000;
array[12758] <= 16'b0000_0000_0000_0000;
array[12759] <= 16'b0000_0000_0000_0000;
array[12760] <= 16'b0000_0000_0000_0000;
array[12761] <= 16'b0000_0000_0000_0000;
array[12762] <= 16'b0000_0000_0000_0000;
array[12763] <= 16'b0000_0000_0000_0000;
array[12764] <= 16'b0000_0000_0000_0000;
array[12765] <= 16'b0000_0000_0000_0000;
array[12766] <= 16'b0000_0000_0000_0000;
array[12767] <= 16'b0000_0000_0000_0000;
array[12768] <= 16'b0000_0000_0000_0000;
array[12769] <= 16'b0000_0000_0000_0000;
array[12770] <= 16'b0000_0000_0000_0000;
array[12771] <= 16'b0000_0000_0000_0000;
array[12772] <= 16'b0000_0000_0000_0000;
array[12773] <= 16'b0000_0000_0000_0000;
array[12774] <= 16'b0000_0000_0000_0000;
array[12775] <= 16'b0000_0000_0000_0000;
array[12776] <= 16'b0000_0000_0000_0000;
array[12777] <= 16'b0000_0000_0000_0000;
array[12778] <= 16'b0000_0000_0000_0000;
array[12779] <= 16'b0000_0000_0000_0000;
array[12780] <= 16'b0000_0000_0000_0000;
array[12781] <= 16'b0000_0000_0000_0000;
array[12782] <= 16'b0000_0000_0000_0000;
array[12783] <= 16'b0000_0000_0000_0000;
array[12784] <= 16'b0000_0000_0000_0000;
array[12785] <= 16'b0000_0000_0000_0000;
array[12786] <= 16'b0000_0000_0000_0000;
array[12787] <= 16'b0000_0000_0000_0000;
array[12788] <= 16'b0000_0000_0000_0000;
array[12789] <= 16'b0000_0000_0000_0000;
array[12790] <= 16'b0000_0000_0000_0000;
array[12791] <= 16'b0000_0000_0000_0000;
array[12792] <= 16'b0000_0000_0000_0000;
array[12793] <= 16'b0000_0000_0000_0000;
array[12794] <= 16'b0000_0000_0000_0000;
array[12795] <= 16'b0000_0000_0000_0000;
array[12796] <= 16'b0000_0000_0000_0000;
array[12797] <= 16'b0000_0000_0000_0000;
array[12798] <= 16'b0000_0000_0000_0000;
array[12799] <= 16'b0000_0000_0000_0000;
array[12800] <= 16'b0000_0000_0000_0000;
array[12801] <= 16'b0000_0000_0000_0000;
array[12802] <= 16'b0000_0000_0000_0000;
array[12803] <= 16'b0000_0000_0000_0000;
array[12804] <= 16'b0000_0000_0000_0000;
array[12805] <= 16'b0000_0000_0000_0000;
array[12806] <= 16'b0000_0000_0000_0000;
array[12807] <= 16'b0000_0000_0000_0000;
array[12808] <= 16'b0000_0000_0000_0000;
array[12809] <= 16'b0000_0000_0000_0000;
array[12810] <= 16'b0000_0000_0000_0000;
array[12811] <= 16'b0000_0000_0000_0000;
array[12812] <= 16'b0000_0000_0000_0000;
array[12813] <= 16'b0000_0000_0000_0000;
array[12814] <= 16'b0000_0000_0000_0000;
array[12815] <= 16'b0000_0000_0000_0000;
array[12816] <= 16'b0000_0000_0000_0000;
array[12817] <= 16'b0000_0000_0000_0000;
array[12818] <= 16'b0000_0000_0000_0000;
array[12819] <= 16'b0000_0000_0000_0000;
array[12820] <= 16'b0000_0000_0000_0000;
array[12821] <= 16'b0000_0000_0000_0000;
array[12822] <= 16'b0000_0000_0000_0000;
array[12823] <= 16'b0000_0000_0000_0000;
array[12824] <= 16'b0000_0000_0000_0000;
array[12825] <= 16'b0000_0000_0000_0000;
array[12826] <= 16'b0000_0000_0000_0000;
array[12827] <= 16'b0000_0000_0000_0000;
array[12828] <= 16'b0000_0000_0000_0000;
array[12829] <= 16'b0000_0000_0000_0000;
array[12830] <= 16'b0000_0000_0000_0000;
array[12831] <= 16'b0000_0000_0000_0000;
array[12832] <= 16'b0000_0000_0000_0000;
array[12833] <= 16'b0000_0000_0000_0000;
array[12834] <= 16'b0000_0000_0000_0000;
array[12835] <= 16'b0000_0000_0000_0000;
array[12836] <= 16'b0000_0000_0000_0000;
array[12837] <= 16'b0000_0000_0000_0000;
array[12838] <= 16'b0000_0000_0000_0000;
array[12839] <= 16'b0000_0000_0000_0000;
array[12840] <= 16'b0000_0000_0000_0000;
array[12841] <= 16'b0000_0000_0000_0000;
array[12842] <= 16'b0000_0000_0000_0000;
array[12843] <= 16'b0000_0000_0000_0000;
array[12844] <= 16'b0000_0000_0000_0000;
array[12845] <= 16'b0000_0000_0000_0000;
array[12846] <= 16'b0000_0000_0000_0000;
array[12847] <= 16'b0000_0000_0000_0000;
array[12848] <= 16'b0000_0000_0000_0000;
array[12849] <= 16'b0000_0000_0000_0000;
array[12850] <= 16'b0000_0000_0000_0000;
array[12851] <= 16'b0000_0000_0000_0000;
array[12852] <= 16'b0000_0000_0000_0000;
array[12853] <= 16'b0000_0000_0000_0000;
array[12854] <= 16'b0000_0000_0000_0000;
array[12855] <= 16'b0000_0000_0000_0000;
array[12856] <= 16'b0000_0000_0000_0000;
array[12857] <= 16'b0000_0000_0000_0000;
array[12858] <= 16'b0000_0000_0000_0000;
array[12859] <= 16'b0000_0000_0000_0000;
array[12860] <= 16'b0000_0000_0000_0000;
array[12861] <= 16'b0000_0000_0000_0000;
array[12862] <= 16'b0000_0000_0000_0000;
array[12863] <= 16'b0000_0000_0000_0000;
array[12864] <= 16'b0000_0000_0000_0000;
array[12865] <= 16'b0000_0000_0000_0000;
array[12866] <= 16'b0000_0000_0000_0000;
array[12867] <= 16'b0000_0000_0000_0000;
array[12868] <= 16'b0000_0000_0000_0000;
array[12869] <= 16'b0000_0000_0000_0000;
array[12870] <= 16'b0000_0000_0000_0000;
array[12871] <= 16'b0000_0000_0000_0000;
array[12872] <= 16'b0000_0000_0000_0000;
array[12873] <= 16'b0000_0000_0000_0000;
array[12874] <= 16'b0000_0000_0000_0000;
array[12875] <= 16'b0000_0000_0000_0000;
array[12876] <= 16'b0000_0000_0000_0000;
array[12877] <= 16'b0000_0000_0000_0000;
array[12878] <= 16'b0000_0000_0000_0000;
array[12879] <= 16'b0000_0000_0000_0000;
array[12880] <= 16'b0000_0000_0000_0000;
array[12881] <= 16'b0000_0000_0000_0000;
array[12882] <= 16'b0000_0000_0000_0000;
array[12883] <= 16'b0000_0000_0000_0000;
array[12884] <= 16'b0000_0000_0000_0000;
array[12885] <= 16'b0000_0000_0000_0000;
array[12886] <= 16'b0000_0000_0000_0000;
array[12887] <= 16'b0000_0000_0000_0000;
array[12888] <= 16'b0000_0000_0000_0000;
array[12889] <= 16'b0000_0000_0000_0000;
array[12890] <= 16'b0000_0000_0000_0000;
array[12891] <= 16'b0000_0000_0000_0000;
array[12892] <= 16'b0000_0000_0000_0000;
array[12893] <= 16'b0000_0000_0000_0000;
array[12894] <= 16'b0000_0000_0000_0000;
array[12895] <= 16'b0000_0000_0000_0000;
array[12896] <= 16'b0000_0000_0000_0000;
array[12897] <= 16'b0000_0000_0000_0000;
array[12898] <= 16'b0000_0000_0000_0000;
array[12899] <= 16'b0000_0000_0000_0000;
array[12900] <= 16'b0000_0000_0000_0000;
array[12901] <= 16'b0000_0000_0000_0000;
array[12902] <= 16'b0000_0000_0000_0000;
array[12903] <= 16'b0000_0000_0000_0000;
array[12904] <= 16'b0000_0000_0000_0000;
array[12905] <= 16'b0000_0000_0000_0000;
array[12906] <= 16'b0000_0000_0000_0000;
array[12907] <= 16'b0000_0000_0000_0000;
array[12908] <= 16'b0000_0000_0000_0000;
array[12909] <= 16'b0000_0000_0000_0000;
array[12910] <= 16'b0000_0000_0000_0000;
array[12911] <= 16'b0000_0000_0000_0000;
array[12912] <= 16'b0000_0000_0000_0000;
array[12913] <= 16'b0000_0000_0000_0000;
array[12914] <= 16'b0000_0000_0000_0000;
array[12915] <= 16'b0000_0000_0000_0000;
array[12916] <= 16'b0000_0000_0000_0000;
array[12917] <= 16'b0000_0000_0000_0000;
array[12918] <= 16'b0000_0000_0000_0000;
array[12919] <= 16'b0000_0000_0000_0000;
array[12920] <= 16'b0000_0000_0000_0000;
array[12921] <= 16'b0000_0000_0000_0000;
array[12922] <= 16'b0000_0000_0000_0000;
array[12923] <= 16'b0000_0000_0000_0000;
array[12924] <= 16'b0000_0000_0000_0000;
array[12925] <= 16'b0000_0000_0000_0000;
array[12926] <= 16'b0000_0000_0000_0000;
array[12927] <= 16'b0000_0000_0000_0000;
array[12928] <= 16'b0000_0000_0000_0000;
array[12929] <= 16'b0000_0000_0000_0000;
array[12930] <= 16'b0000_0000_0000_0000;
array[12931] <= 16'b0000_0000_0000_0000;
array[12932] <= 16'b0000_0000_0000_0000;
array[12933] <= 16'b0000_0000_0000_0000;
array[12934] <= 16'b0000_0000_0000_0000;
array[12935] <= 16'b0000_0000_0000_0000;
array[12936] <= 16'b0000_0000_0000_0000;
array[12937] <= 16'b0000_0000_0000_0000;
array[12938] <= 16'b0000_0000_0000_0000;
array[12939] <= 16'b0000_0000_0000_0000;
array[12940] <= 16'b0000_0000_0000_0000;
array[12941] <= 16'b0000_0000_0000_0000;
array[12942] <= 16'b0000_0000_0000_0000;
array[12943] <= 16'b0000_0000_0000_0000;
array[12944] <= 16'b0000_0000_0000_0000;
array[12945] <= 16'b0000_0000_0000_0000;
array[12946] <= 16'b0000_0000_0000_0000;
array[12947] <= 16'b0000_0000_0000_0000;
array[12948] <= 16'b0000_0000_0000_0000;
array[12949] <= 16'b0000_0000_0000_0000;
array[12950] <= 16'b0000_0000_0000_0000;
array[12951] <= 16'b0000_0000_0000_0000;
array[12952] <= 16'b0000_0000_0000_0000;
array[12953] <= 16'b0000_0000_0000_0000;
array[12954] <= 16'b0000_0000_0000_0000;
array[12955] <= 16'b0000_0000_0000_0000;
array[12956] <= 16'b0000_0000_0000_0000;
array[12957] <= 16'b0000_0000_0000_0000;
array[12958] <= 16'b0000_0000_0000_0000;
array[12959] <= 16'b0000_0000_0000_0000;
array[12960] <= 16'b0000_0000_0000_0000;
array[12961] <= 16'b0000_0000_0000_0000;
array[12962] <= 16'b0000_0000_0000_0000;
array[12963] <= 16'b0000_0000_0000_0000;
array[12964] <= 16'b0000_0000_0000_0000;
array[12965] <= 16'b0000_0000_0000_0000;
array[12966] <= 16'b0000_0000_0000_0000;
array[12967] <= 16'b0000_0000_0000_0000;
array[12968] <= 16'b0000_0000_0000_0000;
array[12969] <= 16'b0000_0000_0000_0000;
array[12970] <= 16'b0000_0000_0000_0000;
array[12971] <= 16'b0000_0000_0000_0000;
array[12972] <= 16'b0000_0000_0000_0000;
array[12973] <= 16'b0000_0000_0000_0000;
array[12974] <= 16'b0000_0000_0000_0000;
array[12975] <= 16'b0000_0000_0000_0000;
array[12976] <= 16'b0000_0000_0000_0000;
array[12977] <= 16'b0000_0000_0000_0000;
array[12978] <= 16'b0000_0000_0000_0000;
array[12979] <= 16'b0000_0000_0000_0000;
array[12980] <= 16'b0000_0000_0000_0000;
array[12981] <= 16'b0000_0000_0000_0000;
array[12982] <= 16'b0000_0000_0000_0000;
array[12983] <= 16'b0000_0000_0000_0000;
array[12984] <= 16'b0000_0000_0000_0000;
array[12985] <= 16'b0000_0000_0000_0000;
array[12986] <= 16'b0000_0000_0000_0000;
array[12987] <= 16'b0000_0000_0000_0000;
array[12988] <= 16'b0000_0000_0000_0000;
array[12989] <= 16'b0000_0000_0000_0000;
array[12990] <= 16'b0000_0000_0000_0000;
array[12991] <= 16'b0000_0000_0000_0000;
array[12992] <= 16'b0000_0000_0000_0000;
array[12993] <= 16'b0000_0000_0000_0000;
array[12994] <= 16'b0000_0000_0000_0000;
array[12995] <= 16'b0000_0000_0000_0000;
array[12996] <= 16'b0000_0000_0000_0000;
array[12997] <= 16'b0000_0000_0000_0000;
array[12998] <= 16'b0000_0000_0000_0000;
array[12999] <= 16'b0000_0000_0000_0000;
array[13000] <= 16'b0000_0000_0000_0000;
array[13001] <= 16'b0000_0000_0000_0000;
array[13002] <= 16'b0000_0000_0000_0000;
array[13003] <= 16'b0000_0000_0000_0000;
array[13004] <= 16'b0000_0000_0000_0000;
array[13005] <= 16'b0000_0000_0000_0000;
array[13006] <= 16'b0000_0000_0000_0000;
array[13007] <= 16'b0000_0000_0000_0000;
array[13008] <= 16'b0000_0000_0000_0000;
array[13009] <= 16'b0000_0000_0000_0000;
array[13010] <= 16'b0000_0000_0000_0000;
array[13011] <= 16'b0000_0000_0000_0000;
array[13012] <= 16'b0000_0000_0000_0000;
array[13013] <= 16'b0000_0000_0000_0000;
array[13014] <= 16'b0000_0000_0000_0000;
array[13015] <= 16'b0000_0000_0000_0000;
array[13016] <= 16'b0000_0000_0000_0000;
array[13017] <= 16'b0000_0000_0000_0000;
array[13018] <= 16'b0000_0000_0000_0000;
array[13019] <= 16'b0000_0000_0000_0000;
array[13020] <= 16'b0000_0000_0000_0000;
array[13021] <= 16'b0000_0000_0000_0000;
array[13022] <= 16'b0000_0000_0000_0000;
array[13023] <= 16'b0000_0000_0000_0000;
array[13024] <= 16'b0000_0000_0000_0000;
array[13025] <= 16'b0000_0000_0000_0000;
array[13026] <= 16'b0000_0000_0000_0000;
array[13027] <= 16'b0000_0000_0000_0000;
array[13028] <= 16'b0000_0000_0000_0000;
array[13029] <= 16'b0000_0000_0000_0000;
array[13030] <= 16'b0000_0000_0000_0000;
array[13031] <= 16'b0000_0000_0000_0000;
array[13032] <= 16'b0000_0000_0000_0000;
array[13033] <= 16'b0000_0000_0000_0000;
array[13034] <= 16'b0000_0000_0000_0000;
array[13035] <= 16'b0000_0000_0000_0000;
array[13036] <= 16'b0000_0000_0000_0000;
array[13037] <= 16'b0000_0000_0000_0000;
array[13038] <= 16'b0000_0000_0000_0000;
array[13039] <= 16'b0000_0000_0000_0000;
array[13040] <= 16'b0000_0000_0000_0000;
array[13041] <= 16'b0000_0000_0000_0000;
array[13042] <= 16'b0000_0000_0000_0000;
array[13043] <= 16'b0000_0000_0000_0000;
array[13044] <= 16'b0000_0000_0000_0000;
array[13045] <= 16'b0000_0000_0000_0000;
array[13046] <= 16'b0000_0000_0000_0000;
array[13047] <= 16'b0000_0000_0000_0000;
array[13048] <= 16'b0000_0000_0000_0000;
array[13049] <= 16'b0000_0000_0000_0000;
array[13050] <= 16'b0000_0000_0000_0000;
array[13051] <= 16'b0000_0000_0000_0000;
array[13052] <= 16'b0000_0000_0000_0000;
array[13053] <= 16'b0000_0000_0000_0000;
array[13054] <= 16'b0000_0000_0000_0000;
array[13055] <= 16'b0000_0000_0000_0000;
array[13056] <= 16'b0000_0000_0000_0000;
array[13057] <= 16'b0000_0000_0000_0000;
array[13058] <= 16'b0000_0000_0000_0000;
array[13059] <= 16'b0000_0000_0000_0000;
array[13060] <= 16'b0000_0000_0000_0000;
array[13061] <= 16'b0000_0000_0000_0000;
array[13062] <= 16'b0000_0000_0000_0000;
array[13063] <= 16'b0000_0000_0000_0000;
array[13064] <= 16'b0000_0000_0000_0000;
array[13065] <= 16'b0000_0000_0000_0000;
array[13066] <= 16'b0000_0000_0000_0000;
array[13067] <= 16'b0000_0000_0000_0000;
array[13068] <= 16'b0000_0000_0000_0000;
array[13069] <= 16'b0000_0000_0000_0000;
array[13070] <= 16'b0000_0000_0000_0000;
array[13071] <= 16'b0000_0000_0000_0000;
array[13072] <= 16'b0000_0000_0000_0000;
array[13073] <= 16'b0000_0000_0000_0000;
array[13074] <= 16'b0000_0000_0000_0000;
array[13075] <= 16'b0000_0000_0000_0000;
array[13076] <= 16'b0000_0000_0000_0000;
array[13077] <= 16'b0000_0000_0000_0000;
array[13078] <= 16'b0000_0000_0000_0000;
array[13079] <= 16'b0000_0000_0000_0000;
array[13080] <= 16'b0000_0000_0000_0000;
array[13081] <= 16'b0000_0000_0000_0000;
array[13082] <= 16'b0000_0000_0000_0000;
array[13083] <= 16'b0000_0000_0000_0000;
array[13084] <= 16'b0000_0000_0000_0000;
array[13085] <= 16'b0000_0000_0000_0000;
array[13086] <= 16'b0000_0000_0000_0000;
array[13087] <= 16'b0000_0000_0000_0000;
array[13088] <= 16'b0000_0000_0000_0000;
array[13089] <= 16'b0000_0000_0000_0000;
array[13090] <= 16'b0000_0000_0000_0000;
array[13091] <= 16'b0000_0000_0000_0000;
array[13092] <= 16'b0000_0000_0000_0000;
array[13093] <= 16'b0000_0000_0000_0000;
array[13094] <= 16'b0000_0000_0000_0000;
array[13095] <= 16'b0000_0000_0000_0000;
array[13096] <= 16'b0000_0000_0000_0000;
array[13097] <= 16'b0000_0000_0000_0000;
array[13098] <= 16'b0000_0000_0000_0000;
array[13099] <= 16'b0000_0000_0000_0000;
array[13100] <= 16'b0000_0000_0000_0000;
array[13101] <= 16'b0000_0000_0000_0000;
array[13102] <= 16'b0000_0000_0000_0000;
array[13103] <= 16'b0000_0000_0000_0000;
array[13104] <= 16'b0000_0000_0000_0000;
array[13105] <= 16'b0000_0000_0000_0000;
array[13106] <= 16'b0000_0000_0000_0000;
array[13107] <= 16'b0000_0000_0000_0000;
array[13108] <= 16'b0000_0000_0000_0000;
array[13109] <= 16'b0000_0000_0000_0000;
array[13110] <= 16'b0000_0000_0000_0000;
array[13111] <= 16'b0000_0000_0000_0000;
array[13112] <= 16'b0000_0000_0000_0000;
array[13113] <= 16'b0000_0000_0000_0000;
array[13114] <= 16'b0000_0000_0000_0000;
array[13115] <= 16'b0000_0000_0000_0000;
array[13116] <= 16'b0000_0000_0000_0000;
array[13117] <= 16'b0000_0000_0000_0000;
array[13118] <= 16'b0000_0000_0000_0000;
array[13119] <= 16'b0000_0000_0000_0000;
array[13120] <= 16'b0000_0000_0000_0000;
array[13121] <= 16'b0000_0000_0000_0000;
array[13122] <= 16'b0000_0000_0000_0000;
array[13123] <= 16'b0000_0000_0000_0000;
array[13124] <= 16'b0000_0000_0000_0000;
array[13125] <= 16'b0000_0000_0000_0000;
array[13126] <= 16'b0000_0000_0000_0000;
array[13127] <= 16'b0000_0000_0000_0000;
array[13128] <= 16'b0000_0000_0000_0000;
array[13129] <= 16'b0000_0000_0000_0000;
array[13130] <= 16'b0000_0000_0000_0000;
array[13131] <= 16'b0000_0000_0000_0000;
array[13132] <= 16'b0000_0000_0000_0000;
array[13133] <= 16'b0000_0000_0000_0000;
array[13134] <= 16'b0000_0000_0000_0000;
array[13135] <= 16'b0000_0000_0000_0000;
array[13136] <= 16'b0000_0000_0000_0000;
array[13137] <= 16'b0000_0000_0000_0000;
array[13138] <= 16'b0000_0000_0000_0000;
array[13139] <= 16'b0000_0000_0000_0000;
array[13140] <= 16'b0000_0000_0000_0000;
array[13141] <= 16'b0000_0000_0000_0000;
array[13142] <= 16'b0000_0000_0000_0000;
array[13143] <= 16'b0000_0000_0000_0000;
array[13144] <= 16'b0000_0000_0000_0000;
array[13145] <= 16'b0000_0000_0000_0000;
array[13146] <= 16'b0000_0000_0000_0000;
array[13147] <= 16'b0000_0000_0000_0000;
array[13148] <= 16'b0000_0000_0000_0000;
array[13149] <= 16'b0000_0000_0000_0000;
array[13150] <= 16'b0000_0000_0000_0000;
array[13151] <= 16'b0000_0000_0000_0000;
array[13152] <= 16'b0000_0000_0000_0000;
array[13153] <= 16'b0000_0000_0000_0000;
array[13154] <= 16'b0000_0000_0000_0000;
array[13155] <= 16'b0000_0000_0000_0000;
array[13156] <= 16'b0000_0000_0000_0000;
array[13157] <= 16'b0000_0000_0000_0000;
array[13158] <= 16'b0000_0000_0000_0000;
array[13159] <= 16'b0000_0000_0000_0000;
array[13160] <= 16'b0000_0000_0000_0000;
array[13161] <= 16'b0000_0000_0000_0000;
array[13162] <= 16'b0000_0000_0000_0000;
array[13163] <= 16'b0000_0000_0000_0000;
array[13164] <= 16'b0000_0000_0000_0000;
array[13165] <= 16'b0000_0000_0000_0000;
array[13166] <= 16'b0000_0000_0000_0000;
array[13167] <= 16'b0000_0000_0000_0000;
array[13168] <= 16'b0000_0000_0000_0000;
array[13169] <= 16'b0000_0000_0000_0000;
array[13170] <= 16'b0000_0000_0000_0000;
array[13171] <= 16'b0000_0000_0000_0000;
array[13172] <= 16'b0000_0000_0000_0000;
array[13173] <= 16'b0000_0000_0000_0000;
array[13174] <= 16'b0000_0000_0000_0000;
array[13175] <= 16'b0000_0000_0000_0000;
array[13176] <= 16'b0000_0000_0000_0000;
array[13177] <= 16'b0000_0000_0000_0000;
array[13178] <= 16'b0000_0000_0000_0000;
array[13179] <= 16'b0000_0000_0000_0000;
array[13180] <= 16'b0000_0000_0000_0000;
array[13181] <= 16'b0000_0000_0000_0000;
array[13182] <= 16'b0000_0000_0000_0000;
array[13183] <= 16'b0000_0000_0000_0000;
array[13184] <= 16'b0000_0000_0000_0000;
array[13185] <= 16'b0000_0000_0000_0000;
array[13186] <= 16'b0000_0000_0000_0000;
array[13187] <= 16'b0000_0000_0000_0000;
array[13188] <= 16'b0000_0000_0000_0000;
array[13189] <= 16'b0000_0000_0000_0000;
array[13190] <= 16'b0000_0000_0000_0000;
array[13191] <= 16'b0000_0000_0000_0000;
array[13192] <= 16'b0000_0000_0000_0000;
array[13193] <= 16'b0000_0000_0000_0000;
array[13194] <= 16'b0000_0000_0000_0000;
array[13195] <= 16'b0000_0000_0000_0000;
array[13196] <= 16'b0000_0000_0000_0000;
array[13197] <= 16'b0000_0000_0000_0000;
array[13198] <= 16'b0000_0000_0000_0000;
array[13199] <= 16'b0000_0000_0000_0000;
array[13200] <= 16'b0000_0000_0000_0000;
array[13201] <= 16'b0000_0000_0000_0000;
array[13202] <= 16'b0000_0000_0000_0000;
array[13203] <= 16'b0000_0000_0000_0000;
array[13204] <= 16'b0000_0000_0000_0000;
array[13205] <= 16'b0000_0000_0000_0000;
array[13206] <= 16'b0000_0000_0000_0000;
array[13207] <= 16'b0000_0000_0000_0000;
array[13208] <= 16'b0000_0000_0000_0000;
array[13209] <= 16'b0000_0000_0000_0000;
array[13210] <= 16'b0000_0000_0000_0000;
array[13211] <= 16'b0000_0000_0000_0000;
array[13212] <= 16'b0000_0000_0000_0000;
array[13213] <= 16'b0000_0000_0000_0000;
array[13214] <= 16'b0000_0000_0000_0000;
array[13215] <= 16'b0000_0000_0000_0000;
array[13216] <= 16'b0000_0000_0000_0000;
array[13217] <= 16'b0000_0000_0000_0000;
array[13218] <= 16'b0000_0000_0000_0000;
array[13219] <= 16'b0000_0000_0000_0000;
array[13220] <= 16'b0000_0000_0000_0000;
array[13221] <= 16'b0000_0000_0000_0000;
array[13222] <= 16'b0000_0000_0000_0000;
array[13223] <= 16'b0000_0000_0000_0000;
array[13224] <= 16'b0000_0000_0000_0000;
array[13225] <= 16'b0000_0000_0000_0000;
array[13226] <= 16'b0000_0000_0000_0000;
array[13227] <= 16'b0000_0000_0000_0000;
array[13228] <= 16'b0000_0000_0000_0000;
array[13229] <= 16'b0000_0000_0000_0000;
array[13230] <= 16'b0000_0000_0000_0000;
array[13231] <= 16'b0000_0000_0000_0000;
array[13232] <= 16'b0000_0000_0000_0000;
array[13233] <= 16'b0000_0000_0000_0000;
array[13234] <= 16'b0000_0000_0000_0000;
array[13235] <= 16'b0000_0000_0000_0000;
array[13236] <= 16'b0000_0000_0000_0000;
array[13237] <= 16'b0000_0000_0000_0000;
array[13238] <= 16'b0000_0000_0000_0000;
array[13239] <= 16'b0000_0000_0000_0000;
array[13240] <= 16'b0000_0000_0000_0000;
array[13241] <= 16'b0000_0000_0000_0000;
array[13242] <= 16'b0000_0000_0000_0000;
array[13243] <= 16'b0000_0000_0000_0000;
array[13244] <= 16'b0000_0000_0000_0000;
array[13245] <= 16'b0000_0000_0000_0000;
array[13246] <= 16'b0000_0000_0000_0000;
array[13247] <= 16'b0000_0000_0000_0000;
array[13248] <= 16'b0000_0000_0000_0000;
array[13249] <= 16'b0000_0000_0000_0000;
array[13250] <= 16'b0000_0000_0000_0000;
array[13251] <= 16'b0000_0000_0000_0000;
array[13252] <= 16'b0000_0000_0000_0000;
array[13253] <= 16'b0000_0000_0000_0000;
array[13254] <= 16'b0000_0000_0000_0000;
array[13255] <= 16'b0000_0000_0000_0000;
array[13256] <= 16'b0000_0000_0000_0000;
array[13257] <= 16'b0000_0000_0000_0000;
array[13258] <= 16'b0000_0000_0000_0000;
array[13259] <= 16'b0000_0000_0000_0000;
array[13260] <= 16'b0000_0000_0000_0000;
array[13261] <= 16'b0000_0000_0000_0000;
array[13262] <= 16'b0000_0000_0000_0000;
array[13263] <= 16'b0000_0000_0000_0000;
array[13264] <= 16'b0000_0000_0000_0000;
array[13265] <= 16'b0000_0000_0000_0000;
array[13266] <= 16'b0000_0000_0000_0000;
array[13267] <= 16'b0000_0000_0000_0000;
array[13268] <= 16'b0000_0000_0000_0000;
array[13269] <= 16'b0000_0000_0000_0000;
array[13270] <= 16'b0000_0000_0000_0000;
array[13271] <= 16'b0000_0000_0000_0000;
array[13272] <= 16'b0000_0000_0000_0000;
array[13273] <= 16'b0000_0000_0000_0000;
array[13274] <= 16'b0000_0000_0000_0000;
array[13275] <= 16'b0000_0000_0000_0000;
array[13276] <= 16'b0000_0000_0000_0000;
array[13277] <= 16'b0000_0000_0000_0000;
array[13278] <= 16'b0000_0000_0000_0000;
array[13279] <= 16'b0000_0000_0000_0000;
array[13280] <= 16'b0000_0000_0000_0000;
array[13281] <= 16'b0000_0000_0000_0000;
array[13282] <= 16'b0000_0000_0000_0000;
array[13283] <= 16'b0000_0000_0000_0000;
array[13284] <= 16'b0000_0000_0000_0000;
array[13285] <= 16'b0000_0000_0000_0000;
array[13286] <= 16'b0000_0000_0000_0000;
array[13287] <= 16'b0000_0000_0000_0000;
array[13288] <= 16'b0000_0000_0000_0000;
array[13289] <= 16'b0000_0000_0000_0000;
array[13290] <= 16'b0000_0000_0000_0000;
array[13291] <= 16'b0000_0000_0000_0000;
array[13292] <= 16'b0000_0000_0000_0000;
array[13293] <= 16'b0000_0000_0000_0000;
array[13294] <= 16'b0000_0000_0000_0000;
array[13295] <= 16'b0000_0000_0000_0000;
array[13296] <= 16'b0000_0000_0000_0000;
array[13297] <= 16'b0000_0000_0000_0000;
array[13298] <= 16'b0000_0000_0000_0000;
array[13299] <= 16'b0000_0000_0000_0000;
array[13300] <= 16'b0000_0000_0000_0000;
array[13301] <= 16'b0000_0000_0000_0000;
array[13302] <= 16'b0000_0000_0000_0000;
array[13303] <= 16'b0000_0000_0000_0000;
array[13304] <= 16'b0000_0000_0000_0000;
array[13305] <= 16'b0000_0000_0000_0000;
array[13306] <= 16'b0000_0000_0000_0000;
array[13307] <= 16'b0000_0000_0000_0000;
array[13308] <= 16'b0000_0000_0000_0000;
array[13309] <= 16'b0000_0000_0000_0000;
array[13310] <= 16'b0000_0000_0000_0000;
array[13311] <= 16'b0000_0000_0000_0000;
array[13312] <= 16'b0000_0000_0000_0000;
array[13313] <= 16'b0000_0000_0000_0000;
array[13314] <= 16'b0000_0000_0000_0000;
array[13315] <= 16'b0000_0000_0000_0000;
array[13316] <= 16'b0000_0000_0000_0000;
array[13317] <= 16'b0000_0000_0000_0000;
array[13318] <= 16'b0000_0000_0000_0000;
array[13319] <= 16'b0000_0000_0000_0000;
array[13320] <= 16'b0000_0000_0000_0000;
array[13321] <= 16'b0000_0000_0000_0000;
array[13322] <= 16'b0000_0000_0000_0000;
array[13323] <= 16'b0000_0000_0000_0000;
array[13324] <= 16'b0000_0000_0000_0000;
array[13325] <= 16'b0000_0000_0000_0000;
array[13326] <= 16'b0000_0000_0000_0000;
array[13327] <= 16'b0000_0000_0000_0000;
array[13328] <= 16'b0000_0000_0000_0000;
array[13329] <= 16'b0000_0000_0000_0000;
array[13330] <= 16'b0000_0000_0000_0000;
array[13331] <= 16'b0000_0000_0000_0000;
array[13332] <= 16'b0000_0000_0000_0000;
array[13333] <= 16'b0000_0000_0000_0000;
array[13334] <= 16'b0000_0000_0000_0000;
array[13335] <= 16'b0000_0000_0000_0000;
array[13336] <= 16'b0000_0000_0000_0000;
array[13337] <= 16'b0000_0000_0000_0000;
array[13338] <= 16'b0000_0000_0000_0000;
array[13339] <= 16'b0000_0000_0000_0000;
array[13340] <= 16'b0000_0000_0000_0000;
array[13341] <= 16'b0000_0000_0000_0000;
array[13342] <= 16'b0000_0000_0000_0000;
array[13343] <= 16'b0000_0000_0000_0000;
array[13344] <= 16'b0000_0000_0000_0000;
array[13345] <= 16'b0000_0000_0000_0000;
array[13346] <= 16'b0000_0000_0000_0000;
array[13347] <= 16'b0000_0000_0000_0000;
array[13348] <= 16'b0000_0000_0000_0000;
array[13349] <= 16'b0000_0000_0000_0000;
array[13350] <= 16'b0000_0000_0000_0000;
array[13351] <= 16'b0000_0000_0000_0000;
array[13352] <= 16'b0000_0000_0000_0000;
array[13353] <= 16'b0000_0000_0000_0000;
array[13354] <= 16'b0000_0000_0000_0000;
array[13355] <= 16'b0000_0000_0000_0000;
array[13356] <= 16'b0000_0000_0000_0000;
array[13357] <= 16'b0000_0000_0000_0000;
array[13358] <= 16'b0000_0000_0000_0000;
array[13359] <= 16'b0000_0000_0000_0000;
array[13360] <= 16'b0000_0000_0000_0000;
array[13361] <= 16'b0000_0000_0000_0000;
array[13362] <= 16'b0000_0000_0000_0000;
array[13363] <= 16'b0000_0000_0000_0000;
array[13364] <= 16'b0000_0000_0000_0000;
array[13365] <= 16'b0000_0000_0000_0000;
array[13366] <= 16'b0000_0000_0000_0000;
array[13367] <= 16'b0000_0000_0000_0000;
array[13368] <= 16'b0000_0000_0000_0000;
array[13369] <= 16'b0000_0000_0000_0000;
array[13370] <= 16'b0000_0000_0000_0000;
array[13371] <= 16'b0000_0000_0000_0000;
array[13372] <= 16'b0000_0000_0000_0000;
array[13373] <= 16'b0000_0000_0000_0000;
array[13374] <= 16'b0000_0000_0000_0000;
array[13375] <= 16'b0000_0000_0000_0000;
array[13376] <= 16'b0000_0000_0000_0000;
array[13377] <= 16'b0000_0000_0000_0000;
array[13378] <= 16'b0000_0000_0000_0000;
array[13379] <= 16'b0000_0000_0000_0000;
array[13380] <= 16'b0000_0000_0000_0000;
array[13381] <= 16'b0000_0000_0000_0000;
array[13382] <= 16'b0000_0000_0000_0000;
array[13383] <= 16'b0000_0000_0000_0000;
array[13384] <= 16'b0000_0000_0000_0000;
array[13385] <= 16'b0000_0000_0000_0000;
array[13386] <= 16'b0000_0000_0000_0000;
array[13387] <= 16'b0000_0000_0000_0000;
array[13388] <= 16'b0000_0000_0000_0000;
array[13389] <= 16'b0000_0000_0000_0000;
array[13390] <= 16'b0000_0000_0000_0000;
array[13391] <= 16'b0000_0000_0000_0000;
array[13392] <= 16'b0000_0000_0000_0000;
array[13393] <= 16'b0000_0000_0000_0000;
array[13394] <= 16'b0000_0000_0000_0000;
array[13395] <= 16'b0000_0000_0000_0000;
array[13396] <= 16'b0000_0000_0000_0000;
array[13397] <= 16'b0000_0000_0000_0000;
array[13398] <= 16'b0000_0000_0000_0000;
array[13399] <= 16'b0000_0000_0000_0000;
array[13400] <= 16'b0000_0000_0000_0000;
array[13401] <= 16'b0000_0000_0000_0000;
array[13402] <= 16'b0000_0000_0000_0000;
array[13403] <= 16'b0000_0000_0000_0000;
array[13404] <= 16'b0000_0000_0000_0000;
array[13405] <= 16'b0000_0000_0000_0000;
array[13406] <= 16'b0000_0000_0000_0000;
array[13407] <= 16'b0000_0000_0000_0000;
array[13408] <= 16'b0000_0000_0000_0000;
array[13409] <= 16'b0000_0000_0000_0000;
array[13410] <= 16'b0000_0000_0000_0000;
array[13411] <= 16'b0000_0000_0000_0000;
array[13412] <= 16'b0000_0000_0000_0000;
array[13413] <= 16'b0000_0000_0000_0000;
array[13414] <= 16'b0000_0000_0000_0000;
array[13415] <= 16'b0000_0000_0000_0000;
array[13416] <= 16'b0000_0000_0000_0000;
array[13417] <= 16'b0000_0000_0000_0000;
array[13418] <= 16'b0000_0000_0000_0000;
array[13419] <= 16'b0000_0000_0000_0000;
array[13420] <= 16'b0000_0000_0000_0000;
array[13421] <= 16'b0000_0000_0000_0000;
array[13422] <= 16'b0000_0000_0000_0000;
array[13423] <= 16'b0000_0000_0000_0000;
array[13424] <= 16'b0000_0000_0000_0000;
array[13425] <= 16'b0000_0000_0000_0000;
array[13426] <= 16'b0000_0000_0000_0000;
array[13427] <= 16'b0000_0000_0000_0000;
array[13428] <= 16'b0000_0000_0000_0000;
array[13429] <= 16'b0000_0000_0000_0000;
array[13430] <= 16'b0000_0000_0000_0000;
array[13431] <= 16'b0000_0000_0000_0000;
array[13432] <= 16'b0000_0000_0000_0000;
array[13433] <= 16'b0000_0000_0000_0000;
array[13434] <= 16'b0000_0000_0000_0000;
array[13435] <= 16'b0000_0000_0000_0000;
array[13436] <= 16'b0000_0000_0000_0000;
array[13437] <= 16'b0000_0000_0000_0000;
array[13438] <= 16'b0000_0000_0000_0000;
array[13439] <= 16'b0000_0000_0000_0000;
array[13440] <= 16'b0000_0000_0000_0000;
array[13441] <= 16'b0000_0000_0000_0000;
array[13442] <= 16'b0000_0000_0000_0000;
array[13443] <= 16'b0000_0000_0000_0000;
array[13444] <= 16'b0000_0000_0000_0000;
array[13445] <= 16'b0000_0000_0000_0000;
array[13446] <= 16'b0000_0000_0000_0000;
array[13447] <= 16'b0000_0000_0000_0000;
array[13448] <= 16'b0000_0000_0000_0000;
array[13449] <= 16'b0000_0000_0000_0000;
array[13450] <= 16'b0000_0000_0000_0000;
array[13451] <= 16'b0000_0000_0000_0000;
array[13452] <= 16'b0000_0000_0000_0000;
array[13453] <= 16'b0000_0000_0000_0000;
array[13454] <= 16'b0000_0000_0000_0000;
array[13455] <= 16'b0000_0000_0000_0000;
array[13456] <= 16'b0000_0000_0000_0000;
array[13457] <= 16'b0000_0000_0000_0000;
array[13458] <= 16'b0000_0000_0000_0000;
array[13459] <= 16'b0000_0000_0000_0000;
array[13460] <= 16'b0000_0000_0000_0000;
array[13461] <= 16'b0000_0000_0000_0000;
array[13462] <= 16'b0000_0000_0000_0000;
array[13463] <= 16'b0000_0000_0000_0000;
array[13464] <= 16'b0000_0000_0000_0000;
array[13465] <= 16'b0000_0000_0000_0000;
array[13466] <= 16'b0000_0000_0000_0000;
array[13467] <= 16'b0000_0000_0000_0000;
array[13468] <= 16'b0000_0000_0000_0000;
array[13469] <= 16'b0000_0000_0000_0000;
array[13470] <= 16'b0000_0000_0000_0000;
array[13471] <= 16'b0000_0000_0000_0000;
array[13472] <= 16'b0000_0000_0000_0000;
array[13473] <= 16'b0000_0000_0000_0000;
array[13474] <= 16'b0000_0000_0000_0000;
array[13475] <= 16'b0000_0000_0000_0000;
array[13476] <= 16'b0000_0000_0000_0000;
array[13477] <= 16'b0000_0000_0000_0000;
array[13478] <= 16'b0000_0000_0000_0000;
array[13479] <= 16'b0000_0000_0000_0000;
array[13480] <= 16'b0000_0000_0000_0000;
array[13481] <= 16'b0000_0000_0000_0000;
array[13482] <= 16'b0000_0000_0000_0000;
array[13483] <= 16'b0000_0000_0000_0000;
array[13484] <= 16'b0000_0000_0000_0000;
array[13485] <= 16'b0000_0000_0000_0000;
array[13486] <= 16'b0000_0000_0000_0000;
array[13487] <= 16'b0000_0000_0000_0000;
array[13488] <= 16'b0000_0000_0000_0000;
array[13489] <= 16'b0000_0000_0000_0000;
array[13490] <= 16'b0000_0000_0000_0000;
array[13491] <= 16'b0000_0000_0000_0000;
array[13492] <= 16'b0000_0000_0000_0000;
array[13493] <= 16'b0000_0000_0000_0000;
array[13494] <= 16'b0000_0000_0000_0000;
array[13495] <= 16'b0000_0000_0000_0000;
array[13496] <= 16'b0000_0000_0000_0000;
array[13497] <= 16'b0000_0000_0000_0000;
array[13498] <= 16'b0000_0000_0000_0000;
array[13499] <= 16'b0000_0000_0000_0000;
array[13500] <= 16'b0000_0000_0000_0000;
array[13501] <= 16'b0000_0000_0000_0000;
array[13502] <= 16'b0000_0000_0000_0000;
array[13503] <= 16'b0000_0000_0000_0000;
array[13504] <= 16'b0000_0000_0000_0000;
array[13505] <= 16'b0000_0000_0000_0000;
array[13506] <= 16'b0000_0000_0000_0000;
array[13507] <= 16'b0000_0000_0000_0000;
array[13508] <= 16'b0000_0000_0000_0000;
array[13509] <= 16'b0000_0000_0000_0000;
array[13510] <= 16'b0000_0000_0000_0000;
array[13511] <= 16'b0000_0000_0000_0000;
array[13512] <= 16'b0000_0000_0000_0000;
array[13513] <= 16'b0000_0000_0000_0000;
array[13514] <= 16'b0000_0000_0000_0000;
array[13515] <= 16'b0000_0000_0000_0000;
array[13516] <= 16'b0000_0000_0000_0000;
array[13517] <= 16'b0000_0000_0000_0000;
array[13518] <= 16'b0000_0000_0000_0000;
array[13519] <= 16'b0000_0000_0000_0000;
array[13520] <= 16'b0000_0000_0000_0000;
array[13521] <= 16'b0000_0000_0000_0000;
array[13522] <= 16'b0000_0000_0000_0000;
array[13523] <= 16'b0000_0000_0000_0000;
array[13524] <= 16'b0000_0000_0000_0000;
array[13525] <= 16'b0000_0000_0000_0000;
array[13526] <= 16'b0000_0000_0000_0000;
array[13527] <= 16'b0000_0000_0000_0000;
array[13528] <= 16'b0000_0000_0000_0000;
array[13529] <= 16'b0000_0000_0000_0000;
array[13530] <= 16'b0000_0000_0000_0000;
array[13531] <= 16'b0000_0000_0000_0000;
array[13532] <= 16'b0000_0000_0000_0000;
array[13533] <= 16'b0000_0000_0000_0000;
array[13534] <= 16'b0000_0000_0000_0000;
array[13535] <= 16'b0000_0000_0000_0000;
array[13536] <= 16'b0000_0000_0000_0000;
array[13537] <= 16'b0000_0000_0000_0000;
array[13538] <= 16'b0000_0000_0000_0000;
array[13539] <= 16'b0000_0000_0000_0000;
array[13540] <= 16'b0000_0000_0000_0000;
array[13541] <= 16'b0000_0000_0000_0000;
array[13542] <= 16'b0000_0000_0000_0000;
array[13543] <= 16'b0000_0000_0000_0000;
array[13544] <= 16'b0000_0000_0000_0000;
array[13545] <= 16'b0000_0000_0000_0000;
array[13546] <= 16'b0000_0000_0000_0000;
array[13547] <= 16'b0000_0000_0000_0000;
array[13548] <= 16'b0000_0000_0000_0000;
array[13549] <= 16'b0000_0000_0000_0000;
array[13550] <= 16'b0000_0000_0000_0000;
array[13551] <= 16'b0000_0000_0000_0000;
array[13552] <= 16'b0000_0000_0000_0000;
array[13553] <= 16'b0000_0000_0000_0000;
array[13554] <= 16'b0000_0000_0000_0000;
array[13555] <= 16'b0000_0000_0000_0000;
array[13556] <= 16'b0000_0000_0000_0000;
array[13557] <= 16'b0000_0000_0000_0000;
array[13558] <= 16'b0000_0000_0000_0000;
array[13559] <= 16'b0000_0000_0000_0000;
array[13560] <= 16'b0000_0000_0000_0000;
array[13561] <= 16'b0000_0000_0000_0000;
array[13562] <= 16'b0000_0000_0000_0000;
array[13563] <= 16'b0000_0000_0000_0000;
array[13564] <= 16'b0000_0000_0000_0000;
array[13565] <= 16'b0000_0000_0000_0000;
array[13566] <= 16'b0000_0000_0000_0000;
array[13567] <= 16'b0000_0000_0000_0000;
array[13568] <= 16'b0000_0000_0000_0000;
array[13569] <= 16'b0000_0000_0000_0000;
array[13570] <= 16'b0000_0000_0000_0000;
array[13571] <= 16'b0000_0000_0000_0000;
array[13572] <= 16'b0000_0000_0000_0000;
array[13573] <= 16'b0000_0000_0000_0000;
array[13574] <= 16'b0000_0000_0000_0000;
array[13575] <= 16'b0000_0000_0000_0000;
array[13576] <= 16'b0000_0000_0000_0000;
array[13577] <= 16'b0000_0000_0000_0000;
array[13578] <= 16'b0000_0000_0000_0000;
array[13579] <= 16'b0000_0000_0000_0000;
array[13580] <= 16'b0000_0000_0000_0000;
array[13581] <= 16'b0000_0000_0000_0000;
array[13582] <= 16'b0000_0000_0000_0000;
array[13583] <= 16'b0000_0000_0000_0000;
array[13584] <= 16'b0000_0000_0000_0000;
array[13585] <= 16'b0000_0000_0000_0000;
array[13586] <= 16'b0000_0000_0000_0000;
array[13587] <= 16'b0000_0000_0000_0000;
array[13588] <= 16'b0000_0000_0000_0000;
array[13589] <= 16'b0000_0000_0000_0000;
array[13590] <= 16'b0000_0000_0000_0000;
array[13591] <= 16'b0000_0000_0000_0000;
array[13592] <= 16'b0000_0000_0000_0000;
array[13593] <= 16'b0000_0000_0000_0000;
array[13594] <= 16'b0000_0000_0000_0000;
array[13595] <= 16'b0000_0000_0000_0000;
array[13596] <= 16'b0000_0000_0000_0000;
array[13597] <= 16'b0000_0000_0000_0000;
array[13598] <= 16'b0000_0000_0000_0000;
array[13599] <= 16'b0000_0000_0000_0000;
array[13600] <= 16'b0000_0000_0000_0000;
array[13601] <= 16'b0000_0000_0000_0000;
array[13602] <= 16'b0000_0000_0000_0000;
array[13603] <= 16'b0000_0000_0000_0000;
array[13604] <= 16'b0000_0000_0000_0000;
array[13605] <= 16'b0000_0000_0000_0000;
array[13606] <= 16'b0000_0000_0000_0000;
array[13607] <= 16'b0000_0000_0000_0000;
array[13608] <= 16'b0000_0000_0000_0000;
array[13609] <= 16'b0000_0000_0000_0000;
array[13610] <= 16'b0000_0000_0000_0000;
array[13611] <= 16'b0000_0000_0000_0000;
array[13612] <= 16'b0000_0000_0000_0000;
array[13613] <= 16'b0000_0000_0000_0000;
array[13614] <= 16'b0000_0000_0000_0000;
array[13615] <= 16'b0000_0000_0000_0000;
array[13616] <= 16'b0000_0000_0000_0000;
array[13617] <= 16'b0000_0000_0000_0000;
array[13618] <= 16'b0000_0000_0000_0000;
array[13619] <= 16'b0000_0000_0000_0000;
array[13620] <= 16'b0000_0000_0000_0000;
array[13621] <= 16'b0000_0000_0000_0000;
array[13622] <= 16'b0000_0000_0000_0000;
array[13623] <= 16'b0000_0000_0000_0000;
array[13624] <= 16'b0000_0000_0000_0000;
array[13625] <= 16'b0000_0000_0000_0000;
array[13626] <= 16'b0000_0000_0000_0000;
array[13627] <= 16'b0000_0000_0000_0000;
array[13628] <= 16'b0000_0000_0000_0000;
array[13629] <= 16'b0000_0000_0000_0000;
array[13630] <= 16'b0000_0000_0000_0000;
array[13631] <= 16'b0000_0000_0000_0000;
array[13632] <= 16'b0000_0000_0000_0000;
array[13633] <= 16'b0000_0000_0000_0000;
array[13634] <= 16'b0000_0000_0000_0000;
array[13635] <= 16'b0000_0000_0000_0000;
array[13636] <= 16'b0000_0000_0000_0000;
array[13637] <= 16'b0000_0000_0000_0000;
array[13638] <= 16'b0000_0000_0000_0000;
array[13639] <= 16'b0000_0000_0000_0000;
array[13640] <= 16'b0000_0000_0000_0000;
array[13641] <= 16'b0000_0000_0000_0000;
array[13642] <= 16'b0000_0000_0000_0000;
array[13643] <= 16'b0000_0000_0000_0000;
array[13644] <= 16'b0000_0000_0000_0000;
array[13645] <= 16'b0000_0000_0000_0000;
array[13646] <= 16'b0000_0000_0000_0000;
array[13647] <= 16'b0000_0000_0000_0000;
array[13648] <= 16'b0000_0000_0000_0000;
array[13649] <= 16'b0000_0000_0000_0000;
array[13650] <= 16'b0000_0000_0000_0000;
array[13651] <= 16'b0000_0000_0000_0000;
array[13652] <= 16'b0000_0000_0000_0000;
array[13653] <= 16'b0000_0000_0000_0000;
array[13654] <= 16'b0000_0000_0000_0000;
array[13655] <= 16'b0000_0000_0000_0000;
array[13656] <= 16'b0000_0000_0000_0000;
array[13657] <= 16'b0000_0000_0000_0000;
array[13658] <= 16'b0000_0000_0000_0000;
array[13659] <= 16'b0000_0000_0000_0000;
array[13660] <= 16'b0000_0000_0000_0000;
array[13661] <= 16'b0000_0000_0000_0000;
array[13662] <= 16'b0000_0000_0000_0000;
array[13663] <= 16'b0000_0000_0000_0000;
array[13664] <= 16'b0000_0000_0000_0000;
array[13665] <= 16'b0000_0000_0000_0000;
array[13666] <= 16'b0000_0000_0000_0000;
array[13667] <= 16'b0000_0000_0000_0000;
array[13668] <= 16'b0000_0000_0000_0000;
array[13669] <= 16'b0000_0000_0000_0000;
array[13670] <= 16'b0000_0000_0000_0000;
array[13671] <= 16'b0000_0000_0000_0000;
array[13672] <= 16'b0000_0000_0000_0000;
array[13673] <= 16'b0000_0000_0000_0000;
array[13674] <= 16'b0000_0000_0000_0000;
array[13675] <= 16'b0000_0000_0000_0000;
array[13676] <= 16'b0000_0000_0000_0000;
array[13677] <= 16'b0000_0000_0000_0000;
array[13678] <= 16'b0000_0000_0000_0000;
array[13679] <= 16'b0000_0000_0000_0000;
array[13680] <= 16'b0000_0000_0000_0000;
array[13681] <= 16'b0000_0000_0000_0000;
array[13682] <= 16'b0000_0000_0000_0000;
array[13683] <= 16'b0000_0000_0000_0000;
array[13684] <= 16'b0000_0000_0000_0000;
array[13685] <= 16'b0000_0000_0000_0000;
array[13686] <= 16'b0000_0000_0000_0000;
array[13687] <= 16'b0000_0000_0000_0000;
array[13688] <= 16'b0000_0000_0000_0000;
array[13689] <= 16'b0000_0000_0000_0000;
array[13690] <= 16'b0000_0000_0000_0000;
array[13691] <= 16'b0000_0000_0000_0000;
array[13692] <= 16'b0000_0000_0000_0000;
array[13693] <= 16'b0000_0000_0000_0000;
array[13694] <= 16'b0000_0000_0000_0000;
array[13695] <= 16'b0000_0000_0000_0000;
array[13696] <= 16'b0000_0000_0000_0000;
array[13697] <= 16'b0000_0000_0000_0000;
array[13698] <= 16'b0000_0000_0000_0000;
array[13699] <= 16'b0000_0000_0000_0000;
array[13700] <= 16'b0000_0000_0000_0000;
array[13701] <= 16'b0000_0000_0000_0000;
array[13702] <= 16'b0000_0000_0000_0000;
array[13703] <= 16'b0000_0000_0000_0000;
array[13704] <= 16'b0000_0000_0000_0000;
array[13705] <= 16'b0000_0000_0000_0000;
array[13706] <= 16'b0000_0000_0000_0000;
array[13707] <= 16'b0000_0000_0000_0000;
array[13708] <= 16'b0000_0000_0000_0000;
array[13709] <= 16'b0000_0000_0000_0000;
array[13710] <= 16'b0000_0000_0000_0000;
array[13711] <= 16'b0000_0000_0000_0000;
array[13712] <= 16'b0000_0000_0000_0000;
array[13713] <= 16'b0000_0000_0000_0000;
array[13714] <= 16'b0000_0000_0000_0000;
array[13715] <= 16'b0000_0000_0000_0000;
array[13716] <= 16'b0000_0000_0000_0000;
array[13717] <= 16'b0000_0000_0000_0000;
array[13718] <= 16'b0000_0000_0000_0000;
array[13719] <= 16'b0000_0000_0000_0000;
array[13720] <= 16'b0000_0000_0000_0000;
array[13721] <= 16'b0000_0000_0000_0000;
array[13722] <= 16'b0000_0000_0000_0000;
array[13723] <= 16'b0000_0000_0000_0000;
array[13724] <= 16'b0000_0000_0000_0000;
array[13725] <= 16'b0000_0000_0000_0000;
array[13726] <= 16'b0000_0000_0000_0000;
array[13727] <= 16'b0000_0000_0000_0000;
array[13728] <= 16'b0000_0000_0000_0000;
array[13729] <= 16'b0000_0000_0000_0000;
array[13730] <= 16'b0000_0000_0000_0000;
array[13731] <= 16'b0000_0000_0000_0000;
array[13732] <= 16'b0000_0000_0000_0000;
array[13733] <= 16'b0000_0000_0000_0000;
array[13734] <= 16'b0000_0000_0000_0000;
array[13735] <= 16'b0000_0000_0000_0000;
array[13736] <= 16'b0000_0000_0000_0000;
array[13737] <= 16'b0000_0000_0000_0000;
array[13738] <= 16'b0000_0000_0000_0000;
array[13739] <= 16'b0000_0000_0000_0000;
array[13740] <= 16'b0000_0000_0000_0000;
array[13741] <= 16'b0000_0000_0000_0000;
array[13742] <= 16'b0000_0000_0000_0000;
array[13743] <= 16'b0000_0000_0000_0000;
array[13744] <= 16'b0000_0000_0000_0000;
array[13745] <= 16'b0000_0000_0000_0000;
array[13746] <= 16'b0000_0000_0000_0000;
array[13747] <= 16'b0000_0000_0000_0000;
array[13748] <= 16'b0000_0000_0000_0000;
array[13749] <= 16'b0000_0000_0000_0000;
array[13750] <= 16'b0000_0000_0000_0000;
array[13751] <= 16'b0000_0000_0000_0000;
array[13752] <= 16'b0000_0000_0000_0000;
array[13753] <= 16'b0000_0000_0000_0000;
array[13754] <= 16'b0000_0000_0000_0000;
array[13755] <= 16'b0000_0000_0000_0000;
array[13756] <= 16'b0000_0000_0000_0000;
array[13757] <= 16'b0000_0000_0000_0000;
array[13758] <= 16'b0000_0000_0000_0000;
array[13759] <= 16'b0000_0000_0000_0000;
array[13760] <= 16'b0000_0000_0000_0000;
array[13761] <= 16'b0000_0000_0000_0000;
array[13762] <= 16'b0000_0000_0000_0000;
array[13763] <= 16'b0000_0000_0000_0000;
array[13764] <= 16'b0000_0000_0000_0000;
array[13765] <= 16'b0000_0000_0000_0000;
array[13766] <= 16'b0000_0000_0000_0000;
array[13767] <= 16'b0000_0000_0000_0000;
array[13768] <= 16'b0000_0000_0000_0000;
array[13769] <= 16'b0000_0000_0000_0000;
array[13770] <= 16'b0000_0000_0000_0000;
array[13771] <= 16'b0000_0000_0000_0000;
array[13772] <= 16'b0000_0000_0000_0000;
array[13773] <= 16'b0000_0000_0000_0000;
array[13774] <= 16'b0000_0000_0000_0000;
array[13775] <= 16'b0000_0000_0000_0000;
array[13776] <= 16'b0000_0000_0000_0000;
array[13777] <= 16'b0000_0000_0000_0000;
array[13778] <= 16'b0000_0000_0000_0000;
array[13779] <= 16'b0000_0000_0000_0000;
array[13780] <= 16'b0000_0000_0000_0000;
array[13781] <= 16'b0000_0000_0000_0000;
array[13782] <= 16'b0000_0000_0000_0000;
array[13783] <= 16'b0000_0000_0000_0000;
array[13784] <= 16'b0000_0000_0000_0000;
array[13785] <= 16'b0000_0000_0000_0000;
array[13786] <= 16'b0000_0000_0000_0000;
array[13787] <= 16'b0000_0000_0000_0000;
array[13788] <= 16'b0000_0000_0000_0000;
array[13789] <= 16'b0000_0000_0000_0000;
array[13790] <= 16'b0000_0000_0000_0000;
array[13791] <= 16'b0000_0000_0000_0000;
array[13792] <= 16'b0000_0000_0000_0000;
array[13793] <= 16'b0000_0000_0000_0000;
array[13794] <= 16'b0000_0000_0000_0000;
array[13795] <= 16'b0000_0000_0000_0000;
array[13796] <= 16'b0000_0000_0000_0000;
array[13797] <= 16'b0000_0000_0000_0000;
array[13798] <= 16'b0000_0000_0000_0000;
array[13799] <= 16'b0000_0000_0000_0000;
array[13800] <= 16'b0000_0000_0000_0000;
array[13801] <= 16'b0000_0000_0000_0000;
array[13802] <= 16'b0000_0000_0000_0000;
array[13803] <= 16'b0000_0000_0000_0000;
array[13804] <= 16'b0000_0000_0000_0000;
array[13805] <= 16'b0000_0000_0000_0000;
array[13806] <= 16'b0000_0000_0000_0000;
array[13807] <= 16'b0000_0000_0000_0000;
array[13808] <= 16'b0000_0000_0000_0000;
array[13809] <= 16'b0000_0000_0000_0000;
array[13810] <= 16'b0000_0000_0000_0000;
array[13811] <= 16'b0000_0000_0000_0000;
array[13812] <= 16'b0000_0000_0000_0000;
array[13813] <= 16'b0000_0000_0000_0000;
array[13814] <= 16'b0000_0000_0000_0000;
array[13815] <= 16'b0000_0000_0000_0000;
array[13816] <= 16'b0000_0000_0000_0000;
array[13817] <= 16'b0000_0000_0000_0000;
array[13818] <= 16'b0000_0000_0000_0000;
array[13819] <= 16'b0000_0000_0000_0000;
array[13820] <= 16'b0000_0000_0000_0000;
array[13821] <= 16'b0000_0000_0000_0000;
array[13822] <= 16'b0000_0000_0000_0000;
array[13823] <= 16'b0000_0000_0000_0000;
array[13824] <= 16'b0000_0000_0000_0000;
array[13825] <= 16'b0000_0000_0000_0000;
array[13826] <= 16'b0000_0000_0000_0000;
array[13827] <= 16'b0000_0000_0000_0000;
array[13828] <= 16'b0000_0000_0000_0000;
array[13829] <= 16'b0000_0000_0000_0000;
array[13830] <= 16'b0000_0000_0000_0000;
array[13831] <= 16'b0000_0000_0000_0000;
array[13832] <= 16'b0000_0000_0000_0000;
array[13833] <= 16'b0000_0000_0000_0000;
array[13834] <= 16'b0000_0000_0000_0000;
array[13835] <= 16'b0000_0000_0000_0000;
array[13836] <= 16'b0000_0000_0000_0000;
array[13837] <= 16'b0000_0000_0000_0000;
array[13838] <= 16'b0000_0000_0000_0000;
array[13839] <= 16'b0000_0000_0000_0000;
array[13840] <= 16'b0000_0000_0000_0000;
array[13841] <= 16'b0000_0000_0000_0000;
array[13842] <= 16'b0000_0000_0000_0000;
array[13843] <= 16'b0000_0000_0000_0000;
array[13844] <= 16'b0000_0000_0000_0000;
array[13845] <= 16'b0000_0000_0000_0000;
array[13846] <= 16'b0000_0000_0000_0000;
array[13847] <= 16'b0000_0000_0000_0000;
array[13848] <= 16'b0000_0000_0000_0000;
array[13849] <= 16'b0000_0000_0000_0000;
array[13850] <= 16'b0000_0000_0000_0000;
array[13851] <= 16'b0000_0000_0000_0000;
array[13852] <= 16'b0000_0000_0000_0000;
array[13853] <= 16'b0000_0000_0000_0000;
array[13854] <= 16'b0000_0000_0000_0000;
array[13855] <= 16'b0000_0000_0000_0000;
array[13856] <= 16'b0000_0000_0000_0000;
array[13857] <= 16'b0000_0000_0000_0000;
array[13858] <= 16'b0000_0000_0000_0000;
array[13859] <= 16'b0000_0000_0000_0000;
array[13860] <= 16'b0000_0000_0000_0000;
array[13861] <= 16'b0000_0000_0000_0000;
array[13862] <= 16'b0000_0000_0000_0000;
array[13863] <= 16'b0000_0000_0000_0000;
array[13864] <= 16'b0000_0000_0000_0000;
array[13865] <= 16'b0000_0000_0000_0000;
array[13866] <= 16'b0000_0000_0000_0000;
array[13867] <= 16'b0000_0000_0000_0000;
array[13868] <= 16'b0000_0000_0000_0000;
array[13869] <= 16'b0000_0000_0000_0000;
array[13870] <= 16'b0000_0000_0000_0000;
array[13871] <= 16'b0000_0000_0000_0000;
array[13872] <= 16'b0000_0000_0000_0000;
array[13873] <= 16'b0000_0000_0000_0000;
array[13874] <= 16'b0000_0000_0000_0000;
array[13875] <= 16'b0000_0000_0000_0000;
array[13876] <= 16'b0000_0000_0000_0000;
array[13877] <= 16'b0000_0000_0000_0000;
array[13878] <= 16'b0000_0000_0000_0000;
array[13879] <= 16'b0000_0000_0000_0000;
array[13880] <= 16'b0000_0000_0000_0000;
array[13881] <= 16'b0000_0000_0000_0000;
array[13882] <= 16'b0000_0000_0000_0000;
array[13883] <= 16'b0000_0000_0000_0000;
array[13884] <= 16'b0000_0000_0000_0000;
array[13885] <= 16'b0000_0000_0000_0000;
array[13886] <= 16'b0000_0000_0000_0000;
array[13887] <= 16'b0000_0000_0000_0000;
array[13888] <= 16'b0000_0000_0000_0000;
array[13889] <= 16'b0000_0000_0000_0000;
array[13890] <= 16'b0000_0000_0000_0000;
array[13891] <= 16'b0000_0000_0000_0000;
array[13892] <= 16'b0000_0000_0000_0000;
array[13893] <= 16'b0000_0000_0000_0000;
array[13894] <= 16'b0000_0000_0000_0000;
array[13895] <= 16'b0000_0000_0000_0000;
array[13896] <= 16'b0000_0000_0000_0000;
array[13897] <= 16'b0000_0000_0000_0000;
array[13898] <= 16'b0000_0000_0000_0000;
array[13899] <= 16'b0000_0000_0000_0000;
array[13900] <= 16'b0000_0000_0000_0000;
array[13901] <= 16'b0000_0000_0000_0000;
array[13902] <= 16'b0000_0000_0000_0000;
array[13903] <= 16'b0000_0000_0000_0000;
array[13904] <= 16'b0000_0000_0000_0000;
array[13905] <= 16'b0000_0000_0000_0000;
array[13906] <= 16'b0000_0000_0000_0000;
array[13907] <= 16'b0000_0000_0000_0000;
array[13908] <= 16'b0000_0000_0000_0000;
array[13909] <= 16'b0000_0000_0000_0000;
array[13910] <= 16'b0000_0000_0000_0000;
array[13911] <= 16'b0000_0000_0000_0000;
array[13912] <= 16'b0000_0000_0000_0000;
array[13913] <= 16'b0000_0000_0000_0000;
array[13914] <= 16'b0000_0000_0000_0000;
array[13915] <= 16'b0000_0000_0000_0000;
array[13916] <= 16'b0000_0000_0000_0000;
array[13917] <= 16'b0000_0000_0000_0000;
array[13918] <= 16'b0000_0000_0000_0000;
array[13919] <= 16'b0000_0000_0000_0000;
array[13920] <= 16'b0000_0000_0000_0000;
array[13921] <= 16'b0000_0000_0000_0000;
array[13922] <= 16'b0000_0000_0000_0000;
array[13923] <= 16'b0000_0000_0000_0000;
array[13924] <= 16'b0000_0000_0000_0000;
array[13925] <= 16'b0000_0000_0000_0000;
array[13926] <= 16'b0000_0000_0000_0000;
array[13927] <= 16'b0000_0000_0000_0000;
array[13928] <= 16'b0000_0000_0000_0000;
array[13929] <= 16'b0000_0000_0000_0000;
array[13930] <= 16'b0000_0000_0000_0000;
array[13931] <= 16'b0000_0000_0000_0000;
array[13932] <= 16'b0000_0000_0000_0000;
array[13933] <= 16'b0000_0000_0000_0000;
array[13934] <= 16'b0000_0000_0000_0000;
array[13935] <= 16'b0000_0000_0000_0000;
array[13936] <= 16'b0000_0000_0000_0000;
array[13937] <= 16'b0000_0000_0000_0000;
array[13938] <= 16'b0000_0000_0000_0000;
array[13939] <= 16'b0000_0000_0000_0000;
array[13940] <= 16'b0000_0000_0000_0000;
array[13941] <= 16'b0000_0000_0000_0000;
array[13942] <= 16'b0000_0000_0000_0000;
array[13943] <= 16'b0000_0000_0000_0000;
array[13944] <= 16'b0000_0000_0000_0000;
array[13945] <= 16'b0000_0000_0000_0000;
array[13946] <= 16'b0000_0000_0000_0000;
array[13947] <= 16'b0000_0000_0000_0000;
array[13948] <= 16'b0000_0000_0000_0000;
array[13949] <= 16'b0000_0000_0000_0000;
array[13950] <= 16'b0000_0000_0000_0000;
array[13951] <= 16'b0000_0000_0000_0000;
array[13952] <= 16'b0000_0000_0000_0000;
array[13953] <= 16'b0000_0000_0000_0000;
array[13954] <= 16'b0000_0000_0000_0000;
array[13955] <= 16'b0000_0000_0000_0000;
array[13956] <= 16'b0000_0000_0000_0000;
array[13957] <= 16'b0000_0000_0000_0000;
array[13958] <= 16'b0000_0000_0000_0000;
array[13959] <= 16'b0000_0000_0000_0000;
array[13960] <= 16'b0000_0000_0000_0000;
array[13961] <= 16'b0000_0000_0000_0000;
array[13962] <= 16'b0000_0000_0000_0000;
array[13963] <= 16'b0000_0000_0000_0000;
array[13964] <= 16'b0000_0000_0000_0000;
array[13965] <= 16'b0000_0000_0000_0000;
array[13966] <= 16'b0000_0000_0000_0000;
array[13967] <= 16'b0000_0000_0000_0000;
array[13968] <= 16'b0000_0000_0000_0000;
array[13969] <= 16'b0000_0000_0000_0000;
array[13970] <= 16'b0000_0000_0000_0000;
array[13971] <= 16'b0000_0000_0000_0000;
array[13972] <= 16'b0000_0000_0000_0000;
array[13973] <= 16'b0000_0000_0000_0000;
array[13974] <= 16'b0000_0000_0000_0000;
array[13975] <= 16'b0000_0000_0000_0000;
array[13976] <= 16'b0000_0000_0000_0000;
array[13977] <= 16'b0000_0000_0000_0000;
array[13978] <= 16'b0000_0000_0000_0000;
array[13979] <= 16'b0000_0000_0000_0000;
array[13980] <= 16'b0000_0000_0000_0000;
array[13981] <= 16'b0000_0000_0000_0000;
array[13982] <= 16'b0000_0000_0000_0000;
array[13983] <= 16'b0000_0000_0000_0000;
array[13984] <= 16'b0000_0000_0000_0000;
array[13985] <= 16'b0000_0000_0000_0000;
array[13986] <= 16'b0000_0000_0000_0000;
array[13987] <= 16'b0000_0000_0000_0000;
array[13988] <= 16'b0000_0000_0000_0000;
array[13989] <= 16'b0000_0000_0000_0000;
array[13990] <= 16'b0000_0000_0000_0000;
array[13991] <= 16'b0000_0000_0000_0000;
array[13992] <= 16'b0000_0000_0000_0000;
array[13993] <= 16'b0000_0000_0000_0000;
array[13994] <= 16'b0000_0000_0000_0000;
array[13995] <= 16'b0000_0000_0000_0000;
array[13996] <= 16'b0000_0000_0000_0000;
array[13997] <= 16'b0000_0000_0000_0000;
array[13998] <= 16'b0000_0000_0000_0000;
array[13999] <= 16'b0000_0000_0000_0000;
array[14000] <= 16'b0000_0000_0000_0000;
array[14001] <= 16'b0000_0000_0000_0000;
array[14002] <= 16'b0000_0000_0000_0000;
array[14003] <= 16'b0000_0000_0000_0000;
array[14004] <= 16'b0000_0000_0000_0000;
array[14005] <= 16'b0000_0000_0000_0000;
array[14006] <= 16'b0000_0000_0000_0000;
array[14007] <= 16'b0000_0000_0000_0000;
array[14008] <= 16'b0000_0000_0000_0000;
array[14009] <= 16'b0000_0000_0000_0000;
array[14010] <= 16'b0000_0000_0000_0000;
array[14011] <= 16'b0000_0000_0000_0000;
array[14012] <= 16'b0000_0000_0000_0000;
array[14013] <= 16'b0000_0000_0000_0000;
array[14014] <= 16'b0000_0000_0000_0000;
array[14015] <= 16'b0000_0000_0000_0000;
array[14016] <= 16'b0000_0000_0000_0000;
array[14017] <= 16'b0000_0000_0000_0000;
array[14018] <= 16'b0000_0000_0000_0000;
array[14019] <= 16'b0000_0000_0000_0000;
array[14020] <= 16'b0000_0000_0000_0000;
array[14021] <= 16'b0000_0000_0000_0000;
array[14022] <= 16'b0000_0000_0000_0000;
array[14023] <= 16'b0000_0000_0000_0000;
array[14024] <= 16'b0000_0000_0000_0000;
array[14025] <= 16'b0000_0000_0000_0000;
array[14026] <= 16'b0000_0000_0000_0000;
array[14027] <= 16'b0000_0000_0000_0000;
array[14028] <= 16'b0000_0000_0000_0000;
array[14029] <= 16'b0000_0000_0000_0000;
array[14030] <= 16'b0000_0000_0000_0000;
array[14031] <= 16'b0000_0000_0000_0000;
array[14032] <= 16'b0000_0000_0000_0000;
array[14033] <= 16'b0000_0000_0000_0000;
array[14034] <= 16'b0000_0000_0000_0000;
array[14035] <= 16'b0000_0000_0000_0000;
array[14036] <= 16'b0000_0000_0000_0000;
array[14037] <= 16'b0000_0000_0000_0000;
array[14038] <= 16'b0000_0000_0000_0000;
array[14039] <= 16'b0000_0000_0000_0000;
array[14040] <= 16'b0000_0000_0000_0000;
array[14041] <= 16'b0000_0000_0000_0000;
array[14042] <= 16'b0000_0000_0000_0000;
array[14043] <= 16'b0000_0000_0000_0000;
array[14044] <= 16'b0000_0000_0000_0000;
array[14045] <= 16'b0000_0000_0000_0000;
array[14046] <= 16'b0000_0000_0000_0000;
array[14047] <= 16'b0000_0000_0000_0000;
array[14048] <= 16'b0000_0000_0000_0000;
array[14049] <= 16'b0000_0000_0000_0000;
array[14050] <= 16'b0000_0000_0000_0000;
array[14051] <= 16'b0000_0000_0000_0000;
array[14052] <= 16'b0000_0000_0000_0000;
array[14053] <= 16'b0000_0000_0000_0000;
array[14054] <= 16'b0000_0000_0000_0000;
array[14055] <= 16'b0000_0000_0000_0000;
array[14056] <= 16'b0000_0000_0000_0000;
array[14057] <= 16'b0000_0000_0000_0000;
array[14058] <= 16'b0000_0000_0000_0000;
array[14059] <= 16'b0000_0000_0000_0000;
array[14060] <= 16'b0000_0000_0000_0000;
array[14061] <= 16'b0000_0000_0000_0000;
array[14062] <= 16'b0000_0000_0000_0000;
array[14063] <= 16'b0000_0000_0000_0000;
array[14064] <= 16'b0000_0000_0000_0000;
array[14065] <= 16'b0000_0000_0000_0000;
array[14066] <= 16'b0000_0000_0000_0000;
array[14067] <= 16'b0000_0000_0000_0000;
array[14068] <= 16'b0000_0000_0000_0000;
array[14069] <= 16'b0000_0000_0000_0000;
array[14070] <= 16'b0000_0000_0000_0000;
array[14071] <= 16'b0000_0000_0000_0000;
array[14072] <= 16'b0000_0000_0000_0000;
array[14073] <= 16'b0000_0000_0000_0000;
array[14074] <= 16'b0000_0000_0000_0000;
array[14075] <= 16'b0000_0000_0000_0000;
array[14076] <= 16'b0000_0000_0000_0000;
array[14077] <= 16'b0000_0000_0000_0000;
array[14078] <= 16'b0000_0000_0000_0000;
array[14079] <= 16'b0000_0000_0000_0000;
array[14080] <= 16'b0000_0000_0000_0000;
array[14081] <= 16'b0000_0000_0000_0000;
array[14082] <= 16'b0000_0000_0000_0000;
array[14083] <= 16'b0000_0000_0000_0000;
array[14084] <= 16'b0000_0000_0000_0000;
array[14085] <= 16'b0000_0000_0000_0000;
array[14086] <= 16'b0000_0000_0000_0000;
array[14087] <= 16'b0000_0000_0000_0000;
array[14088] <= 16'b0000_0000_0000_0000;
array[14089] <= 16'b0000_0000_0000_0000;
array[14090] <= 16'b0000_0000_0000_0000;
array[14091] <= 16'b0000_0000_0000_0000;
array[14092] <= 16'b0000_0000_0000_0000;
array[14093] <= 16'b0000_0000_0000_0000;
array[14094] <= 16'b0000_0000_0000_0000;
array[14095] <= 16'b0000_0000_0000_0000;
array[14096] <= 16'b0000_0000_0000_0000;
array[14097] <= 16'b0000_0000_0000_0000;
array[14098] <= 16'b0000_0000_0000_0000;
array[14099] <= 16'b0000_0000_0000_0000;
array[14100] <= 16'b0000_0000_0000_0000;
array[14101] <= 16'b0000_0000_0000_0000;
array[14102] <= 16'b0000_0000_0000_0000;
array[14103] <= 16'b0000_0000_0000_0000;
array[14104] <= 16'b0000_0000_0000_0000;
array[14105] <= 16'b0000_0000_0000_0000;
array[14106] <= 16'b0000_0000_0000_0000;
array[14107] <= 16'b0000_0000_0000_0000;
array[14108] <= 16'b0000_0000_0000_0000;
array[14109] <= 16'b0000_0000_0000_0000;
array[14110] <= 16'b0000_0000_0000_0000;
array[14111] <= 16'b0000_0000_0000_0000;
array[14112] <= 16'b0000_0000_0000_0000;
array[14113] <= 16'b0000_0000_0000_0000;
array[14114] <= 16'b0000_0000_0000_0000;
array[14115] <= 16'b0000_0000_0000_0000;
array[14116] <= 16'b0000_0000_0000_0000;
array[14117] <= 16'b0000_0000_0000_0000;
array[14118] <= 16'b0000_0000_0000_0000;
array[14119] <= 16'b0000_0000_0000_0000;
array[14120] <= 16'b0000_0000_0000_0000;
array[14121] <= 16'b0000_0000_0000_0000;
array[14122] <= 16'b0000_0000_0000_0000;
array[14123] <= 16'b0000_0000_0000_0000;
array[14124] <= 16'b0000_0000_0000_0000;
array[14125] <= 16'b0000_0000_0000_0000;
array[14126] <= 16'b0000_0000_0000_0000;
array[14127] <= 16'b0000_0000_0000_0000;
array[14128] <= 16'b0000_0000_0000_0000;
array[14129] <= 16'b0000_0000_0000_0000;
array[14130] <= 16'b0000_0000_0000_0000;
array[14131] <= 16'b0000_0000_0000_0000;
array[14132] <= 16'b0000_0000_0000_0000;
array[14133] <= 16'b0000_0000_0000_0000;
array[14134] <= 16'b0000_0000_0000_0000;
array[14135] <= 16'b0000_0000_0000_0000;
array[14136] <= 16'b0000_0000_0000_0000;
array[14137] <= 16'b0000_0000_0000_0000;
array[14138] <= 16'b0000_0000_0000_0000;
array[14139] <= 16'b0000_0000_0000_0000;
array[14140] <= 16'b0000_0000_0000_0000;
array[14141] <= 16'b0000_0000_0000_0000;
array[14142] <= 16'b0000_0000_0000_0000;
array[14143] <= 16'b0000_0000_0000_0000;
array[14144] <= 16'b0000_0000_0000_0000;
array[14145] <= 16'b0000_0000_0000_0000;
array[14146] <= 16'b0000_0000_0000_0000;
array[14147] <= 16'b0000_0000_0000_0000;
array[14148] <= 16'b0000_0000_0000_0000;
array[14149] <= 16'b0000_0000_0000_0000;
array[14150] <= 16'b0000_0000_0000_0000;
array[14151] <= 16'b0000_0000_0000_0000;
array[14152] <= 16'b0000_0000_0000_0000;
array[14153] <= 16'b0000_0000_0000_0000;
array[14154] <= 16'b0000_0000_0000_0000;
array[14155] <= 16'b0000_0000_0000_0000;
array[14156] <= 16'b0000_0000_0000_0000;
array[14157] <= 16'b0000_0000_0000_0000;
array[14158] <= 16'b0000_0000_0000_0000;
array[14159] <= 16'b0000_0000_0000_0000;
array[14160] <= 16'b0000_0000_0000_0000;
array[14161] <= 16'b0000_0000_0000_0000;
array[14162] <= 16'b0000_0000_0000_0000;
array[14163] <= 16'b0000_0000_0000_0000;
array[14164] <= 16'b0000_0000_0000_0000;
array[14165] <= 16'b0000_0000_0000_0000;
array[14166] <= 16'b0000_0000_0000_0000;
array[14167] <= 16'b0000_0000_0000_0000;
array[14168] <= 16'b0000_0000_0000_0000;
array[14169] <= 16'b0000_0000_0000_0000;
array[14170] <= 16'b0000_0000_0000_0000;
array[14171] <= 16'b0000_0000_0000_0000;
array[14172] <= 16'b0000_0000_0000_0000;
array[14173] <= 16'b0000_0000_0000_0000;
array[14174] <= 16'b0000_0000_0000_0000;
array[14175] <= 16'b0000_0000_0000_0000;
array[14176] <= 16'b0000_0000_0000_0000;
array[14177] <= 16'b0000_0000_0000_0000;
array[14178] <= 16'b0000_0000_0000_0000;
array[14179] <= 16'b0000_0000_0000_0000;
array[14180] <= 16'b0000_0000_0000_0000;
array[14181] <= 16'b0000_0000_0000_0000;
array[14182] <= 16'b0000_0000_0000_0000;
array[14183] <= 16'b0000_0000_0000_0000;
array[14184] <= 16'b0000_0000_0000_0000;
array[14185] <= 16'b0000_0000_0000_0000;
array[14186] <= 16'b0000_0000_0000_0000;
array[14187] <= 16'b0000_0000_0000_0000;
array[14188] <= 16'b0000_0000_0000_0000;
array[14189] <= 16'b0000_0000_0000_0000;
array[14190] <= 16'b0000_0000_0000_0000;
array[14191] <= 16'b0000_0000_0000_0000;
array[14192] <= 16'b0000_0000_0000_0000;
array[14193] <= 16'b0000_0000_0000_0000;
array[14194] <= 16'b0000_0000_0000_0000;
array[14195] <= 16'b0000_0000_0000_0000;
array[14196] <= 16'b0000_0000_0000_0000;
array[14197] <= 16'b0000_0000_0000_0000;
array[14198] <= 16'b0000_0000_0000_0000;
array[14199] <= 16'b0000_0000_0000_0000;
array[14200] <= 16'b0000_0000_0000_0000;
array[14201] <= 16'b0000_0000_0000_0000;
array[14202] <= 16'b0000_0000_0000_0000;
array[14203] <= 16'b0000_0000_0000_0000;
array[14204] <= 16'b0000_0000_0000_0000;
array[14205] <= 16'b0000_0000_0000_0000;
array[14206] <= 16'b0000_0000_0000_0000;
array[14207] <= 16'b0000_0000_0000_0000;
array[14208] <= 16'b0000_0000_0000_0000;
array[14209] <= 16'b0000_0000_0000_0000;
array[14210] <= 16'b0000_0000_0000_0000;
array[14211] <= 16'b0000_0000_0000_0000;
array[14212] <= 16'b0000_0000_0000_0000;
array[14213] <= 16'b0000_0000_0000_0000;
array[14214] <= 16'b0000_0000_0000_0000;
array[14215] <= 16'b0000_0000_0000_0000;
array[14216] <= 16'b0000_0000_0000_0000;
array[14217] <= 16'b0000_0000_0000_0000;
array[14218] <= 16'b0000_0000_0000_0000;
array[14219] <= 16'b0000_0000_0000_0000;
array[14220] <= 16'b0000_0000_0000_0000;
array[14221] <= 16'b0000_0000_0000_0000;
array[14222] <= 16'b0000_0000_0000_0000;
array[14223] <= 16'b0000_0000_0000_0000;
array[14224] <= 16'b0000_0000_0000_0000;
array[14225] <= 16'b0000_0000_0000_0000;
array[14226] <= 16'b0000_0000_0000_0000;
array[14227] <= 16'b0000_0000_0000_0000;
array[14228] <= 16'b0000_0000_0000_0000;
array[14229] <= 16'b0000_0000_0000_0000;
array[14230] <= 16'b0000_0000_0000_0000;
array[14231] <= 16'b0000_0000_0000_0000;
array[14232] <= 16'b0000_0000_0000_0000;
array[14233] <= 16'b0000_0000_0000_0000;
array[14234] <= 16'b0000_0000_0000_0000;
array[14235] <= 16'b0000_0000_0000_0000;
array[14236] <= 16'b0000_0000_0000_0000;
array[14237] <= 16'b0000_0000_0000_0000;
array[14238] <= 16'b0000_0000_0000_0000;
array[14239] <= 16'b0000_0000_0000_0000;
array[14240] <= 16'b0000_0000_0000_0000;
array[14241] <= 16'b0000_0000_0000_0000;
array[14242] <= 16'b0000_0000_0000_0000;
array[14243] <= 16'b0000_0000_0000_0000;
array[14244] <= 16'b0000_0000_0000_0000;
array[14245] <= 16'b0000_0000_0000_0000;
array[14246] <= 16'b0000_0000_0000_0000;
array[14247] <= 16'b0000_0000_0000_0000;
array[14248] <= 16'b0000_0000_0000_0000;
array[14249] <= 16'b0000_0000_0000_0000;
array[14250] <= 16'b0000_0000_0000_0000;
array[14251] <= 16'b0000_0000_0000_0000;
array[14252] <= 16'b0000_0000_0000_0000;
array[14253] <= 16'b0000_0000_0000_0000;
array[14254] <= 16'b0000_0000_0000_0000;
array[14255] <= 16'b0000_0000_0000_0000;
array[14256] <= 16'b0000_0000_0000_0000;
array[14257] <= 16'b0000_0000_0000_0000;
array[14258] <= 16'b0000_0000_0000_0000;
array[14259] <= 16'b0000_0000_0000_0000;
array[14260] <= 16'b0000_0000_0000_0000;
array[14261] <= 16'b0000_0000_0000_0000;
array[14262] <= 16'b0000_0000_0000_0000;
array[14263] <= 16'b0000_0000_0000_0000;
array[14264] <= 16'b0000_0000_0000_0000;
array[14265] <= 16'b0000_0000_0000_0000;
array[14266] <= 16'b0000_0000_0000_0000;
array[14267] <= 16'b0000_0000_0000_0000;
array[14268] <= 16'b0000_0000_0000_0000;
array[14269] <= 16'b0000_0000_0000_0000;
array[14270] <= 16'b0000_0000_0000_0000;
array[14271] <= 16'b0000_0000_0000_0000;
array[14272] <= 16'b0000_0000_0000_0000;
array[14273] <= 16'b0000_0000_0000_0000;
array[14274] <= 16'b0000_0000_0000_0000;
array[14275] <= 16'b0000_0000_0000_0000;
array[14276] <= 16'b0000_0000_0000_0000;
array[14277] <= 16'b0000_0000_0000_0000;
array[14278] <= 16'b0000_0000_0000_0000;
array[14279] <= 16'b0000_0000_0000_0000;
array[14280] <= 16'b0000_0000_0000_0000;
array[14281] <= 16'b0000_0000_0000_0000;
array[14282] <= 16'b0000_0000_0000_0000;
array[14283] <= 16'b0000_0000_0000_0000;
array[14284] <= 16'b0000_0000_0000_0000;
array[14285] <= 16'b0000_0000_0000_0000;
array[14286] <= 16'b0000_0000_0000_0000;
array[14287] <= 16'b0000_0000_0000_0000;
array[14288] <= 16'b0000_0000_0000_0000;
array[14289] <= 16'b0000_0000_0000_0000;
array[14290] <= 16'b0000_0000_0000_0000;
array[14291] <= 16'b0000_0000_0000_0000;
array[14292] <= 16'b0000_0000_0000_0000;
array[14293] <= 16'b0000_0000_0000_0000;
array[14294] <= 16'b0000_0000_0000_0000;
array[14295] <= 16'b0000_0000_0000_0000;
array[14296] <= 16'b0000_0000_0000_0000;
array[14297] <= 16'b0000_0000_0000_0000;
array[14298] <= 16'b0000_0000_0000_0000;
array[14299] <= 16'b0000_0000_0000_0000;
array[14300] <= 16'b0000_0000_0000_0000;
array[14301] <= 16'b0000_0000_0000_0000;
array[14302] <= 16'b0000_0000_0000_0000;
array[14303] <= 16'b0000_0000_0000_0000;
array[14304] <= 16'b0000_0000_0000_0000;
array[14305] <= 16'b0000_0000_0000_0000;
array[14306] <= 16'b0000_0000_0000_0000;
array[14307] <= 16'b0000_0000_0000_0000;
array[14308] <= 16'b0000_0000_0000_0000;
array[14309] <= 16'b0000_0000_0000_0000;
array[14310] <= 16'b0000_0000_0000_0000;
array[14311] <= 16'b0000_0000_0000_0000;
array[14312] <= 16'b0000_0000_0000_0000;
array[14313] <= 16'b0000_0000_0000_0000;
array[14314] <= 16'b0000_0000_0000_0000;
array[14315] <= 16'b0000_0000_0000_0000;
array[14316] <= 16'b0000_0000_0000_0000;
array[14317] <= 16'b0000_0000_0000_0000;
array[14318] <= 16'b0000_0000_0000_0000;
array[14319] <= 16'b0000_0000_0000_0000;
array[14320] <= 16'b0000_0000_0000_0000;
array[14321] <= 16'b0000_0000_0000_0000;
array[14322] <= 16'b0000_0000_0000_0000;
array[14323] <= 16'b0000_0000_0000_0000;
array[14324] <= 16'b0000_0000_0000_0000;
array[14325] <= 16'b0000_0000_0000_0000;
array[14326] <= 16'b0000_0000_0000_0000;
array[14327] <= 16'b0000_0000_0000_0000;
array[14328] <= 16'b0000_0000_0000_0000;
array[14329] <= 16'b0000_0000_0000_0000;
array[14330] <= 16'b0000_0000_0000_0000;
array[14331] <= 16'b0000_0000_0000_0000;
array[14332] <= 16'b0000_0000_0000_0000;
array[14333] <= 16'b0000_0000_0000_0000;
array[14334] <= 16'b0000_0000_0000_0000;
array[14335] <= 16'b0000_0000_0000_0000;
array[14336] <= 16'b0000_0000_0000_0000;
array[14337] <= 16'b0000_0000_0000_0000;
array[14338] <= 16'b0000_0000_0000_0000;
array[14339] <= 16'b0000_0000_0000_0000;
array[14340] <= 16'b0000_0000_0000_0000;
array[14341] <= 16'b0000_0000_0000_0000;
array[14342] <= 16'b0000_0000_0000_0000;
array[14343] <= 16'b0000_0000_0000_0000;
array[14344] <= 16'b0000_0000_0000_0000;
array[14345] <= 16'b0000_0000_0000_0000;
array[14346] <= 16'b0000_0000_0000_0000;
array[14347] <= 16'b0000_0000_0000_0000;
array[14348] <= 16'b0000_0000_0000_0000;
array[14349] <= 16'b0000_0000_0000_0000;
array[14350] <= 16'b0000_0000_0000_0000;
array[14351] <= 16'b0000_0000_0000_0000;
array[14352] <= 16'b0000_0000_0000_0000;
array[14353] <= 16'b0000_0000_0000_0000;
array[14354] <= 16'b0000_0000_0000_0000;
array[14355] <= 16'b0000_0000_0000_0000;
array[14356] <= 16'b0000_0000_0000_0000;
array[14357] <= 16'b0000_0000_0000_0000;
array[14358] <= 16'b0000_0000_0000_0000;
array[14359] <= 16'b0000_0000_0000_0000;
array[14360] <= 16'b0000_0000_0000_0000;
array[14361] <= 16'b0000_0000_0000_0000;
array[14362] <= 16'b0000_0000_0000_0000;
array[14363] <= 16'b0000_0000_0000_0000;
array[14364] <= 16'b0000_0000_0000_0000;
array[14365] <= 16'b0000_0000_0000_0000;
array[14366] <= 16'b0000_0000_0000_0000;
array[14367] <= 16'b0000_0000_0000_0000;
array[14368] <= 16'b0000_0000_0000_0000;
array[14369] <= 16'b0000_0000_0000_0000;
array[14370] <= 16'b0000_0000_0000_0000;
array[14371] <= 16'b0000_0000_0000_0000;
array[14372] <= 16'b0000_0000_0000_0000;
array[14373] <= 16'b0000_0000_0000_0000;
array[14374] <= 16'b0000_0000_0000_0000;
array[14375] <= 16'b0000_0000_0000_0000;
array[14376] <= 16'b0000_0000_0000_0000;
array[14377] <= 16'b0000_0000_0000_0000;
array[14378] <= 16'b0000_0000_0000_0000;
array[14379] <= 16'b0000_0000_0000_0000;
array[14380] <= 16'b0000_0000_0000_0000;
array[14381] <= 16'b0000_0000_0000_0000;
array[14382] <= 16'b0000_0000_0000_0000;
array[14383] <= 16'b0000_0000_0000_0000;
array[14384] <= 16'b0000_0000_0000_0000;
array[14385] <= 16'b0000_0000_0000_0000;
array[14386] <= 16'b0000_0000_0000_0000;
array[14387] <= 16'b0000_0000_0000_0000;
array[14388] <= 16'b0000_0000_0000_0000;
array[14389] <= 16'b0000_0000_0000_0000;
array[14390] <= 16'b0000_0000_0000_0000;
array[14391] <= 16'b0000_0000_0000_0000;
array[14392] <= 16'b0000_0000_0000_0000;
array[14393] <= 16'b0000_0000_0000_0000;
array[14394] <= 16'b0000_0000_0000_0000;
array[14395] <= 16'b0000_0000_0000_0000;
array[14396] <= 16'b0000_0000_0000_0000;
array[14397] <= 16'b0000_0000_0000_0000;
array[14398] <= 16'b0000_0000_0000_0000;
array[14399] <= 16'b0000_0000_0000_0000;
array[14400] <= 16'b0000_0000_0000_0000;
array[14401] <= 16'b0000_0000_0000_0000;
array[14402] <= 16'b0000_0000_0000_0000;
array[14403] <= 16'b0000_0000_0000_0000;
array[14404] <= 16'b0000_0000_0000_0000;
array[14405] <= 16'b0000_0000_0000_0000;
array[14406] <= 16'b0000_0000_0000_0000;
array[14407] <= 16'b0000_0000_0000_0000;
array[14408] <= 16'b0000_0000_0000_0000;
array[14409] <= 16'b0000_0000_0000_0000;
array[14410] <= 16'b0000_0000_0000_0000;
array[14411] <= 16'b0000_0000_0000_0000;
array[14412] <= 16'b0000_0000_0000_0000;
array[14413] <= 16'b0000_0000_0000_0000;
array[14414] <= 16'b0000_0000_0000_0000;
array[14415] <= 16'b0000_0000_0000_0000;
array[14416] <= 16'b0000_0000_0000_0000;
array[14417] <= 16'b0000_0000_0000_0000;
array[14418] <= 16'b0000_0000_0000_0000;
array[14419] <= 16'b0000_0000_0000_0000;
array[14420] <= 16'b0000_0000_0000_0000;
array[14421] <= 16'b0000_0000_0000_0000;
array[14422] <= 16'b0000_0000_0000_0000;
array[14423] <= 16'b0000_0000_0000_0000;
array[14424] <= 16'b0000_0000_0000_0000;
array[14425] <= 16'b0000_0000_0000_0000;
array[14426] <= 16'b0000_0000_0000_0000;
array[14427] <= 16'b0000_0000_0000_0000;
array[14428] <= 16'b0000_0000_0000_0000;
array[14429] <= 16'b0000_0000_0000_0000;
array[14430] <= 16'b0000_0000_0000_0000;
array[14431] <= 16'b0000_0000_0000_0000;
array[14432] <= 16'b0000_0000_0000_0000;
array[14433] <= 16'b0000_0000_0000_0000;
array[14434] <= 16'b0000_0000_0000_0000;
array[14435] <= 16'b0000_0000_0000_0000;
array[14436] <= 16'b0000_0000_0000_0000;
array[14437] <= 16'b0000_0000_0000_0000;
array[14438] <= 16'b0000_0000_0000_0000;
array[14439] <= 16'b0000_0000_0000_0000;
array[14440] <= 16'b0000_0000_0000_0000;
array[14441] <= 16'b0000_0000_0000_0000;
array[14442] <= 16'b0000_0000_0000_0000;
array[14443] <= 16'b0000_0000_0000_0000;
array[14444] <= 16'b0000_0000_0000_0000;
array[14445] <= 16'b0000_0000_0000_0000;
array[14446] <= 16'b0000_0000_0000_0000;
array[14447] <= 16'b0000_0000_0000_0000;
array[14448] <= 16'b0000_0000_0000_0000;
array[14449] <= 16'b0000_0000_0000_0000;
array[14450] <= 16'b0000_0000_0000_0000;
array[14451] <= 16'b0000_0000_0000_0000;
array[14452] <= 16'b0000_0000_0000_0000;
array[14453] <= 16'b0000_0000_0000_0000;
array[14454] <= 16'b0000_0000_0000_0000;
array[14455] <= 16'b0000_0000_0000_0000;
array[14456] <= 16'b0000_0000_0000_0000;
array[14457] <= 16'b0000_0000_0000_0000;
array[14458] <= 16'b0000_0000_0000_0000;
array[14459] <= 16'b0000_0000_0000_0000;
array[14460] <= 16'b0000_0000_0000_0000;
array[14461] <= 16'b0000_0000_0000_0000;
array[14462] <= 16'b0000_0000_0000_0000;
array[14463] <= 16'b0000_0000_0000_0000;
array[14464] <= 16'b0000_0000_0000_0000;
array[14465] <= 16'b0000_0000_0000_0000;
array[14466] <= 16'b0000_0000_0000_0000;
array[14467] <= 16'b0000_0000_0000_0000;
array[14468] <= 16'b0000_0000_0000_0000;
array[14469] <= 16'b0000_0000_0000_0000;
array[14470] <= 16'b0000_0000_0000_0000;
array[14471] <= 16'b0000_0000_0000_0000;
array[14472] <= 16'b0000_0000_0000_0000;
array[14473] <= 16'b0000_0000_0000_0000;
array[14474] <= 16'b0000_0000_0000_0000;
array[14475] <= 16'b0000_0000_0000_0000;
array[14476] <= 16'b0000_0000_0000_0000;
array[14477] <= 16'b0000_0000_0000_0000;
array[14478] <= 16'b0000_0000_0000_0000;
array[14479] <= 16'b0000_0000_0000_0000;
array[14480] <= 16'b0000_0000_0000_0000;
array[14481] <= 16'b0000_0000_0000_0000;
array[14482] <= 16'b0000_0000_0000_0000;
array[14483] <= 16'b0000_0000_0000_0000;
array[14484] <= 16'b0000_0000_0000_0000;
array[14485] <= 16'b0000_0000_0000_0000;
array[14486] <= 16'b0000_0000_0000_0000;
array[14487] <= 16'b0000_0000_0000_0000;
array[14488] <= 16'b0000_0000_0000_0000;
array[14489] <= 16'b0000_0000_0000_0000;
array[14490] <= 16'b0000_0000_0000_0000;
array[14491] <= 16'b0000_0000_0000_0000;
array[14492] <= 16'b0000_0000_0000_0000;
array[14493] <= 16'b0000_0000_0000_0000;
array[14494] <= 16'b0000_0000_0000_0000;
array[14495] <= 16'b0000_0000_0000_0000;
array[14496] <= 16'b0000_0000_0000_0000;
array[14497] <= 16'b0000_0000_0000_0000;
array[14498] <= 16'b0000_0000_0000_0000;
array[14499] <= 16'b0000_0000_0000_0000;
array[14500] <= 16'b0000_0000_0000_0000;
array[14501] <= 16'b0000_0000_0000_0000;
array[14502] <= 16'b0000_0000_0000_0000;
array[14503] <= 16'b0000_0000_0000_0000;
array[14504] <= 16'b0000_0000_0000_0000;
array[14505] <= 16'b0000_0000_0000_0000;
array[14506] <= 16'b0000_0000_0000_0000;
array[14507] <= 16'b0000_0000_0000_0000;
array[14508] <= 16'b0000_0000_0000_0000;
array[14509] <= 16'b0000_0000_0000_0000;
array[14510] <= 16'b0000_0000_0000_0000;
array[14511] <= 16'b0000_0000_0000_0000;
array[14512] <= 16'b0000_0000_0000_0000;
array[14513] <= 16'b0000_0000_0000_0000;
array[14514] <= 16'b0000_0000_0000_0000;
array[14515] <= 16'b0000_0000_0000_0000;
array[14516] <= 16'b0000_0000_0000_0000;
array[14517] <= 16'b0000_0000_0000_0000;
array[14518] <= 16'b0000_0000_0000_0000;
array[14519] <= 16'b0000_0000_0000_0000;
array[14520] <= 16'b0000_0000_0000_0000;
array[14521] <= 16'b0000_0000_0000_0000;
array[14522] <= 16'b0000_0000_0000_0000;
array[14523] <= 16'b0000_0000_0000_0000;
array[14524] <= 16'b0000_0000_0000_0000;
array[14525] <= 16'b0000_0000_0000_0000;
array[14526] <= 16'b0000_0000_0000_0000;
array[14527] <= 16'b0000_0000_0000_0000;
array[14528] <= 16'b0000_0000_0000_0000;
array[14529] <= 16'b0000_0000_0000_0000;
array[14530] <= 16'b0000_0000_0000_0000;
array[14531] <= 16'b0000_0000_0000_0000;
array[14532] <= 16'b0000_0000_0000_0000;
array[14533] <= 16'b0000_0000_0000_0000;
array[14534] <= 16'b0000_0000_0000_0000;
array[14535] <= 16'b0000_0000_0000_0000;
array[14536] <= 16'b0000_0000_0000_0000;
array[14537] <= 16'b0000_0000_0000_0000;
array[14538] <= 16'b0000_0000_0000_0000;
array[14539] <= 16'b0000_0000_0000_0000;
array[14540] <= 16'b0000_0000_0000_0000;
array[14541] <= 16'b0000_0000_0000_0000;
array[14542] <= 16'b0000_0000_0000_0000;
array[14543] <= 16'b0000_0000_0000_0000;
array[14544] <= 16'b0000_0000_0000_0000;
array[14545] <= 16'b0000_0000_0000_0000;
array[14546] <= 16'b0000_0000_0000_0000;
array[14547] <= 16'b0000_0000_0000_0000;
array[14548] <= 16'b0000_0000_0000_0000;
array[14549] <= 16'b0000_0000_0000_0000;
array[14550] <= 16'b0000_0000_0000_0000;
array[14551] <= 16'b0000_0000_0000_0000;
array[14552] <= 16'b0000_0000_0000_0000;
array[14553] <= 16'b0000_0000_0000_0000;
array[14554] <= 16'b0000_0000_0000_0000;
array[14555] <= 16'b0000_0000_0000_0000;
array[14556] <= 16'b0000_0000_0000_0000;
array[14557] <= 16'b0000_0000_0000_0000;
array[14558] <= 16'b0000_0000_0000_0000;
array[14559] <= 16'b0000_0000_0000_0000;
array[14560] <= 16'b0000_0000_0000_0000;
array[14561] <= 16'b0000_0000_0000_0000;
array[14562] <= 16'b0000_0000_0000_0000;
array[14563] <= 16'b0000_0000_0000_0000;
array[14564] <= 16'b0000_0000_0000_0000;
array[14565] <= 16'b0000_0000_0000_0000;
array[14566] <= 16'b0000_0000_0000_0000;
array[14567] <= 16'b0000_0000_0000_0000;
array[14568] <= 16'b0000_0000_0000_0000;
array[14569] <= 16'b0000_0000_0000_0000;
array[14570] <= 16'b0000_0000_0000_0000;
array[14571] <= 16'b0000_0000_0000_0000;
array[14572] <= 16'b0000_0000_0000_0000;
array[14573] <= 16'b0000_0000_0000_0000;
array[14574] <= 16'b0000_0000_0000_0000;
array[14575] <= 16'b0000_0000_0000_0000;
array[14576] <= 16'b0000_0000_0000_0000;
array[14577] <= 16'b0000_0000_0000_0000;
array[14578] <= 16'b0000_0000_0000_0000;
array[14579] <= 16'b0000_0000_0000_0000;
array[14580] <= 16'b0000_0000_0000_0000;
array[14581] <= 16'b0000_0000_0000_0000;
array[14582] <= 16'b0000_0000_0000_0000;
array[14583] <= 16'b0000_0000_0000_0000;
array[14584] <= 16'b0000_0000_0000_0000;
array[14585] <= 16'b0000_0000_0000_0000;
array[14586] <= 16'b0000_0000_0000_0000;
array[14587] <= 16'b0000_0000_0000_0000;
array[14588] <= 16'b0000_0000_0000_0000;
array[14589] <= 16'b0000_0000_0000_0000;
array[14590] <= 16'b0000_0000_0000_0000;
array[14591] <= 16'b0000_0000_0000_0000;
array[14592] <= 16'b0000_0000_0000_0000;
array[14593] <= 16'b0000_0000_0000_0000;
array[14594] <= 16'b0000_0000_0000_0000;
array[14595] <= 16'b0000_0000_0000_0000;
array[14596] <= 16'b0000_0000_0000_0000;
array[14597] <= 16'b0000_0000_0000_0000;
array[14598] <= 16'b0000_0000_0000_0000;
array[14599] <= 16'b0000_0000_0000_0000;
array[14600] <= 16'b0000_0000_0000_0000;
array[14601] <= 16'b0000_0000_0000_0000;
array[14602] <= 16'b0000_0000_0000_0000;
array[14603] <= 16'b0000_0000_0000_0000;
array[14604] <= 16'b0000_0000_0000_0000;
array[14605] <= 16'b0000_0000_0000_0000;
array[14606] <= 16'b0000_0000_0000_0000;
array[14607] <= 16'b0000_0000_0000_0000;
array[14608] <= 16'b0000_0000_0000_0000;
array[14609] <= 16'b0000_0000_0000_0000;
array[14610] <= 16'b0000_0000_0000_0000;
array[14611] <= 16'b0000_0000_0000_0000;
array[14612] <= 16'b0000_0000_0000_0000;
array[14613] <= 16'b0000_0000_0000_0000;
array[14614] <= 16'b0000_0000_0000_0000;
array[14615] <= 16'b0000_0000_0000_0000;
array[14616] <= 16'b0000_0000_0000_0000;
array[14617] <= 16'b0000_0000_0000_0000;
array[14618] <= 16'b0000_0000_0000_0000;
array[14619] <= 16'b0000_0000_0000_0000;
array[14620] <= 16'b0000_0000_0000_0000;
array[14621] <= 16'b0000_0000_0000_0000;
array[14622] <= 16'b0000_0000_0000_0000;
array[14623] <= 16'b0000_0000_0000_0000;
array[14624] <= 16'b0000_0000_0000_0000;
array[14625] <= 16'b0000_0000_0000_0000;
array[14626] <= 16'b0000_0000_0000_0000;
array[14627] <= 16'b0000_0000_0000_0000;
array[14628] <= 16'b0000_0000_0000_0000;
array[14629] <= 16'b0000_0000_0000_0000;
array[14630] <= 16'b0000_0000_0000_0000;
array[14631] <= 16'b0000_0000_0000_0000;
array[14632] <= 16'b0000_0000_0000_0000;
array[14633] <= 16'b0000_0000_0000_0000;
array[14634] <= 16'b0000_0000_0000_0000;
array[14635] <= 16'b0000_0000_0000_0000;
array[14636] <= 16'b0000_0000_0000_0000;
array[14637] <= 16'b0000_0000_0000_0000;
array[14638] <= 16'b0000_0000_0000_0000;
array[14639] <= 16'b0000_0000_0000_0000;
array[14640] <= 16'b0000_0000_0000_0000;
array[14641] <= 16'b0000_0000_0000_0000;
array[14642] <= 16'b0000_0000_0000_0000;
array[14643] <= 16'b0000_0000_0000_0000;
array[14644] <= 16'b0000_0000_0000_0000;
array[14645] <= 16'b0000_0000_0000_0000;
array[14646] <= 16'b0000_0000_0000_0000;
array[14647] <= 16'b0000_0000_0000_0000;
array[14648] <= 16'b0000_0000_0000_0000;
array[14649] <= 16'b0000_0000_0000_0000;
array[14650] <= 16'b0000_0000_0000_0000;
array[14651] <= 16'b0000_0000_0000_0000;
array[14652] <= 16'b0000_0000_0000_0000;
array[14653] <= 16'b0000_0000_0000_0000;
array[14654] <= 16'b0000_0000_0000_0000;
array[14655] <= 16'b0000_0000_0000_0000;
array[14656] <= 16'b0000_0000_0000_0000;
array[14657] <= 16'b0000_0000_0000_0000;
array[14658] <= 16'b0000_0000_0000_0000;
array[14659] <= 16'b0000_0000_0000_0000;
array[14660] <= 16'b0000_0000_0000_0000;
array[14661] <= 16'b0000_0000_0000_0000;
array[14662] <= 16'b0000_0000_0000_0000;
array[14663] <= 16'b0000_0000_0000_0000;
array[14664] <= 16'b0000_0000_0000_0000;
array[14665] <= 16'b0000_0000_0000_0000;
array[14666] <= 16'b0000_0000_0000_0000;
array[14667] <= 16'b0000_0000_0000_0000;
array[14668] <= 16'b0000_0000_0000_0000;
array[14669] <= 16'b0000_0000_0000_0000;
array[14670] <= 16'b0000_0000_0000_0000;
array[14671] <= 16'b0000_0000_0000_0000;
array[14672] <= 16'b0000_0000_0000_0000;
array[14673] <= 16'b0000_0000_0000_0000;
array[14674] <= 16'b0000_0000_0000_0000;
array[14675] <= 16'b0000_0000_0000_0000;
array[14676] <= 16'b0000_0000_0000_0000;
array[14677] <= 16'b0000_0000_0000_0000;
array[14678] <= 16'b0000_0000_0000_0000;
array[14679] <= 16'b0000_0000_0000_0000;
array[14680] <= 16'b0000_0000_0000_0000;
array[14681] <= 16'b0000_0000_0000_0000;
array[14682] <= 16'b0000_0000_0000_0000;
array[14683] <= 16'b0000_0000_0000_0000;
array[14684] <= 16'b0000_0000_0000_0000;
array[14685] <= 16'b0000_0000_0000_0000;
array[14686] <= 16'b0000_0000_0000_0000;
array[14687] <= 16'b0000_0000_0000_0000;
array[14688] <= 16'b0000_0000_0000_0000;
array[14689] <= 16'b0000_0000_0000_0000;
array[14690] <= 16'b0000_0000_0000_0000;
array[14691] <= 16'b0000_0000_0000_0000;
array[14692] <= 16'b0000_0000_0000_0000;
array[14693] <= 16'b0000_0000_0000_0000;
array[14694] <= 16'b0000_0000_0000_0000;
array[14695] <= 16'b0000_0000_0000_0000;
array[14696] <= 16'b0000_0000_0000_0000;
array[14697] <= 16'b0000_0000_0000_0000;
array[14698] <= 16'b0000_0000_0000_0000;
array[14699] <= 16'b0000_0000_0000_0000;
array[14700] <= 16'b0000_0000_0000_0000;
array[14701] <= 16'b0000_0000_0000_0000;
array[14702] <= 16'b0000_0000_0000_0000;
array[14703] <= 16'b0000_0000_0000_0000;
array[14704] <= 16'b0000_0000_0000_0000;
array[14705] <= 16'b0000_0000_0000_0000;
array[14706] <= 16'b0000_0000_0000_0000;
array[14707] <= 16'b0000_0000_0000_0000;
array[14708] <= 16'b0000_0000_0000_0000;
array[14709] <= 16'b0000_0000_0000_0000;
array[14710] <= 16'b0000_0000_0000_0000;
array[14711] <= 16'b0000_0000_0000_0000;
array[14712] <= 16'b0000_0000_0000_0000;
array[14713] <= 16'b0000_0000_0000_0000;
array[14714] <= 16'b0000_0000_0000_0000;
array[14715] <= 16'b0000_0000_0000_0000;
array[14716] <= 16'b0000_0000_0000_0000;
array[14717] <= 16'b0000_0000_0000_0000;
array[14718] <= 16'b0000_0000_0000_0000;
array[14719] <= 16'b0000_0000_0000_0000;
array[14720] <= 16'b0000_0000_0000_0000;
array[14721] <= 16'b0000_0000_0000_0000;
array[14722] <= 16'b0000_0000_0000_0000;
array[14723] <= 16'b0000_0000_0000_0000;
array[14724] <= 16'b0000_0000_0000_0000;
array[14725] <= 16'b0000_0000_0000_0000;
array[14726] <= 16'b0000_0000_0000_0000;
array[14727] <= 16'b0000_0000_0000_0000;
array[14728] <= 16'b0000_0000_0000_0000;
array[14729] <= 16'b0000_0000_0000_0000;
array[14730] <= 16'b0000_0000_0000_0000;
array[14731] <= 16'b0000_0000_0000_0000;
array[14732] <= 16'b0000_0000_0000_0000;
array[14733] <= 16'b0000_0000_0000_0000;
array[14734] <= 16'b0000_0000_0000_0000;
array[14735] <= 16'b0000_0000_0000_0000;
array[14736] <= 16'b0000_0000_0000_0000;
array[14737] <= 16'b0000_0000_0000_0000;
array[14738] <= 16'b0000_0000_0000_0000;
array[14739] <= 16'b0000_0000_0000_0000;
array[14740] <= 16'b0000_0000_0000_0000;
array[14741] <= 16'b0000_0000_0000_0000;
array[14742] <= 16'b0000_0000_0000_0000;
array[14743] <= 16'b0000_0000_0000_0000;
array[14744] <= 16'b0000_0000_0000_0000;
array[14745] <= 16'b0000_0000_0000_0000;
array[14746] <= 16'b0000_0000_0000_0000;
array[14747] <= 16'b0000_0000_0000_0000;
array[14748] <= 16'b0000_0000_0000_0000;
array[14749] <= 16'b0000_0000_0000_0000;
array[14750] <= 16'b0000_0000_0000_0000;
array[14751] <= 16'b0000_0000_0000_0000;
array[14752] <= 16'b0000_0000_0000_0000;
array[14753] <= 16'b0000_0000_0000_0000;
array[14754] <= 16'b0000_0000_0000_0000;
array[14755] <= 16'b0000_0000_0000_0000;
array[14756] <= 16'b0000_0000_0000_0000;
array[14757] <= 16'b0000_0000_0000_0000;
array[14758] <= 16'b0000_0000_0000_0000;
array[14759] <= 16'b0000_0000_0000_0000;
array[14760] <= 16'b0000_0000_0000_0000;
array[14761] <= 16'b0000_0000_0000_0000;
array[14762] <= 16'b0000_0000_0000_0000;
array[14763] <= 16'b0000_0000_0000_0000;
array[14764] <= 16'b0000_0000_0000_0000;
array[14765] <= 16'b0000_0000_0000_0000;
array[14766] <= 16'b0000_0000_0000_0000;
array[14767] <= 16'b0000_0000_0000_0000;
array[14768] <= 16'b0000_0000_0000_0000;
array[14769] <= 16'b0000_0000_0000_0000;
array[14770] <= 16'b0000_0000_0000_0000;
array[14771] <= 16'b0000_0000_0000_0000;
array[14772] <= 16'b0000_0000_0000_0000;
array[14773] <= 16'b0000_0000_0000_0000;
array[14774] <= 16'b0000_0000_0000_0000;
array[14775] <= 16'b0000_0000_0000_0000;
array[14776] <= 16'b0000_0000_0000_0000;
array[14777] <= 16'b0000_0000_0000_0000;
array[14778] <= 16'b0000_0000_0000_0000;
array[14779] <= 16'b0000_0000_0000_0000;
array[14780] <= 16'b0000_0000_0000_0000;
array[14781] <= 16'b0000_0000_0000_0000;
array[14782] <= 16'b0000_0000_0000_0000;
array[14783] <= 16'b0000_0000_0000_0000;
array[14784] <= 16'b0000_0000_0000_0000;
array[14785] <= 16'b0000_0000_0000_0000;
array[14786] <= 16'b0000_0000_0000_0000;
array[14787] <= 16'b0000_0000_0000_0000;
array[14788] <= 16'b0000_0000_0000_0000;
array[14789] <= 16'b0000_0000_0000_0000;
array[14790] <= 16'b0000_0000_0000_0000;
array[14791] <= 16'b0000_0000_0000_0000;
array[14792] <= 16'b0000_0000_0000_0000;
array[14793] <= 16'b0000_0000_0000_0000;
array[14794] <= 16'b0000_0000_0000_0000;
array[14795] <= 16'b0000_0000_0000_0000;
array[14796] <= 16'b0000_0000_0000_0000;
array[14797] <= 16'b0000_0000_0000_0000;
array[14798] <= 16'b0000_0000_0000_0000;
array[14799] <= 16'b0000_0000_0000_0000;
array[14800] <= 16'b0000_0000_0000_0000;
array[14801] <= 16'b0000_0000_0000_0000;
array[14802] <= 16'b0000_0000_0000_0000;
array[14803] <= 16'b0000_0000_0000_0000;
array[14804] <= 16'b0000_0000_0000_0000;
array[14805] <= 16'b0000_0000_0000_0000;
array[14806] <= 16'b0000_0000_0000_0000;
array[14807] <= 16'b0000_0000_0000_0000;
array[14808] <= 16'b0000_0000_0000_0000;
array[14809] <= 16'b0000_0000_0000_0000;
array[14810] <= 16'b0000_0000_0000_0000;
array[14811] <= 16'b0000_0000_0000_0000;
array[14812] <= 16'b0000_0000_0000_0000;
array[14813] <= 16'b0000_0000_0000_0000;
array[14814] <= 16'b0000_0000_0000_0000;
array[14815] <= 16'b0000_0000_0000_0000;
array[14816] <= 16'b0000_0000_0000_0000;
array[14817] <= 16'b0000_0000_0000_0000;
array[14818] <= 16'b0000_0000_0000_0000;
array[14819] <= 16'b0000_0000_0000_0000;
array[14820] <= 16'b0000_0000_0000_0000;
array[14821] <= 16'b0000_0000_0000_0000;
array[14822] <= 16'b0000_0000_0000_0000;
array[14823] <= 16'b0000_0000_0000_0000;
array[14824] <= 16'b0000_0000_0000_0000;
array[14825] <= 16'b0000_0000_0000_0000;
array[14826] <= 16'b0000_0000_0000_0000;
array[14827] <= 16'b0000_0000_0000_0000;
array[14828] <= 16'b0000_0000_0000_0000;
array[14829] <= 16'b0000_0000_0000_0000;
array[14830] <= 16'b0000_0000_0000_0000;
array[14831] <= 16'b0000_0000_0000_0000;
array[14832] <= 16'b0000_0000_0000_0000;
array[14833] <= 16'b0000_0000_0000_0000;
array[14834] <= 16'b0000_0000_0000_0000;
array[14835] <= 16'b0000_0000_0000_0000;
array[14836] <= 16'b0000_0000_0000_0000;
array[14837] <= 16'b0000_0000_0000_0000;
array[14838] <= 16'b0000_0000_0000_0000;
array[14839] <= 16'b0000_0000_0000_0000;
array[14840] <= 16'b0000_0000_0000_0000;
array[14841] <= 16'b0000_0000_0000_0000;
array[14842] <= 16'b0000_0000_0000_0000;
array[14843] <= 16'b0000_0000_0000_0000;
array[14844] <= 16'b0000_0000_0000_0000;
array[14845] <= 16'b0000_0000_0000_0000;
array[14846] <= 16'b0000_0000_0000_0000;
array[14847] <= 16'b0000_0000_0000_0000;
array[14848] <= 16'b0000_0000_0000_0000;
array[14849] <= 16'b0000_0000_0000_0000;
array[14850] <= 16'b0000_0000_0000_0000;
array[14851] <= 16'b0000_0000_0000_0000;
array[14852] <= 16'b0000_0000_0000_0000;
array[14853] <= 16'b0000_0000_0000_0000;
array[14854] <= 16'b0000_0000_0000_0000;
array[14855] <= 16'b0000_0000_0000_0000;
array[14856] <= 16'b0000_0000_0000_0000;
array[14857] <= 16'b0000_0000_0000_0000;
array[14858] <= 16'b0000_0000_0000_0000;
array[14859] <= 16'b0000_0000_0000_0000;
array[14860] <= 16'b0000_0000_0000_0000;
array[14861] <= 16'b0000_0000_0000_0000;
array[14862] <= 16'b0000_0000_0000_0000;
array[14863] <= 16'b0000_0000_0000_0000;
array[14864] <= 16'b0000_0000_0000_0000;
array[14865] <= 16'b0000_0000_0000_0000;
array[14866] <= 16'b0000_0000_0000_0000;
array[14867] <= 16'b0000_0000_0000_0000;
array[14868] <= 16'b0000_0000_0000_0000;
array[14869] <= 16'b0000_0000_0000_0000;
array[14870] <= 16'b0000_0000_0000_0000;
array[14871] <= 16'b0000_0000_0000_0000;
array[14872] <= 16'b0000_0000_0000_0000;
array[14873] <= 16'b0000_0000_0000_0000;
array[14874] <= 16'b0000_0000_0000_0000;
array[14875] <= 16'b0000_0000_0000_0000;
array[14876] <= 16'b0000_0000_0000_0000;
array[14877] <= 16'b0000_0000_0000_0000;
array[14878] <= 16'b0000_0000_0000_0000;
array[14879] <= 16'b0000_0000_0000_0000;
array[14880] <= 16'b0000_0000_0000_0000;
array[14881] <= 16'b0000_0000_0000_0000;
array[14882] <= 16'b0000_0000_0000_0000;
array[14883] <= 16'b0000_0000_0000_0000;
array[14884] <= 16'b0000_0000_0000_0000;
array[14885] <= 16'b0000_0000_0000_0000;
array[14886] <= 16'b0000_0000_0000_0000;
array[14887] <= 16'b0000_0000_0000_0000;
array[14888] <= 16'b0000_0000_0000_0000;
array[14889] <= 16'b0000_0000_0000_0000;
array[14890] <= 16'b0000_0000_0000_0000;
array[14891] <= 16'b0000_0000_0000_0000;
array[14892] <= 16'b0000_0000_0000_0000;
array[14893] <= 16'b0000_0000_0000_0000;
array[14894] <= 16'b0000_0000_0000_0000;
array[14895] <= 16'b0000_0000_0000_0000;
array[14896] <= 16'b0000_0000_0000_0000;
array[14897] <= 16'b0000_0000_0000_0000;
array[14898] <= 16'b0000_0000_0000_0000;
array[14899] <= 16'b0000_0000_0000_0000;
array[14900] <= 16'b0000_0000_0000_0000;
array[14901] <= 16'b0000_0000_0000_0000;
array[14902] <= 16'b0000_0000_0000_0000;
array[14903] <= 16'b0000_0000_0000_0000;
array[14904] <= 16'b0000_0000_0000_0000;
array[14905] <= 16'b0000_0000_0000_0000;
array[14906] <= 16'b0000_0000_0000_0000;
array[14907] <= 16'b0000_0000_0000_0000;
array[14908] <= 16'b0000_0000_0000_0000;
array[14909] <= 16'b0000_0000_0000_0000;
array[14910] <= 16'b0000_0000_0000_0000;
array[14911] <= 16'b0000_0000_0000_0000;
array[14912] <= 16'b0000_0000_0000_0000;
array[14913] <= 16'b0000_0000_0000_0000;
array[14914] <= 16'b0000_0000_0000_0000;
array[14915] <= 16'b0000_0000_0000_0000;
array[14916] <= 16'b0000_0000_0000_0000;
array[14917] <= 16'b0000_0000_0000_0000;
array[14918] <= 16'b0000_0000_0000_0000;
array[14919] <= 16'b0000_0000_0000_0000;
array[14920] <= 16'b0000_0000_0000_0000;
array[14921] <= 16'b0000_0000_0000_0000;
array[14922] <= 16'b0000_0000_0000_0000;
array[14923] <= 16'b0000_0000_0000_0000;
array[14924] <= 16'b0000_0000_0000_0000;
array[14925] <= 16'b0000_0000_0000_0000;
array[14926] <= 16'b0000_0000_0000_0000;
array[14927] <= 16'b0000_0000_0000_0000;
array[14928] <= 16'b0000_0000_0000_0000;
array[14929] <= 16'b0000_0000_0000_0000;
array[14930] <= 16'b0000_0000_0000_0000;
array[14931] <= 16'b0000_0000_0000_0000;
array[14932] <= 16'b0000_0000_0000_0000;
array[14933] <= 16'b0000_0000_0000_0000;
array[14934] <= 16'b0000_0000_0000_0000;
array[14935] <= 16'b0000_0000_0000_0000;
array[14936] <= 16'b0000_0000_0000_0000;
array[14937] <= 16'b0000_0000_0000_0000;
array[14938] <= 16'b0000_0000_0000_0000;
array[14939] <= 16'b0000_0000_0000_0000;
array[14940] <= 16'b0000_0000_0000_0000;
array[14941] <= 16'b0000_0000_0000_0000;
array[14942] <= 16'b0000_0000_0000_0000;
array[14943] <= 16'b0000_0000_0000_0000;
array[14944] <= 16'b0000_0000_0000_0000;
array[14945] <= 16'b0000_0000_0000_0000;
array[14946] <= 16'b0000_0000_0000_0000;
array[14947] <= 16'b0000_0000_0000_0000;
array[14948] <= 16'b0000_0000_0000_0000;
array[14949] <= 16'b0000_0000_0000_0000;
array[14950] <= 16'b0000_0000_0000_0000;
array[14951] <= 16'b0000_0000_0000_0000;
array[14952] <= 16'b0000_0000_0000_0000;
array[14953] <= 16'b0000_0000_0000_0000;
array[14954] <= 16'b0000_0000_0000_0000;
array[14955] <= 16'b0000_0000_0000_0000;
array[14956] <= 16'b0000_0000_0000_0000;
array[14957] <= 16'b0000_0000_0000_0000;
array[14958] <= 16'b0000_0000_0000_0000;
array[14959] <= 16'b0000_0000_0000_0000;
array[14960] <= 16'b0000_0000_0000_0000;
array[14961] <= 16'b0000_0000_0000_0000;
array[14962] <= 16'b0000_0000_0000_0000;
array[14963] <= 16'b0000_0000_0000_0000;
array[14964] <= 16'b0000_0000_0000_0000;
array[14965] <= 16'b0000_0000_0000_0000;
array[14966] <= 16'b0000_0000_0000_0000;
array[14967] <= 16'b0000_0000_0000_0000;
array[14968] <= 16'b0000_0000_0000_0000;
array[14969] <= 16'b0000_0000_0000_0000;
array[14970] <= 16'b0000_0000_0000_0000;
array[14971] <= 16'b0000_0000_0000_0000;
array[14972] <= 16'b0000_0000_0000_0000;
array[14973] <= 16'b0000_0000_0000_0000;
array[14974] <= 16'b0000_0000_0000_0000;
array[14975] <= 16'b0000_0000_0000_0000;
array[14976] <= 16'b0000_0000_0000_0000;
array[14977] <= 16'b0000_0000_0000_0000;
array[14978] <= 16'b0000_0000_0000_0000;
array[14979] <= 16'b0000_0000_0000_0000;
array[14980] <= 16'b0000_0000_0000_0000;
array[14981] <= 16'b0000_0000_0000_0000;
array[14982] <= 16'b0000_0000_0000_0000;
array[14983] <= 16'b0000_0000_0000_0000;
array[14984] <= 16'b0000_0000_0000_0000;
array[14985] <= 16'b0000_0000_0000_0000;
array[14986] <= 16'b0000_0000_0000_0000;
array[14987] <= 16'b0000_0000_0000_0000;
array[14988] <= 16'b0000_0000_0000_0000;
array[14989] <= 16'b0000_0000_0000_0000;
array[14990] <= 16'b0000_0000_0000_0000;
array[14991] <= 16'b0000_0000_0000_0000;
array[14992] <= 16'b0000_0000_0000_0000;
array[14993] <= 16'b0000_0000_0000_0000;
array[14994] <= 16'b0000_0000_0000_0000;
array[14995] <= 16'b0000_0000_0000_0000;
array[14996] <= 16'b0000_0000_0000_0000;
array[14997] <= 16'b0000_0000_0000_0000;
array[14998] <= 16'b0000_0000_0000_0000;
array[14999] <= 16'b0000_0000_0000_0000;
array[15000] <= 16'b0000_0000_0000_0000;
array[15001] <= 16'b0000_0000_0000_0000;
array[15002] <= 16'b0000_0000_0000_0000;
array[15003] <= 16'b0000_0000_0000_0000;
array[15004] <= 16'b0000_0000_0000_0000;
array[15005] <= 16'b0000_0000_0000_0000;
array[15006] <= 16'b0000_0000_0000_0000;
array[15007] <= 16'b0000_0000_0000_0000;
array[15008] <= 16'b0000_0000_0000_0000;
array[15009] <= 16'b0000_0000_0000_0000;
array[15010] <= 16'b0000_0000_0000_0000;
array[15011] <= 16'b0000_0000_0000_0000;
array[15012] <= 16'b0000_0000_0000_0000;
array[15013] <= 16'b0000_0000_0000_0000;
array[15014] <= 16'b0000_0000_0000_0000;
array[15015] <= 16'b0000_0000_0000_0000;
array[15016] <= 16'b0000_0000_0000_0000;
array[15017] <= 16'b0000_0000_0000_0000;
array[15018] <= 16'b0000_0000_0000_0000;
array[15019] <= 16'b0000_0000_0000_0000;
array[15020] <= 16'b0000_0000_0000_0000;
array[15021] <= 16'b0000_0000_0000_0000;
array[15022] <= 16'b0000_0000_0000_0000;
array[15023] <= 16'b0000_0000_0000_0000;
array[15024] <= 16'b0000_0000_0000_0000;
array[15025] <= 16'b0000_0000_0000_0000;
array[15026] <= 16'b0000_0000_0000_0000;
array[15027] <= 16'b0000_0000_0000_0000;
array[15028] <= 16'b0000_0000_0000_0000;
array[15029] <= 16'b0000_0000_0000_0000;
array[15030] <= 16'b0000_0000_0000_0000;
array[15031] <= 16'b0000_0000_0000_0000;
array[15032] <= 16'b0000_0000_0000_0000;
array[15033] <= 16'b0000_0000_0000_0000;
array[15034] <= 16'b0000_0000_0000_0000;
array[15035] <= 16'b0000_0000_0000_0000;
array[15036] <= 16'b0000_0000_0000_0000;
array[15037] <= 16'b0000_0000_0000_0000;
array[15038] <= 16'b0000_0000_0000_0000;
array[15039] <= 16'b0000_0000_0000_0000;
array[15040] <= 16'b0000_0000_0000_0000;
array[15041] <= 16'b0000_0000_0000_0000;
array[15042] <= 16'b0000_0000_0000_0000;
array[15043] <= 16'b0000_0000_0000_0000;
array[15044] <= 16'b0000_0000_0000_0000;
array[15045] <= 16'b0000_0000_0000_0000;
array[15046] <= 16'b0000_0000_0000_0000;
array[15047] <= 16'b0000_0000_0000_0000;
array[15048] <= 16'b0000_0000_0000_0000;
array[15049] <= 16'b0000_0000_0000_0000;
array[15050] <= 16'b0000_0000_0000_0000;
array[15051] <= 16'b0000_0000_0000_0000;
array[15052] <= 16'b0000_0000_0000_0000;
array[15053] <= 16'b0000_0000_0000_0000;
array[15054] <= 16'b0000_0000_0000_0000;
array[15055] <= 16'b0000_0000_0000_0000;
array[15056] <= 16'b0000_0000_0000_0000;
array[15057] <= 16'b0000_0000_0000_0000;
array[15058] <= 16'b0000_0000_0000_0000;
array[15059] <= 16'b0000_0000_0000_0000;
array[15060] <= 16'b0000_0000_0000_0000;
array[15061] <= 16'b0000_0000_0000_0000;
array[15062] <= 16'b0000_0000_0000_0000;
array[15063] <= 16'b0000_0000_0000_0000;
array[15064] <= 16'b0000_0000_0000_0000;
array[15065] <= 16'b0000_0000_0000_0000;
array[15066] <= 16'b0000_0000_0000_0000;
array[15067] <= 16'b0000_0000_0000_0000;
array[15068] <= 16'b0000_0000_0000_0000;
array[15069] <= 16'b0000_0000_0000_0000;
array[15070] <= 16'b0000_0000_0000_0000;
array[15071] <= 16'b0000_0000_0000_0000;
array[15072] <= 16'b0000_0000_0000_0000;
array[15073] <= 16'b0000_0000_0000_0000;
array[15074] <= 16'b0000_0000_0000_0000;
array[15075] <= 16'b0000_0000_0000_0000;
array[15076] <= 16'b0000_0000_0000_0000;
array[15077] <= 16'b0000_0000_0000_0000;
array[15078] <= 16'b0000_0000_0000_0000;
array[15079] <= 16'b0000_0000_0000_0000;
array[15080] <= 16'b0000_0000_0000_0000;
array[15081] <= 16'b0000_0000_0000_0000;
array[15082] <= 16'b0000_0000_0000_0000;
array[15083] <= 16'b0000_0000_0000_0000;
array[15084] <= 16'b0000_0000_0000_0000;
array[15085] <= 16'b0000_0000_0000_0000;
array[15086] <= 16'b0000_0000_0000_0000;
array[15087] <= 16'b0000_0000_0000_0000;
array[15088] <= 16'b0000_0000_0000_0000;
array[15089] <= 16'b0000_0000_0000_0000;
array[15090] <= 16'b0000_0000_0000_0000;
array[15091] <= 16'b0000_0000_0000_0000;
array[15092] <= 16'b0000_0000_0000_0000;
array[15093] <= 16'b0000_0000_0000_0000;
array[15094] <= 16'b0000_0000_0000_0000;
array[15095] <= 16'b0000_0000_0000_0000;
array[15096] <= 16'b0000_0000_0000_0000;
array[15097] <= 16'b0000_0000_0000_0000;
array[15098] <= 16'b0000_0000_0000_0000;
array[15099] <= 16'b0000_0000_0000_0000;
array[15100] <= 16'b0000_0000_0000_0000;
array[15101] <= 16'b0000_0000_0000_0000;
array[15102] <= 16'b0000_0000_0000_0000;
array[15103] <= 16'b0000_0000_0000_0000;
array[15104] <= 16'b0000_0000_0000_0000;
array[15105] <= 16'b0000_0000_0000_0000;
array[15106] <= 16'b0000_0000_0000_0000;
array[15107] <= 16'b0000_0000_0000_0000;
array[15108] <= 16'b0000_0000_0000_0000;
array[15109] <= 16'b0000_0000_0000_0000;
array[15110] <= 16'b0000_0000_0000_0000;
array[15111] <= 16'b0000_0000_0000_0000;
array[15112] <= 16'b0000_0000_0000_0000;
array[15113] <= 16'b0000_0000_0000_0000;
array[15114] <= 16'b0000_0000_0000_0000;
array[15115] <= 16'b0000_0000_0000_0000;
array[15116] <= 16'b0000_0000_0000_0000;
array[15117] <= 16'b0000_0000_0000_0000;
array[15118] <= 16'b0000_0000_0000_0000;
array[15119] <= 16'b0000_0000_0000_0000;
array[15120] <= 16'b0000_0000_0000_0000;
array[15121] <= 16'b0000_0000_0000_0000;
array[15122] <= 16'b0000_0000_0000_0000;
array[15123] <= 16'b0000_0000_0000_0000;
array[15124] <= 16'b0000_0000_0000_0000;
array[15125] <= 16'b0000_0000_0000_0000;
array[15126] <= 16'b0000_0000_0000_0000;
array[15127] <= 16'b0000_0000_0000_0000;
array[15128] <= 16'b0000_0000_0000_0000;
array[15129] <= 16'b0000_0000_0000_0000;
array[15130] <= 16'b0000_0000_0000_0000;
array[15131] <= 16'b0000_0000_0000_0000;
array[15132] <= 16'b0000_0000_0000_0000;
array[15133] <= 16'b0000_0000_0000_0000;
array[15134] <= 16'b0000_0000_0000_0000;
array[15135] <= 16'b0000_0000_0000_0000;
array[15136] <= 16'b0000_0000_0000_0000;
array[15137] <= 16'b0000_0000_0000_0000;
array[15138] <= 16'b0000_0000_0000_0000;
array[15139] <= 16'b0000_0000_0000_0000;
array[15140] <= 16'b0000_0000_0000_0000;
array[15141] <= 16'b0000_0000_0000_0000;
array[15142] <= 16'b0000_0000_0000_0000;
array[15143] <= 16'b0000_0000_0000_0000;
array[15144] <= 16'b0000_0000_0000_0000;
array[15145] <= 16'b0000_0000_0000_0000;
array[15146] <= 16'b0000_0000_0000_0000;
array[15147] <= 16'b0000_0000_0000_0000;
array[15148] <= 16'b0000_0000_0000_0000;
array[15149] <= 16'b0000_0000_0000_0000;
array[15150] <= 16'b0000_0000_0000_0000;
array[15151] <= 16'b0000_0000_0000_0000;
array[15152] <= 16'b0000_0000_0000_0000;
array[15153] <= 16'b0000_0000_0000_0000;
array[15154] <= 16'b0000_0000_0000_0000;
array[15155] <= 16'b0000_0000_0000_0000;
array[15156] <= 16'b0000_0000_0000_0000;
array[15157] <= 16'b0000_0000_0000_0000;
array[15158] <= 16'b0000_0000_0000_0000;
array[15159] <= 16'b0000_0000_0000_0000;
array[15160] <= 16'b0000_0000_0000_0000;
array[15161] <= 16'b0000_0000_0000_0000;
array[15162] <= 16'b0000_0000_0000_0000;
array[15163] <= 16'b0000_0000_0000_0000;
array[15164] <= 16'b0000_0000_0000_0000;
array[15165] <= 16'b0000_0000_0000_0000;
array[15166] <= 16'b0000_0000_0000_0000;
array[15167] <= 16'b0000_0000_0000_0000;
array[15168] <= 16'b0000_0000_0000_0000;
array[15169] <= 16'b0000_0000_0000_0000;
array[15170] <= 16'b0000_0000_0000_0000;
array[15171] <= 16'b0000_0000_0000_0000;
array[15172] <= 16'b0000_0000_0000_0000;
array[15173] <= 16'b0000_0000_0000_0000;
array[15174] <= 16'b0000_0000_0000_0000;
array[15175] <= 16'b0000_0000_0000_0000;
array[15176] <= 16'b0000_0000_0000_0000;
array[15177] <= 16'b0000_0000_0000_0000;
array[15178] <= 16'b0000_0000_0000_0000;
array[15179] <= 16'b0000_0000_0000_0000;
array[15180] <= 16'b0000_0000_0000_0000;
array[15181] <= 16'b0000_0000_0000_0000;
array[15182] <= 16'b0000_0000_0000_0000;
array[15183] <= 16'b0000_0000_0000_0000;
array[15184] <= 16'b0000_0000_0000_0000;
array[15185] <= 16'b0000_0000_0000_0000;
array[15186] <= 16'b0000_0000_0000_0000;
array[15187] <= 16'b0000_0000_0000_0000;
array[15188] <= 16'b0000_0000_0000_0000;
array[15189] <= 16'b0000_0000_0000_0000;
array[15190] <= 16'b0000_0000_0000_0000;
array[15191] <= 16'b0000_0000_0000_0000;
array[15192] <= 16'b0000_0000_0000_0000;
array[15193] <= 16'b0000_0000_0000_0000;
array[15194] <= 16'b0000_0000_0000_0000;
array[15195] <= 16'b0000_0000_0000_0000;
array[15196] <= 16'b0000_0000_0000_0000;
array[15197] <= 16'b0000_0000_0000_0000;
array[15198] <= 16'b0000_0000_0000_0000;
array[15199] <= 16'b0000_0000_0000_0000;
array[15200] <= 16'b0000_0000_0000_0000;
array[15201] <= 16'b0000_0000_0000_0000;
array[15202] <= 16'b0000_0000_0000_0000;
array[15203] <= 16'b0000_0000_0000_0000;
array[15204] <= 16'b0000_0000_0000_0000;
array[15205] <= 16'b0000_0000_0000_0000;
array[15206] <= 16'b0000_0000_0000_0000;
array[15207] <= 16'b0000_0000_0000_0000;
array[15208] <= 16'b0000_0000_0000_0000;
array[15209] <= 16'b0000_0000_0000_0000;
array[15210] <= 16'b0000_0000_0000_0000;
array[15211] <= 16'b0000_0000_0000_0000;
array[15212] <= 16'b0000_0000_0000_0000;
array[15213] <= 16'b0000_0000_0000_0000;
array[15214] <= 16'b0000_0000_0000_0000;
array[15215] <= 16'b0000_0000_0000_0000;
array[15216] <= 16'b0000_0000_0000_0000;
array[15217] <= 16'b0000_0000_0000_0000;
array[15218] <= 16'b0000_0000_0000_0000;
array[15219] <= 16'b0000_0000_0000_0000;
array[15220] <= 16'b0000_0000_0000_0000;
array[15221] <= 16'b0000_0000_0000_0000;
array[15222] <= 16'b0000_0000_0000_0000;
array[15223] <= 16'b0000_0000_0000_0000;
array[15224] <= 16'b0000_0000_0000_0000;
array[15225] <= 16'b0000_0000_0000_0000;
array[15226] <= 16'b0000_0000_0000_0000;
array[15227] <= 16'b0000_0000_0000_0000;
array[15228] <= 16'b0000_0000_0000_0000;
array[15229] <= 16'b0000_0000_0000_0000;
array[15230] <= 16'b0000_0000_0000_0000;
array[15231] <= 16'b0000_0000_0000_0000;
array[15232] <= 16'b0000_0000_0000_0000;
array[15233] <= 16'b0000_0000_0000_0000;
array[15234] <= 16'b0000_0000_0000_0000;
array[15235] <= 16'b0000_0000_0000_0000;
array[15236] <= 16'b0000_0000_0000_0000;
array[15237] <= 16'b0000_0000_0000_0000;
array[15238] <= 16'b0000_0000_0000_0000;
array[15239] <= 16'b0000_0000_0000_0000;
array[15240] <= 16'b0000_0000_0000_0000;
array[15241] <= 16'b0000_0000_0000_0000;
array[15242] <= 16'b0000_0000_0000_0000;
array[15243] <= 16'b0000_0000_0000_0000;
array[15244] <= 16'b0000_0000_0000_0000;
array[15245] <= 16'b0000_0000_0000_0000;
array[15246] <= 16'b0000_0000_0000_0000;
array[15247] <= 16'b0000_0000_0000_0000;
array[15248] <= 16'b0000_0000_0000_0000;
array[15249] <= 16'b0000_0000_0000_0000;
array[15250] <= 16'b0000_0000_0000_0000;
array[15251] <= 16'b0000_0000_0000_0000;
array[15252] <= 16'b0000_0000_0000_0000;
array[15253] <= 16'b0000_0000_0000_0000;
array[15254] <= 16'b0000_0000_0000_0000;
array[15255] <= 16'b0000_0000_0000_0000;
array[15256] <= 16'b0000_0000_0000_0000;
array[15257] <= 16'b0000_0000_0000_0000;
array[15258] <= 16'b0000_0000_0000_0000;
array[15259] <= 16'b0000_0000_0000_0000;
array[15260] <= 16'b0000_0000_0000_0000;
array[15261] <= 16'b0000_0000_0000_0000;
array[15262] <= 16'b0000_0000_0000_0000;
array[15263] <= 16'b0000_0000_0000_0000;
array[15264] <= 16'b0000_0000_0000_0000;
array[15265] <= 16'b0000_0000_0000_0000;
array[15266] <= 16'b0000_0000_0000_0000;
array[15267] <= 16'b0000_0000_0000_0000;
array[15268] <= 16'b0000_0000_0000_0000;
array[15269] <= 16'b0000_0000_0000_0000;
array[15270] <= 16'b0000_0000_0000_0000;
array[15271] <= 16'b0000_0000_0000_0000;
array[15272] <= 16'b0000_0000_0000_0000;
array[15273] <= 16'b0000_0000_0000_0000;
array[15274] <= 16'b0000_0000_0000_0000;
array[15275] <= 16'b0000_0000_0000_0000;
array[15276] <= 16'b0000_0000_0000_0000;
array[15277] <= 16'b0000_0000_0000_0000;
array[15278] <= 16'b0000_0000_0000_0000;
array[15279] <= 16'b0000_0000_0000_0000;
array[15280] <= 16'b0000_0000_0000_0000;
array[15281] <= 16'b0000_0000_0000_0000;
array[15282] <= 16'b0000_0000_0000_0000;
array[15283] <= 16'b0000_0000_0000_0000;
array[15284] <= 16'b0000_0000_0000_0000;
array[15285] <= 16'b0000_0000_0000_0000;
array[15286] <= 16'b0000_0000_0000_0000;
array[15287] <= 16'b0000_0000_0000_0000;
array[15288] <= 16'b0000_0000_0000_0000;
array[15289] <= 16'b0000_0000_0000_0000;
array[15290] <= 16'b0000_0000_0000_0000;
array[15291] <= 16'b0000_0000_0000_0000;
array[15292] <= 16'b0000_0000_0000_0000;
array[15293] <= 16'b0000_0000_0000_0000;
array[15294] <= 16'b0000_0000_0000_0000;
array[15295] <= 16'b0000_0000_0000_0000;
array[15296] <= 16'b0000_0000_0000_0000;
array[15297] <= 16'b0000_0000_0000_0000;
array[15298] <= 16'b0000_0000_0000_0000;
array[15299] <= 16'b0000_0000_0000_0000;
array[15300] <= 16'b0000_0000_0000_0000;
array[15301] <= 16'b0000_0000_0000_0000;
array[15302] <= 16'b0000_0000_0000_0000;
array[15303] <= 16'b0000_0000_0000_0000;
array[15304] <= 16'b0000_0000_0000_0000;
array[15305] <= 16'b0000_0000_0000_0000;
array[15306] <= 16'b0000_0000_0000_0000;
array[15307] <= 16'b0000_0000_0000_0000;
array[15308] <= 16'b0000_0000_0000_0000;
array[15309] <= 16'b0000_0000_0000_0000;
array[15310] <= 16'b0000_0000_0000_0000;
array[15311] <= 16'b0000_0000_0000_0000;
array[15312] <= 16'b0000_0000_0000_0000;
array[15313] <= 16'b0000_0000_0000_0000;
array[15314] <= 16'b0000_0000_0000_0000;
array[15315] <= 16'b0000_0000_0000_0000;
array[15316] <= 16'b0000_0000_0000_0000;
array[15317] <= 16'b0000_0000_0000_0000;
array[15318] <= 16'b0000_0000_0000_0000;
array[15319] <= 16'b0000_0000_0000_0000;
array[15320] <= 16'b0000_0000_0000_0000;
array[15321] <= 16'b0000_0000_0000_0000;
array[15322] <= 16'b0000_0000_0000_0000;
array[15323] <= 16'b0000_0000_0000_0000;
array[15324] <= 16'b0000_0000_0000_0000;
array[15325] <= 16'b0000_0000_0000_0000;
array[15326] <= 16'b0000_0000_0000_0000;
array[15327] <= 16'b0000_0000_0000_0000;
array[15328] <= 16'b0000_0000_0000_0000;
array[15329] <= 16'b0000_0000_0000_0000;
array[15330] <= 16'b0000_0000_0000_0000;
array[15331] <= 16'b0000_0000_0000_0000;
array[15332] <= 16'b0000_0000_0000_0000;
array[15333] <= 16'b0000_0000_0000_0000;
array[15334] <= 16'b0000_0000_0000_0000;
array[15335] <= 16'b0000_0000_0000_0000;
array[15336] <= 16'b0000_0000_0000_0000;
array[15337] <= 16'b0000_0000_0000_0000;
array[15338] <= 16'b0000_0000_0000_0000;
array[15339] <= 16'b0000_0000_0000_0000;
array[15340] <= 16'b0000_0000_0000_0000;
array[15341] <= 16'b0000_0000_0000_0000;
array[15342] <= 16'b0000_0000_0000_0000;
array[15343] <= 16'b0000_0000_0000_0000;
array[15344] <= 16'b0000_0000_0000_0000;
array[15345] <= 16'b0000_0000_0000_0000;
array[15346] <= 16'b0000_0000_0000_0000;
array[15347] <= 16'b0000_0000_0000_0000;
array[15348] <= 16'b0000_0000_0000_0000;
array[15349] <= 16'b0000_0000_0000_0000;
array[15350] <= 16'b0000_0000_0000_0000;
array[15351] <= 16'b0000_0000_0000_0000;
array[15352] <= 16'b0000_0000_0000_0000;
array[15353] <= 16'b0000_0000_0000_0000;
array[15354] <= 16'b0000_0000_0000_0000;
array[15355] <= 16'b0000_0000_0000_0000;
array[15356] <= 16'b0000_0000_0000_0000;
array[15357] <= 16'b0000_0000_0000_0000;
array[15358] <= 16'b0000_0000_0000_0000;
array[15359] <= 16'b0000_0000_0000_0000;
array[15360] <= 16'b0000_0000_0000_0000;
array[15361] <= 16'b0000_0000_0000_0000;
array[15362] <= 16'b0000_0000_0000_0000;
array[15363] <= 16'b0000_0000_0000_0000;
array[15364] <= 16'b0000_0000_0000_0000;
array[15365] <= 16'b0000_0000_0000_0000;
array[15366] <= 16'b0000_0000_0000_0000;
array[15367] <= 16'b0000_0000_0000_0000;
array[15368] <= 16'b0000_0000_0000_0000;
array[15369] <= 16'b0000_0000_0000_0000;
array[15370] <= 16'b0000_0000_0000_0000;
array[15371] <= 16'b0000_0000_0000_0000;
array[15372] <= 16'b0000_0000_0000_0000;
array[15373] <= 16'b0000_0000_0000_0000;
array[15374] <= 16'b0000_0000_0000_0000;
array[15375] <= 16'b0000_0000_0000_0000;
array[15376] <= 16'b0000_0000_0000_0000;
array[15377] <= 16'b0000_0000_0000_0000;
array[15378] <= 16'b0000_0000_0000_0000;
array[15379] <= 16'b0000_0000_0000_0000;
array[15380] <= 16'b0000_0000_0000_0000;
array[15381] <= 16'b0000_0000_0000_0000;
array[15382] <= 16'b0000_0000_0000_0000;
array[15383] <= 16'b0000_0000_0000_0000;
array[15384] <= 16'b0000_0000_0000_0000;
array[15385] <= 16'b0000_0000_0000_0000;
array[15386] <= 16'b0000_0000_0000_0000;
array[15387] <= 16'b0000_0000_0000_0000;
array[15388] <= 16'b0000_0000_0000_0000;
array[15389] <= 16'b0000_0000_0000_0000;
array[15390] <= 16'b0000_0000_0000_0000;
array[15391] <= 16'b0000_0000_0000_0000;
array[15392] <= 16'b0000_0000_0000_0000;
array[15393] <= 16'b0000_0000_0000_0000;
array[15394] <= 16'b0000_0000_0000_0000;
array[15395] <= 16'b0000_0000_0000_0000;
array[15396] <= 16'b0000_0000_0000_0000;
array[15397] <= 16'b0000_0000_0000_0000;
array[15398] <= 16'b0000_0000_0000_0000;
array[15399] <= 16'b0000_0000_0000_0000;
array[15400] <= 16'b0000_0000_0000_0000;
array[15401] <= 16'b0000_0000_0000_0000;
array[15402] <= 16'b0000_0000_0000_0000;
array[15403] <= 16'b0000_0000_0000_0000;
array[15404] <= 16'b0000_0000_0000_0000;
array[15405] <= 16'b0000_0000_0000_0000;
array[15406] <= 16'b0000_0000_0000_0000;
array[15407] <= 16'b0000_0000_0000_0000;
array[15408] <= 16'b0000_0000_0000_0000;
array[15409] <= 16'b0000_0000_0000_0000;
array[15410] <= 16'b0000_0000_0000_0000;
array[15411] <= 16'b0000_0000_0000_0000;
array[15412] <= 16'b0000_0000_0000_0000;
array[15413] <= 16'b0000_0000_0000_0000;
array[15414] <= 16'b0000_0000_0000_0000;
array[15415] <= 16'b0000_0000_0000_0000;
array[15416] <= 16'b0000_0000_0000_0000;
array[15417] <= 16'b0000_0000_0000_0000;
array[15418] <= 16'b0000_0000_0000_0000;
array[15419] <= 16'b0000_0000_0000_0000;
array[15420] <= 16'b0000_0000_0000_0000;
array[15421] <= 16'b0000_0000_0000_0000;
array[15422] <= 16'b0000_0000_0000_0000;
array[15423] <= 16'b0000_0000_0000_0000;
array[15424] <= 16'b0000_0000_0000_0000;
array[15425] <= 16'b0000_0000_0000_0000;
array[15426] <= 16'b0000_0000_0000_0000;
array[15427] <= 16'b0000_0000_0000_0000;
array[15428] <= 16'b0000_0000_0000_0000;
array[15429] <= 16'b0000_0000_0000_0000;
array[15430] <= 16'b0000_0000_0000_0000;
array[15431] <= 16'b0000_0000_0000_0000;
array[15432] <= 16'b0000_0000_0000_0000;
array[15433] <= 16'b0000_0000_0000_0000;
array[15434] <= 16'b0000_0000_0000_0000;
array[15435] <= 16'b0000_0000_0000_0000;
array[15436] <= 16'b0000_0000_0000_0000;
array[15437] <= 16'b0000_0000_0000_0000;
array[15438] <= 16'b0000_0000_0000_0000;
array[15439] <= 16'b0000_0000_0000_0000;
array[15440] <= 16'b0000_0000_0000_0000;
array[15441] <= 16'b0000_0000_0000_0000;
array[15442] <= 16'b0000_0000_0000_0000;
array[15443] <= 16'b0000_0000_0000_0000;
array[15444] <= 16'b0000_0000_0000_0000;
array[15445] <= 16'b0000_0000_0000_0000;
array[15446] <= 16'b0000_0000_0000_0000;
array[15447] <= 16'b0000_0000_0000_0000;
array[15448] <= 16'b0000_0000_0000_0000;
array[15449] <= 16'b0000_0000_0000_0000;
array[15450] <= 16'b0000_0000_0000_0000;
array[15451] <= 16'b0000_0000_0000_0000;
array[15452] <= 16'b0000_0000_0000_0000;
array[15453] <= 16'b0000_0000_0000_0000;
array[15454] <= 16'b0000_0000_0000_0000;
array[15455] <= 16'b0000_0000_0000_0000;
array[15456] <= 16'b0000_0000_0000_0000;
array[15457] <= 16'b0000_0000_0000_0000;
array[15458] <= 16'b0000_0000_0000_0000;
array[15459] <= 16'b0000_0000_0000_0000;
array[15460] <= 16'b0000_0000_0000_0000;
array[15461] <= 16'b0000_0000_0000_0000;
array[15462] <= 16'b0000_0000_0000_0000;
array[15463] <= 16'b0000_0000_0000_0000;
array[15464] <= 16'b0000_0000_0000_0000;
array[15465] <= 16'b0000_0000_0000_0000;
array[15466] <= 16'b0000_0000_0000_0000;
array[15467] <= 16'b0000_0000_0000_0000;
array[15468] <= 16'b0000_0000_0000_0000;
array[15469] <= 16'b0000_0000_0000_0000;
array[15470] <= 16'b0000_0000_0000_0000;
array[15471] <= 16'b0000_0000_0000_0000;
array[15472] <= 16'b0000_0000_0000_0000;
array[15473] <= 16'b0000_0000_0000_0000;
array[15474] <= 16'b0000_0000_0000_0000;
array[15475] <= 16'b0000_0000_0000_0000;
array[15476] <= 16'b0000_0000_0000_0000;
array[15477] <= 16'b0000_0000_0000_0000;
array[15478] <= 16'b0000_0000_0000_0000;
array[15479] <= 16'b0000_0000_0000_0000;
array[15480] <= 16'b0000_0000_0000_0000;
array[15481] <= 16'b0000_0000_0000_0000;
array[15482] <= 16'b0000_0000_0000_0000;
array[15483] <= 16'b0000_0000_0000_0000;
array[15484] <= 16'b0000_0000_0000_0000;
array[15485] <= 16'b0000_0000_0000_0000;
array[15486] <= 16'b0000_0000_0000_0000;
array[15487] <= 16'b0000_0000_0000_0000;
array[15488] <= 16'b0000_0000_0000_0000;
array[15489] <= 16'b0000_0000_0000_0000;
array[15490] <= 16'b0000_0000_0000_0000;
array[15491] <= 16'b0000_0000_0000_0000;
array[15492] <= 16'b0000_0000_0000_0000;
array[15493] <= 16'b0000_0000_0000_0000;
array[15494] <= 16'b0000_0000_0000_0000;
array[15495] <= 16'b0000_0000_0000_0000;
array[15496] <= 16'b0000_0000_0000_0000;
array[15497] <= 16'b0000_0000_0000_0000;
array[15498] <= 16'b0000_0000_0000_0000;
array[15499] <= 16'b0000_0000_0000_0000;
array[15500] <= 16'b0000_0000_0000_0000;
array[15501] <= 16'b0000_0000_0000_0000;
array[15502] <= 16'b0000_0000_0000_0000;
array[15503] <= 16'b0000_0000_0000_0000;
array[15504] <= 16'b0000_0000_0000_0000;
array[15505] <= 16'b0000_0000_0000_0000;
array[15506] <= 16'b0000_0000_0000_0000;
array[15507] <= 16'b0000_0000_0000_0000;
array[15508] <= 16'b0000_0000_0000_0000;
array[15509] <= 16'b0000_0000_0000_0000;
array[15510] <= 16'b0000_0000_0000_0000;
array[15511] <= 16'b0000_0000_0000_0000;
array[15512] <= 16'b0000_0000_0000_0000;
array[15513] <= 16'b0000_0000_0000_0000;
array[15514] <= 16'b0000_0000_0000_0000;
array[15515] <= 16'b0000_0000_0000_0000;
array[15516] <= 16'b0000_0000_0000_0000;
array[15517] <= 16'b0000_0000_0000_0000;
array[15518] <= 16'b0000_0000_0000_0000;
array[15519] <= 16'b0000_0000_0000_0000;
array[15520] <= 16'b0000_0000_0000_0000;
array[15521] <= 16'b0000_0000_0000_0000;
array[15522] <= 16'b0000_0000_0000_0000;
array[15523] <= 16'b0000_0000_0000_0000;
array[15524] <= 16'b0000_0000_0000_0000;
array[15525] <= 16'b0000_0000_0000_0000;
array[15526] <= 16'b0000_0000_0000_0000;
array[15527] <= 16'b0000_0000_0000_0000;
array[15528] <= 16'b0000_0000_0000_0000;
array[15529] <= 16'b0000_0000_0000_0000;
array[15530] <= 16'b0000_0000_0000_0000;
array[15531] <= 16'b0000_0000_0000_0000;
array[15532] <= 16'b0000_0000_0000_0000;
array[15533] <= 16'b0000_0000_0000_0000;
array[15534] <= 16'b0000_0000_0000_0000;
array[15535] <= 16'b0000_0000_0000_0000;
array[15536] <= 16'b0000_0000_0000_0000;
array[15537] <= 16'b0000_0000_0000_0000;
array[15538] <= 16'b0000_0000_0000_0000;
array[15539] <= 16'b0000_0000_0000_0000;
array[15540] <= 16'b0000_0000_0000_0000;
array[15541] <= 16'b0000_0000_0000_0000;
array[15542] <= 16'b0000_0000_0000_0000;
array[15543] <= 16'b0000_0000_0000_0000;
array[15544] <= 16'b0000_0000_0000_0000;
array[15545] <= 16'b0000_0000_0000_0000;
array[15546] <= 16'b0000_0000_0000_0000;
array[15547] <= 16'b0000_0000_0000_0000;
array[15548] <= 16'b0000_0000_0000_0000;
array[15549] <= 16'b0000_0000_0000_0000;
array[15550] <= 16'b0000_0000_0000_0000;
array[15551] <= 16'b0000_0000_0000_0000;
array[15552] <= 16'b0000_0000_0000_0000;
array[15553] <= 16'b0000_0000_0000_0000;
array[15554] <= 16'b0000_0000_0000_0000;
array[15555] <= 16'b0000_0000_0000_0000;
array[15556] <= 16'b0000_0000_0000_0000;
array[15557] <= 16'b0000_0000_0000_0000;
array[15558] <= 16'b0000_0000_0000_0000;
array[15559] <= 16'b0000_0000_0000_0000;
array[15560] <= 16'b0000_0000_0000_0000;
array[15561] <= 16'b0000_0000_0000_0000;
array[15562] <= 16'b0000_0000_0000_0000;
array[15563] <= 16'b0000_0000_0000_0000;
array[15564] <= 16'b0000_0000_0000_0000;
array[15565] <= 16'b0000_0000_0000_0000;
array[15566] <= 16'b0000_0000_0000_0000;
array[15567] <= 16'b0000_0000_0000_0000;
array[15568] <= 16'b0000_0000_0000_0000;
array[15569] <= 16'b0000_0000_0000_0000;
array[15570] <= 16'b0000_0000_0000_0000;
array[15571] <= 16'b0000_0000_0000_0000;
array[15572] <= 16'b0000_0000_0000_0000;
array[15573] <= 16'b0000_0000_0000_0000;
array[15574] <= 16'b0000_0000_0000_0000;
array[15575] <= 16'b0000_0000_0000_0000;
array[15576] <= 16'b0000_0000_0000_0000;
array[15577] <= 16'b0000_0000_0000_0000;
array[15578] <= 16'b0000_0000_0000_0000;
array[15579] <= 16'b0000_0000_0000_0000;
array[15580] <= 16'b0000_0000_0000_0000;
array[15581] <= 16'b0000_0000_0000_0000;
array[15582] <= 16'b0000_0000_0000_0000;
array[15583] <= 16'b0000_0000_0000_0000;
array[15584] <= 16'b0000_0000_0000_0000;
array[15585] <= 16'b0000_0000_0000_0000;
array[15586] <= 16'b0000_0000_0000_0000;
array[15587] <= 16'b0000_0000_0000_0000;
array[15588] <= 16'b0000_0000_0000_0000;
array[15589] <= 16'b0000_0000_0000_0000;
array[15590] <= 16'b0000_0000_0000_0000;
array[15591] <= 16'b0000_0000_0000_0000;
array[15592] <= 16'b0000_0000_0000_0000;
array[15593] <= 16'b0000_0000_0000_0000;
array[15594] <= 16'b0000_0000_0000_0000;
array[15595] <= 16'b0000_0000_0000_0000;
array[15596] <= 16'b0000_0000_0000_0000;
array[15597] <= 16'b0000_0000_0000_0000;
array[15598] <= 16'b0000_0000_0000_0000;
array[15599] <= 16'b0000_0000_0000_0000;
array[15600] <= 16'b0000_0000_0000_0000;
array[15601] <= 16'b0000_0000_0000_0000;
array[15602] <= 16'b0000_0000_0000_0000;
array[15603] <= 16'b0000_0000_0000_0000;
array[15604] <= 16'b0000_0000_0000_0000;
array[15605] <= 16'b0000_0000_0000_0000;
array[15606] <= 16'b0000_0000_0000_0000;
array[15607] <= 16'b0000_0000_0000_0000;
array[15608] <= 16'b0000_0000_0000_0000;
array[15609] <= 16'b0000_0000_0000_0000;
array[15610] <= 16'b0000_0000_0000_0000;
array[15611] <= 16'b0000_0000_0000_0000;
array[15612] <= 16'b0000_0000_0000_0000;
array[15613] <= 16'b0000_0000_0000_0000;
array[15614] <= 16'b0000_0000_0000_0000;
array[15615] <= 16'b0000_0000_0000_0000;
array[15616] <= 16'b0000_0000_0000_0000;
array[15617] <= 16'b0000_0000_0000_0000;
array[15618] <= 16'b0000_0000_0000_0000;
array[15619] <= 16'b0000_0000_0000_0000;
array[15620] <= 16'b0000_0000_0000_0000;
array[15621] <= 16'b0000_0000_0000_0000;
array[15622] <= 16'b0000_0000_0000_0000;
array[15623] <= 16'b0000_0000_0000_0000;
array[15624] <= 16'b0000_0000_0000_0000;
array[15625] <= 16'b0000_0000_0000_0000;
array[15626] <= 16'b0000_0000_0000_0000;
array[15627] <= 16'b0000_0000_0000_0000;
array[15628] <= 16'b0000_0000_0000_0000;
array[15629] <= 16'b0000_0000_0000_0000;
array[15630] <= 16'b0000_0000_0000_0000;
array[15631] <= 16'b0000_0000_0000_0000;
array[15632] <= 16'b0000_0000_0000_0000;
array[15633] <= 16'b0000_0000_0000_0000;
array[15634] <= 16'b0000_0000_0000_0000;
array[15635] <= 16'b0000_0000_0000_0000;
array[15636] <= 16'b0000_0000_0000_0000;
array[15637] <= 16'b0000_0000_0000_0000;
array[15638] <= 16'b0000_0000_0000_0000;
array[15639] <= 16'b0000_0000_0000_0000;
array[15640] <= 16'b0000_0000_0000_0000;
array[15641] <= 16'b0000_0000_0000_0000;
array[15642] <= 16'b0000_0000_0000_0000;
array[15643] <= 16'b0000_0000_0000_0000;
array[15644] <= 16'b0000_0000_0000_0000;
array[15645] <= 16'b0000_0000_0000_0000;
array[15646] <= 16'b0000_0000_0000_0000;
array[15647] <= 16'b0000_0000_0000_0000;
array[15648] <= 16'b0000_0000_0000_0000;
array[15649] <= 16'b0000_0000_0000_0000;
array[15650] <= 16'b0000_0000_0000_0000;
array[15651] <= 16'b0000_0000_0000_0000;
array[15652] <= 16'b0000_0000_0000_0000;
array[15653] <= 16'b0000_0000_0000_0000;
array[15654] <= 16'b0000_0000_0000_0000;
array[15655] <= 16'b0000_0000_0000_0000;
array[15656] <= 16'b0000_0000_0000_0000;
array[15657] <= 16'b0000_0000_0000_0000;
array[15658] <= 16'b0000_0000_0000_0000;
array[15659] <= 16'b0000_0000_0000_0000;
array[15660] <= 16'b0000_0000_0000_0000;
array[15661] <= 16'b0000_0000_0000_0000;
array[15662] <= 16'b0000_0000_0000_0000;
array[15663] <= 16'b0000_0000_0000_0000;
array[15664] <= 16'b0000_0000_0000_0000;
array[15665] <= 16'b0000_0000_0000_0000;
array[15666] <= 16'b0000_0000_0000_0000;
array[15667] <= 16'b0000_0000_0000_0000;
array[15668] <= 16'b0000_0000_0000_0000;
array[15669] <= 16'b0000_0000_0000_0000;
array[15670] <= 16'b0000_0000_0000_0000;
array[15671] <= 16'b0000_0000_0000_0000;
array[15672] <= 16'b0000_0000_0000_0000;
array[15673] <= 16'b0000_0000_0000_0000;
array[15674] <= 16'b0000_0000_0000_0000;
array[15675] <= 16'b0000_0000_0000_0000;
array[15676] <= 16'b0000_0000_0000_0000;
array[15677] <= 16'b0000_0000_0000_0000;
array[15678] <= 16'b0000_0000_0000_0000;
array[15679] <= 16'b0000_0000_0000_0000;
array[15680] <= 16'b0000_0000_0000_0000;
array[15681] <= 16'b0000_0000_0000_0000;
array[15682] <= 16'b0000_0000_0000_0000;
array[15683] <= 16'b0000_0000_0000_0000;
array[15684] <= 16'b0000_0000_0000_0000;
array[15685] <= 16'b0000_0000_0000_0000;
array[15686] <= 16'b0000_0000_0000_0000;
array[15687] <= 16'b0000_0000_0000_0000;
array[15688] <= 16'b0000_0000_0000_0000;
array[15689] <= 16'b0000_0000_0000_0000;
array[15690] <= 16'b0000_0000_0000_0000;
array[15691] <= 16'b0000_0000_0000_0000;
array[15692] <= 16'b0000_0000_0000_0000;
array[15693] <= 16'b0000_0000_0000_0000;
array[15694] <= 16'b0000_0000_0000_0000;
array[15695] <= 16'b0000_0000_0000_0000;
array[15696] <= 16'b0000_0000_0000_0000;
array[15697] <= 16'b0000_0000_0000_0000;
array[15698] <= 16'b0000_0000_0000_0000;
array[15699] <= 16'b0000_0000_0000_0000;
array[15700] <= 16'b0000_0000_0000_0000;
array[15701] <= 16'b0000_0000_0000_0000;
array[15702] <= 16'b0000_0000_0000_0000;
array[15703] <= 16'b0000_0000_0000_0000;
array[15704] <= 16'b0000_0000_0000_0000;
array[15705] <= 16'b0000_0000_0000_0000;
array[15706] <= 16'b0000_0000_0000_0000;
array[15707] <= 16'b0000_0000_0000_0000;
array[15708] <= 16'b0000_0000_0000_0000;
array[15709] <= 16'b0000_0000_0000_0000;
array[15710] <= 16'b0000_0000_0000_0000;
array[15711] <= 16'b0000_0000_0000_0000;
array[15712] <= 16'b0000_0000_0000_0000;
array[15713] <= 16'b0000_0000_0000_0000;
array[15714] <= 16'b0000_0000_0000_0000;
array[15715] <= 16'b0000_0000_0000_0000;
array[15716] <= 16'b0000_0000_0000_0000;
array[15717] <= 16'b0000_0000_0000_0000;
array[15718] <= 16'b0000_0000_0000_0000;
array[15719] <= 16'b0000_0000_0000_0000;
array[15720] <= 16'b0000_0000_0000_0000;
array[15721] <= 16'b0000_0000_0000_0000;
array[15722] <= 16'b0000_0000_0000_0000;
array[15723] <= 16'b0000_0000_0000_0000;
array[15724] <= 16'b0000_0000_0000_0000;
array[15725] <= 16'b0000_0000_0000_0000;
array[15726] <= 16'b0000_0000_0000_0000;
array[15727] <= 16'b0000_0000_0000_0000;
array[15728] <= 16'b0000_0000_0000_0000;
array[15729] <= 16'b0000_0000_0000_0000;
array[15730] <= 16'b0000_0000_0000_0000;
array[15731] <= 16'b0000_0000_0000_0000;
array[15732] <= 16'b0000_0000_0000_0000;
array[15733] <= 16'b0000_0000_0000_0000;
array[15734] <= 16'b0000_0000_0000_0000;
array[15735] <= 16'b0000_0000_0000_0000;
array[15736] <= 16'b0000_0000_0000_0000;
array[15737] <= 16'b0000_0000_0000_0000;
array[15738] <= 16'b0000_0000_0000_0000;
array[15739] <= 16'b0000_0000_0000_0000;
array[15740] <= 16'b0000_0000_0000_0000;
array[15741] <= 16'b0000_0000_0000_0000;
array[15742] <= 16'b0000_0000_0000_0000;
array[15743] <= 16'b0000_0000_0000_0000;
array[15744] <= 16'b0000_0000_0000_0000;
array[15745] <= 16'b0000_0000_0000_0000;
array[15746] <= 16'b0000_0000_0000_0000;
array[15747] <= 16'b0000_0000_0000_0000;
array[15748] <= 16'b0000_0000_0000_0000;
array[15749] <= 16'b0000_0000_0000_0000;
array[15750] <= 16'b0000_0000_0000_0000;
array[15751] <= 16'b0000_0000_0000_0000;
array[15752] <= 16'b0000_0000_0000_0000;
array[15753] <= 16'b0000_0000_0000_0000;
array[15754] <= 16'b0000_0000_0000_0000;
array[15755] <= 16'b0000_0000_0000_0000;
array[15756] <= 16'b0000_0000_0000_0000;
array[15757] <= 16'b0000_0000_0000_0000;
array[15758] <= 16'b0000_0000_0000_0000;
array[15759] <= 16'b0000_0000_0000_0000;
array[15760] <= 16'b0000_0000_0000_0000;
array[15761] <= 16'b0000_0000_0000_0000;
array[15762] <= 16'b0000_0000_0000_0000;
array[15763] <= 16'b0000_0000_0000_0000;
array[15764] <= 16'b0000_0000_0000_0000;
array[15765] <= 16'b0000_0000_0000_0000;
array[15766] <= 16'b0000_0000_0000_0000;
array[15767] <= 16'b0000_0000_0000_0000;
array[15768] <= 16'b0000_0000_0000_0000;
array[15769] <= 16'b0000_0000_0000_0000;
array[15770] <= 16'b0000_0000_0000_0000;
array[15771] <= 16'b0000_0000_0000_0000;
array[15772] <= 16'b0000_0000_0000_0000;
array[15773] <= 16'b0000_0000_0000_0000;
array[15774] <= 16'b0000_0000_0000_0000;
array[15775] <= 16'b0000_0000_0000_0000;
array[15776] <= 16'b0000_0000_0000_0000;
array[15777] <= 16'b0000_0000_0000_0000;
array[15778] <= 16'b0000_0000_0000_0000;
array[15779] <= 16'b0000_0000_0000_0000;
array[15780] <= 16'b0000_0000_0000_0000;
array[15781] <= 16'b0000_0000_0000_0000;
array[15782] <= 16'b0000_0000_0000_0000;
array[15783] <= 16'b0000_0000_0000_0000;
array[15784] <= 16'b0000_0000_0000_0000;
array[15785] <= 16'b0000_0000_0000_0000;
array[15786] <= 16'b0000_0000_0000_0000;
array[15787] <= 16'b0000_0000_0000_0000;
array[15788] <= 16'b0000_0000_0000_0000;
array[15789] <= 16'b0000_0000_0000_0000;
array[15790] <= 16'b0000_0000_0000_0000;
array[15791] <= 16'b0000_0000_0000_0000;
array[15792] <= 16'b0000_0000_0000_0000;
array[15793] <= 16'b0000_0000_0000_0000;
array[15794] <= 16'b0000_0000_0000_0000;
array[15795] <= 16'b0000_0000_0000_0000;
array[15796] <= 16'b0000_0000_0000_0000;
array[15797] <= 16'b0000_0000_0000_0000;
array[15798] <= 16'b0000_0000_0000_0000;
array[15799] <= 16'b0000_0000_0000_0000;
array[15800] <= 16'b0000_0000_0000_0000;
array[15801] <= 16'b0000_0000_0000_0000;
array[15802] <= 16'b0000_0000_0000_0000;
array[15803] <= 16'b0000_0000_0000_0000;
array[15804] <= 16'b0000_0000_0000_0000;
array[15805] <= 16'b0000_0000_0000_0000;
array[15806] <= 16'b0000_0000_0000_0000;
array[15807] <= 16'b0000_0000_0000_0000;
array[15808] <= 16'b0000_0000_0000_0000;
array[15809] <= 16'b0000_0000_0000_0000;
array[15810] <= 16'b0000_0000_0000_0000;
array[15811] <= 16'b0000_0000_0000_0000;
array[15812] <= 16'b0000_0000_0000_0000;
array[15813] <= 16'b0000_0000_0000_0000;
array[15814] <= 16'b0000_0000_0000_0000;
array[15815] <= 16'b0000_0000_0000_0000;
array[15816] <= 16'b0000_0000_0000_0000;
array[15817] <= 16'b0000_0000_0000_0000;
array[15818] <= 16'b0000_0000_0000_0000;
array[15819] <= 16'b0000_0000_0000_0000;
array[15820] <= 16'b0000_0000_0000_0000;
array[15821] <= 16'b0000_0000_0000_0000;
array[15822] <= 16'b0000_0000_0000_0000;
array[15823] <= 16'b0000_0000_0000_0000;
array[15824] <= 16'b0000_0000_0000_0000;
array[15825] <= 16'b0000_0000_0000_0000;
array[15826] <= 16'b0000_0000_0000_0000;
array[15827] <= 16'b0000_0000_0000_0000;
array[15828] <= 16'b0000_0000_0000_0000;
array[15829] <= 16'b0000_0000_0000_0000;
array[15830] <= 16'b0000_0000_0000_0000;
array[15831] <= 16'b0000_0000_0000_0000;
array[15832] <= 16'b0000_0000_0000_0000;
array[15833] <= 16'b0000_0000_0000_0000;
array[15834] <= 16'b0000_0000_0000_0000;
array[15835] <= 16'b0000_0000_0000_0000;
array[15836] <= 16'b0000_0000_0000_0000;
array[15837] <= 16'b0000_0000_0000_0000;
array[15838] <= 16'b0000_0000_0000_0000;
array[15839] <= 16'b0000_0000_0000_0000;
array[15840] <= 16'b0000_0000_0000_0000;
array[15841] <= 16'b0000_0000_0000_0000;
array[15842] <= 16'b0000_0000_0000_0000;
array[15843] <= 16'b0000_0000_0000_0000;
array[15844] <= 16'b0000_0000_0000_0000;
array[15845] <= 16'b0000_0000_0000_0000;
array[15846] <= 16'b0000_0000_0000_0000;
array[15847] <= 16'b0000_0000_0000_0000;
array[15848] <= 16'b0000_0000_0000_0000;
array[15849] <= 16'b0000_0000_0000_0000;
array[15850] <= 16'b0000_0000_0000_0000;
array[15851] <= 16'b0000_0000_0000_0000;
array[15852] <= 16'b0000_0000_0000_0000;
array[15853] <= 16'b0000_0000_0000_0000;
array[15854] <= 16'b0000_0000_0000_0000;
array[15855] <= 16'b0000_0000_0000_0000;
array[15856] <= 16'b0000_0000_0000_0000;
array[15857] <= 16'b0000_0000_0000_0000;
array[15858] <= 16'b0000_0000_0000_0000;
array[15859] <= 16'b0000_0000_0000_0000;
array[15860] <= 16'b0000_0000_0000_0000;
array[15861] <= 16'b0000_0000_0000_0000;
array[15862] <= 16'b0000_0000_0000_0000;
array[15863] <= 16'b0000_0000_0000_0000;
array[15864] <= 16'b0000_0000_0000_0000;
array[15865] <= 16'b0000_0000_0000_0000;
array[15866] <= 16'b0000_0000_0000_0000;
array[15867] <= 16'b0000_0000_0000_0000;
array[15868] <= 16'b0000_0000_0000_0000;
array[15869] <= 16'b0000_0000_0000_0000;
array[15870] <= 16'b0000_0000_0000_0000;
array[15871] <= 16'b0000_0000_0000_0000;
array[15872] <= 16'b0000_0000_0000_0000;
array[15873] <= 16'b0000_0000_0000_0000;
array[15874] <= 16'b0000_0000_0000_0000;
array[15875] <= 16'b0000_0000_0000_0000;
array[15876] <= 16'b0000_0000_0000_0000;
array[15877] <= 16'b0000_0000_0000_0000;
array[15878] <= 16'b0000_0000_0000_0000;
array[15879] <= 16'b0000_0000_0000_0000;
array[15880] <= 16'b0000_0000_0000_0000;
array[15881] <= 16'b0000_0000_0000_0000;
array[15882] <= 16'b0000_0000_0000_0000;
array[15883] <= 16'b0000_0000_0000_0000;
array[15884] <= 16'b0000_0000_0000_0000;
array[15885] <= 16'b0000_0000_0000_0000;
array[15886] <= 16'b0000_0000_0000_0000;
array[15887] <= 16'b0000_0000_0000_0000;
array[15888] <= 16'b0000_0000_0000_0000;
array[15889] <= 16'b0000_0000_0000_0000;
array[15890] <= 16'b0000_0000_0000_0000;
array[15891] <= 16'b0000_0000_0000_0000;
array[15892] <= 16'b0000_0000_0000_0000;
array[15893] <= 16'b0000_0000_0000_0000;
array[15894] <= 16'b0000_0000_0000_0000;
array[15895] <= 16'b0000_0000_0000_0000;
array[15896] <= 16'b0000_0000_0000_0000;
array[15897] <= 16'b0000_0000_0000_0000;
array[15898] <= 16'b0000_0000_0000_0000;
array[15899] <= 16'b0000_0000_0000_0000;
array[15900] <= 16'b0000_0000_0000_0000;
array[15901] <= 16'b0000_0000_0000_0000;
array[15902] <= 16'b0000_0000_0000_0000;
array[15903] <= 16'b0000_0000_0000_0000;
array[15904] <= 16'b0000_0000_0000_0000;
array[15905] <= 16'b0000_0000_0000_0000;
array[15906] <= 16'b0000_0000_0000_0000;
array[15907] <= 16'b0000_0000_0000_0000;
array[15908] <= 16'b0000_0000_0000_0000;
array[15909] <= 16'b0000_0000_0000_0000;
array[15910] <= 16'b0000_0000_0000_0000;
array[15911] <= 16'b0000_0000_0000_0000;
array[15912] <= 16'b0000_0000_0000_0000;
array[15913] <= 16'b0000_0000_0000_0000;
array[15914] <= 16'b0000_0000_0000_0000;
array[15915] <= 16'b0000_0000_0000_0000;
array[15916] <= 16'b0000_0000_0000_0000;
array[15917] <= 16'b0000_0000_0000_0000;
array[15918] <= 16'b0000_0000_0000_0000;
array[15919] <= 16'b0000_0000_0000_0000;
array[15920] <= 16'b0000_0000_0000_0000;
array[15921] <= 16'b0000_0000_0000_0000;
array[15922] <= 16'b0000_0000_0000_0000;
array[15923] <= 16'b0000_0000_0000_0000;
array[15924] <= 16'b0000_0000_0000_0000;
array[15925] <= 16'b0000_0000_0000_0000;
array[15926] <= 16'b0000_0000_0000_0000;
array[15927] <= 16'b0000_0000_0000_0000;
array[15928] <= 16'b0000_0000_0000_0000;
array[15929] <= 16'b0000_0000_0000_0000;
array[15930] <= 16'b0000_0000_0000_0000;
array[15931] <= 16'b0000_0000_0000_0000;
array[15932] <= 16'b0000_0000_0000_0000;
array[15933] <= 16'b0000_0000_0000_0000;
array[15934] <= 16'b0000_0000_0000_0000;
array[15935] <= 16'b0000_0000_0000_0000;
array[15936] <= 16'b0000_0000_0000_0000;
array[15937] <= 16'b0000_0000_0000_0000;
array[15938] <= 16'b0000_0000_0000_0000;
array[15939] <= 16'b0000_0000_0000_0000;
array[15940] <= 16'b0000_0000_0000_0000;
array[15941] <= 16'b0000_0000_0000_0000;
array[15942] <= 16'b0000_0000_0000_0000;
array[15943] <= 16'b0000_0000_0000_0000;
array[15944] <= 16'b0000_0000_0000_0000;
array[15945] <= 16'b0000_0000_0000_0000;
array[15946] <= 16'b0000_0000_0000_0000;
array[15947] <= 16'b0000_0000_0000_0000;
array[15948] <= 16'b0000_0000_0000_0000;
array[15949] <= 16'b0000_0000_0000_0000;
array[15950] <= 16'b0000_0000_0000_0000;
array[15951] <= 16'b0000_0000_0000_0000;
array[15952] <= 16'b0000_0000_0000_0000;
array[15953] <= 16'b0000_0000_0000_0000;
array[15954] <= 16'b0000_0000_0000_0000;
array[15955] <= 16'b0000_0000_0000_0000;
array[15956] <= 16'b0000_0000_0000_0000;
array[15957] <= 16'b0000_0000_0000_0000;
array[15958] <= 16'b0000_0000_0000_0000;
array[15959] <= 16'b0000_0000_0000_0000;
array[15960] <= 16'b0000_0000_0000_0000;
array[15961] <= 16'b0000_0000_0000_0000;
array[15962] <= 16'b0000_0000_0000_0000;
array[15963] <= 16'b0000_0000_0000_0000;
array[15964] <= 16'b0000_0000_0000_0000;
array[15965] <= 16'b0000_0000_0000_0000;
array[15966] <= 16'b0000_0000_0000_0000;
array[15967] <= 16'b0000_0000_0000_0000;
array[15968] <= 16'b0000_0000_0000_0000;
array[15969] <= 16'b0000_0000_0000_0000;
array[15970] <= 16'b0000_0000_0000_0000;
array[15971] <= 16'b0000_0000_0000_0000;
array[15972] <= 16'b0000_0000_0000_0000;
array[15973] <= 16'b0000_0000_0000_0000;
array[15974] <= 16'b0000_0000_0000_0000;
array[15975] <= 16'b0000_0000_0000_0000;
array[15976] <= 16'b0000_0000_0000_0000;
array[15977] <= 16'b0000_0000_0000_0000;
array[15978] <= 16'b0000_0000_0000_0000;
array[15979] <= 16'b0000_0000_0000_0000;
array[15980] <= 16'b0000_0000_0000_0000;
array[15981] <= 16'b0000_0000_0000_0000;
array[15982] <= 16'b0000_0000_0000_0000;
array[15983] <= 16'b0000_0000_0000_0000;
array[15984] <= 16'b0000_0000_0000_0000;
array[15985] <= 16'b0000_0000_0000_0000;
array[15986] <= 16'b0000_0000_0000_0000;
array[15987] <= 16'b0000_0000_0000_0000;
array[15988] <= 16'b0000_0000_0000_0000;
array[15989] <= 16'b0000_0000_0000_0000;
array[15990] <= 16'b0000_0000_0000_0000;
array[15991] <= 16'b0000_0000_0000_0000;
array[15992] <= 16'b0000_0000_0000_0000;
array[15993] <= 16'b0000_0000_0000_0000;
array[15994] <= 16'b0000_0000_0000_0000;
array[15995] <= 16'b0000_0000_0000_0000;
array[15996] <= 16'b0000_0000_0000_0000;
array[15997] <= 16'b0000_0000_0000_0000;
array[15998] <= 16'b0000_0000_0000_0000;
array[15999] <= 16'b0000_0000_0000_0000;
array[16000] <= 16'b0000_0000_0000_0000;
array[16001] <= 16'b0000_0000_0000_0000;
array[16002] <= 16'b0000_0000_0000_0000;
array[16003] <= 16'b0000_0000_0000_0000;
array[16004] <= 16'b0000_0000_0000_0000;
array[16005] <= 16'b0000_0000_0000_0000;
array[16006] <= 16'b0000_0000_0000_0000;
array[16007] <= 16'b0000_0000_0000_0000;
array[16008] <= 16'b0000_0000_0000_0000;
array[16009] <= 16'b0000_0000_0000_0000;
array[16010] <= 16'b0000_0000_0000_0000;
array[16011] <= 16'b0000_0000_0000_0000;
array[16012] <= 16'b0000_0000_0000_0000;
array[16013] <= 16'b0000_0000_0000_0000;
array[16014] <= 16'b0000_0000_0000_0000;
array[16015] <= 16'b0000_0000_0000_0000;
array[16016] <= 16'b0000_0000_0000_0000;
array[16017] <= 16'b0000_0000_0000_0000;
array[16018] <= 16'b0000_0000_0000_0000;
array[16019] <= 16'b0000_0000_0000_0000;
array[16020] <= 16'b0000_0000_0000_0000;
array[16021] <= 16'b0000_0000_0000_0000;
array[16022] <= 16'b0000_0000_0000_0000;
array[16023] <= 16'b0000_0000_0000_0000;
array[16024] <= 16'b0000_0000_0000_0000;
array[16025] <= 16'b0000_0000_0000_0000;
array[16026] <= 16'b0000_0000_0000_0000;
array[16027] <= 16'b0000_0000_0000_0000;
array[16028] <= 16'b0000_0000_0000_0000;
array[16029] <= 16'b0000_0000_0000_0000;
array[16030] <= 16'b0000_0000_0000_0000;
array[16031] <= 16'b0000_0000_0000_0000;
array[16032] <= 16'b0000_0000_0000_0000;
array[16033] <= 16'b0000_0000_0000_0000;
array[16034] <= 16'b0000_0000_0000_0000;
array[16035] <= 16'b0000_0000_0000_0000;
array[16036] <= 16'b0000_0000_0000_0000;
array[16037] <= 16'b0000_0000_0000_0000;
array[16038] <= 16'b0000_0000_0000_0000;
array[16039] <= 16'b0000_0000_0000_0000;
array[16040] <= 16'b0000_0000_0000_0000;
array[16041] <= 16'b0000_0000_0000_0000;
array[16042] <= 16'b0000_0000_0000_0000;
array[16043] <= 16'b0000_0000_0000_0000;
array[16044] <= 16'b0000_0000_0000_0000;
array[16045] <= 16'b0000_0000_0000_0000;
array[16046] <= 16'b0000_0000_0000_0000;
array[16047] <= 16'b0000_0000_0000_0000;
array[16048] <= 16'b0000_0000_0000_0000;
array[16049] <= 16'b0000_0000_0000_0000;
array[16050] <= 16'b0000_0000_0000_0000;
array[16051] <= 16'b0000_0000_0000_0000;
array[16052] <= 16'b0000_0000_0000_0000;
array[16053] <= 16'b0000_0000_0000_0000;
array[16054] <= 16'b0000_0000_0000_0000;
array[16055] <= 16'b0000_0000_0000_0000;
array[16056] <= 16'b0000_0000_0000_0000;
array[16057] <= 16'b0000_0000_0000_0000;
array[16058] <= 16'b0000_0000_0000_0000;
array[16059] <= 16'b0000_0000_0000_0000;
array[16060] <= 16'b0000_0000_0000_0000;
array[16061] <= 16'b0000_0000_0000_0000;
array[16062] <= 16'b0000_0000_0000_0000;
array[16063] <= 16'b0000_0000_0000_0000;
array[16064] <= 16'b0000_0000_0000_0000;
array[16065] <= 16'b0000_0000_0000_0000;
array[16066] <= 16'b0000_0000_0000_0000;
array[16067] <= 16'b0000_0000_0000_0000;
array[16068] <= 16'b0000_0000_0000_0000;
array[16069] <= 16'b0000_0000_0000_0000;
array[16070] <= 16'b0000_0000_0000_0000;
array[16071] <= 16'b0000_0000_0000_0000;
array[16072] <= 16'b0000_0000_0000_0000;
array[16073] <= 16'b0000_0000_0000_0000;
array[16074] <= 16'b0000_0000_0000_0000;
array[16075] <= 16'b0000_0000_0000_0000;
array[16076] <= 16'b0000_0000_0000_0000;
array[16077] <= 16'b0000_0000_0000_0000;
array[16078] <= 16'b0000_0000_0000_0000;
array[16079] <= 16'b0000_0000_0000_0000;
array[16080] <= 16'b0000_0000_0000_0000;
array[16081] <= 16'b0000_0000_0000_0000;
array[16082] <= 16'b0000_0000_0000_0000;
array[16083] <= 16'b0000_0000_0000_0000;
array[16084] <= 16'b0000_0000_0000_0000;
array[16085] <= 16'b0000_0000_0000_0000;
array[16086] <= 16'b0000_0000_0000_0000;
array[16087] <= 16'b0000_0000_0000_0000;
array[16088] <= 16'b0000_0000_0000_0000;
array[16089] <= 16'b0000_0000_0000_0000;
array[16090] <= 16'b0000_0000_0000_0000;
array[16091] <= 16'b0000_0000_0000_0000;
array[16092] <= 16'b0000_0000_0000_0000;
array[16093] <= 16'b0000_0000_0000_0000;
array[16094] <= 16'b0000_0000_0000_0000;
array[16095] <= 16'b0000_0000_0000_0000;
array[16096] <= 16'b0000_0000_0000_0000;
array[16097] <= 16'b0000_0000_0000_0000;
array[16098] <= 16'b0000_0000_0000_0000;
array[16099] <= 16'b0000_0000_0000_0000;
array[16100] <= 16'b0000_0000_0000_0000;
array[16101] <= 16'b0000_0000_0000_0000;
array[16102] <= 16'b0000_0000_0000_0000;
array[16103] <= 16'b0000_0000_0000_0000;
array[16104] <= 16'b0000_0000_0000_0000;
array[16105] <= 16'b0000_0000_0000_0000;
array[16106] <= 16'b0000_0000_0000_0000;
array[16107] <= 16'b0000_0000_0000_0000;
array[16108] <= 16'b0000_0000_0000_0000;
array[16109] <= 16'b0000_0000_0000_0000;
array[16110] <= 16'b0000_0000_0000_0000;
array[16111] <= 16'b0000_0000_0000_0000;
array[16112] <= 16'b0000_0000_0000_0000;
array[16113] <= 16'b0000_0000_0000_0000;
array[16114] <= 16'b0000_0000_0000_0000;
array[16115] <= 16'b0000_0000_0000_0000;
array[16116] <= 16'b0000_0000_0000_0000;
array[16117] <= 16'b0000_0000_0000_0000;
array[16118] <= 16'b0000_0000_0000_0000;
array[16119] <= 16'b0000_0000_0000_0000;
array[16120] <= 16'b0000_0000_0000_0000;
array[16121] <= 16'b0000_0000_0000_0000;
array[16122] <= 16'b0000_0000_0000_0000;
array[16123] <= 16'b0000_0000_0000_0000;
array[16124] <= 16'b0000_0000_0000_0000;
array[16125] <= 16'b0000_0000_0000_0000;
array[16126] <= 16'b0000_0000_0000_0000;
array[16127] <= 16'b0000_0000_0000_0000;
array[16128] <= 16'b0000_0000_0000_0000;
array[16129] <= 16'b0000_0000_0000_0000;
array[16130] <= 16'b0000_0000_0000_0000;
array[16131] <= 16'b0000_0000_0000_0000;
array[16132] <= 16'b0000_0000_0000_0000;
array[16133] <= 16'b0000_0000_0000_0000;
array[16134] <= 16'b0000_0000_0000_0000;
array[16135] <= 16'b0000_0000_0000_0000;
array[16136] <= 16'b0000_0000_0000_0000;
array[16137] <= 16'b0000_0000_0000_0000;
array[16138] <= 16'b0000_0000_0000_0000;
array[16139] <= 16'b0000_0000_0000_0000;
array[16140] <= 16'b0000_0000_0000_0000;
array[16141] <= 16'b0000_0000_0000_0000;
array[16142] <= 16'b0000_0000_0000_0000;
array[16143] <= 16'b0000_0000_0000_0000;
array[16144] <= 16'b0000_0000_0000_0000;
array[16145] <= 16'b0000_0000_0000_0000;
array[16146] <= 16'b0000_0000_0000_0000;
array[16147] <= 16'b0000_0000_0000_0000;
array[16148] <= 16'b0000_0000_0000_0000;
array[16149] <= 16'b0000_0000_0000_0000;
array[16150] <= 16'b0000_0000_0000_0000;
array[16151] <= 16'b0000_0000_0000_0000;
array[16152] <= 16'b0000_0000_0000_0000;
array[16153] <= 16'b0000_0000_0000_0000;
array[16154] <= 16'b0000_0000_0000_0000;
array[16155] <= 16'b0000_0000_0000_0000;
array[16156] <= 16'b0000_0000_0000_0000;
array[16157] <= 16'b0000_0000_0000_0000;
array[16158] <= 16'b0000_0000_0000_0000;
array[16159] <= 16'b0000_0000_0000_0000;
array[16160] <= 16'b0000_0000_0000_0000;
array[16161] <= 16'b0000_0000_0000_0000;
array[16162] <= 16'b0000_0000_0000_0000;
array[16163] <= 16'b0000_0000_0000_0000;
array[16164] <= 16'b0000_0000_0000_0000;
array[16165] <= 16'b0000_0000_0000_0000;
array[16166] <= 16'b0000_0000_0000_0000;
array[16167] <= 16'b0000_0000_0000_0000;
array[16168] <= 16'b0000_0000_0000_0000;
array[16169] <= 16'b0000_0000_0000_0000;
array[16170] <= 16'b0000_0000_0000_0000;
array[16171] <= 16'b0000_0000_0000_0000;
array[16172] <= 16'b0000_0000_0000_0000;
array[16173] <= 16'b0000_0000_0000_0000;
array[16174] <= 16'b0000_0000_0000_0000;
array[16175] <= 16'b0000_0000_0000_0000;
array[16176] <= 16'b0000_0000_0000_0000;
array[16177] <= 16'b0000_0000_0000_0000;
array[16178] <= 16'b0000_0000_0000_0000;
array[16179] <= 16'b0000_0000_0000_0000;
array[16180] <= 16'b0000_0000_0000_0000;
array[16181] <= 16'b0000_0000_0000_0000;
array[16182] <= 16'b0000_0000_0000_0000;
array[16183] <= 16'b0000_0000_0000_0000;
array[16184] <= 16'b0000_0000_0000_0000;
array[16185] <= 16'b0000_0000_0000_0000;
array[16186] <= 16'b0000_0000_0000_0000;
array[16187] <= 16'b0000_0000_0000_0000;
array[16188] <= 16'b0000_0000_0000_0000;
array[16189] <= 16'b0000_0000_0000_0000;
array[16190] <= 16'b0000_0000_0000_0000;
array[16191] <= 16'b0000_0000_0000_0000;
array[16192] <= 16'b0000_0000_0000_0000;
array[16193] <= 16'b0000_0000_0000_0000;
array[16194] <= 16'b0000_0000_0000_0000;
array[16195] <= 16'b0000_0000_0000_0000;
array[16196] <= 16'b0000_0000_0000_0000;
array[16197] <= 16'b0000_0000_0000_0000;
array[16198] <= 16'b0000_0000_0000_0000;
array[16199] <= 16'b0000_0000_0000_0000;
array[16200] <= 16'b0000_0000_0000_0000;
array[16201] <= 16'b0000_0000_0000_0000;
array[16202] <= 16'b0000_0000_0000_0000;
array[16203] <= 16'b0000_0000_0000_0000;
array[16204] <= 16'b0000_0000_0000_0000;
array[16205] <= 16'b0000_0000_0000_0000;
array[16206] <= 16'b0000_0000_0000_0000;
array[16207] <= 16'b0000_0000_0000_0000;
array[16208] <= 16'b0000_0000_0000_0000;
array[16209] <= 16'b0000_0000_0000_0000;
array[16210] <= 16'b0000_0000_0000_0000;
array[16211] <= 16'b0000_0000_0000_0000;
array[16212] <= 16'b0000_0000_0000_0000;
array[16213] <= 16'b0000_0000_0000_0000;
array[16214] <= 16'b0000_0000_0000_0000;
array[16215] <= 16'b0000_0000_0000_0000;
array[16216] <= 16'b0000_0000_0000_0000;
array[16217] <= 16'b0000_0000_0000_0000;
array[16218] <= 16'b0000_0000_0000_0000;
array[16219] <= 16'b0000_0000_0000_0000;
array[16220] <= 16'b0000_0000_0000_0000;
array[16221] <= 16'b0000_0000_0000_0000;
array[16222] <= 16'b0000_0000_0000_0000;
array[16223] <= 16'b0000_0000_0000_0000;
array[16224] <= 16'b0000_0000_0000_0000;
array[16225] <= 16'b0000_0000_0000_0000;
array[16226] <= 16'b0000_0000_0000_0000;
array[16227] <= 16'b0000_0000_0000_0000;
array[16228] <= 16'b0000_0000_0000_0000;
array[16229] <= 16'b0000_0000_0000_0000;
array[16230] <= 16'b0000_0000_0000_0000;
array[16231] <= 16'b0000_0000_0000_0000;
array[16232] <= 16'b0000_0000_0000_0000;
array[16233] <= 16'b0000_0000_0000_0000;
array[16234] <= 16'b0000_0000_0000_0000;
array[16235] <= 16'b0000_0000_0000_0000;
array[16236] <= 16'b0000_0000_0000_0000;
array[16237] <= 16'b0000_0000_0000_0000;
array[16238] <= 16'b0000_0000_0000_0000;
array[16239] <= 16'b0000_0000_0000_0000;
array[16240] <= 16'b0000_0000_0000_0000;
array[16241] <= 16'b0000_0000_0000_0000;
array[16242] <= 16'b0000_0000_0000_0000;
array[16243] <= 16'b0000_0000_0000_0000;
array[16244] <= 16'b0000_0000_0000_0000;
array[16245] <= 16'b0000_0000_0000_0000;
array[16246] <= 16'b0000_0000_0000_0000;
array[16247] <= 16'b0000_0000_0000_0000;
array[16248] <= 16'b0000_0000_0000_0000;
array[16249] <= 16'b0000_0000_0000_0000;
array[16250] <= 16'b0000_0000_0000_0000;
array[16251] <= 16'b0000_0000_0000_0000;
array[16252] <= 16'b0000_0000_0000_0000;
array[16253] <= 16'b0000_0000_0000_0000;
array[16254] <= 16'b0000_0000_0000_0000;
array[16255] <= 16'b0000_0000_0000_0000;
array[16256] <= 16'b0000_0000_0000_0000;
array[16257] <= 16'b0000_0000_0000_0000;
array[16258] <= 16'b0000_0000_0000_0000;
array[16259] <= 16'b0000_0000_0000_0000;
array[16260] <= 16'b0000_0000_0000_0000;
array[16261] <= 16'b0000_0000_0000_0000;
array[16262] <= 16'b0000_0000_0000_0000;
array[16263] <= 16'b0000_0000_0000_0000;
array[16264] <= 16'b0000_0000_0000_0000;
array[16265] <= 16'b0000_0000_0000_0000;
array[16266] <= 16'b0000_0000_0000_0000;
array[16267] <= 16'b0000_0000_0000_0000;
array[16268] <= 16'b0000_0000_0000_0000;
array[16269] <= 16'b0000_0000_0000_0000;
array[16270] <= 16'b0000_0000_0000_0000;
array[16271] <= 16'b0000_0000_0000_0000;
array[16272] <= 16'b0000_0000_0000_0000;
array[16273] <= 16'b0000_0000_0000_0000;
array[16274] <= 16'b0000_0000_0000_0000;
array[16275] <= 16'b0000_0000_0000_0000;
array[16276] <= 16'b0000_0000_0000_0000;
array[16277] <= 16'b0000_0000_0000_0000;
array[16278] <= 16'b0000_0000_0000_0000;
array[16279] <= 16'b0000_0000_0000_0000;
array[16280] <= 16'b0000_0000_0000_0000;
array[16281] <= 16'b0000_0000_0000_0000;
array[16282] <= 16'b0000_0000_0000_0000;
array[16283] <= 16'b0000_0000_0000_0000;
array[16284] <= 16'b0000_0000_0000_0000;
array[16285] <= 16'b0000_0000_0000_0000;
array[16286] <= 16'b0000_0000_0000_0000;
array[16287] <= 16'b0000_0000_0000_0000;
array[16288] <= 16'b0000_0000_0000_0000;
array[16289] <= 16'b0000_0000_0000_0000;
array[16290] <= 16'b0000_0000_0000_0000;
array[16291] <= 16'b0000_0000_0000_0000;
array[16292] <= 16'b0000_0000_0000_0000;
array[16293] <= 16'b0000_0000_0000_0000;
array[16294] <= 16'b0000_0000_0000_0000;
array[16295] <= 16'b0000_0000_0000_0000;
array[16296] <= 16'b0000_0000_0000_0000;
array[16297] <= 16'b0000_0000_0000_0000;
array[16298] <= 16'b0000_0000_0000_0000;
array[16299] <= 16'b0000_0000_0000_0000;
array[16300] <= 16'b0000_0000_0000_0000;
array[16301] <= 16'b0000_0000_0000_0000;
array[16302] <= 16'b0000_0000_0000_0000;
array[16303] <= 16'b0000_0000_0000_0000;
array[16304] <= 16'b0000_0000_0000_0000;
array[16305] <= 16'b0000_0000_0000_0000;
array[16306] <= 16'b0000_0000_0000_0000;
array[16307] <= 16'b0000_0000_0000_0000;
array[16308] <= 16'b0000_0000_0000_0000;
array[16309] <= 16'b0000_0000_0000_0000;
array[16310] <= 16'b0000_0000_0000_0000;
array[16311] <= 16'b0000_0000_0000_0000;
array[16312] <= 16'b0000_0000_0000_0000;
array[16313] <= 16'b0000_0000_0000_0000;
array[16314] <= 16'b0000_0000_0000_0000;
array[16315] <= 16'b0000_0000_0000_0000;
array[16316] <= 16'b0000_0000_0000_0000;
array[16317] <= 16'b0000_0000_0000_0000;
array[16318] <= 16'b0000_0000_0000_0000;
array[16319] <= 16'b0000_0000_0000_0000;
array[16320] <= 16'b0000_0000_0000_0000;
array[16321] <= 16'b0000_0000_0000_0000;
array[16322] <= 16'b0000_0000_0000_0000;
array[16323] <= 16'b0000_0000_0000_0000;
array[16324] <= 16'b0000_0000_0000_0000;
array[16325] <= 16'b0000_0000_0000_0000;
array[16326] <= 16'b0000_0000_0000_0000;
array[16327] <= 16'b0000_0000_0000_0000;
array[16328] <= 16'b0000_0000_0000_0000;
array[16329] <= 16'b0000_0000_0000_0000;
array[16330] <= 16'b0000_0000_0000_0000;
array[16331] <= 16'b0000_0000_0000_0000;
array[16332] <= 16'b0000_0000_0000_0000;
array[16333] <= 16'b0000_0000_0000_0000;
array[16334] <= 16'b0000_0000_0000_0000;
array[16335] <= 16'b0000_0000_0000_0000;
array[16336] <= 16'b0000_0000_0000_0000;
array[16337] <= 16'b0000_0000_0000_0000;
array[16338] <= 16'b0000_0000_0000_0000;
array[16339] <= 16'b0000_0000_0000_0000;
array[16340] <= 16'b0000_0000_0000_0000;
array[16341] <= 16'b0000_0000_0000_0000;
array[16342] <= 16'b0000_0000_0000_0000;
array[16343] <= 16'b0000_0000_0000_0000;
array[16344] <= 16'b0000_0000_0000_0000;
array[16345] <= 16'b0000_0000_0000_0000;
array[16346] <= 16'b0000_0000_0000_0000;
array[16347] <= 16'b0000_0000_0000_0000;
array[16348] <= 16'b0000_0000_0000_0000;
array[16349] <= 16'b0000_0000_0000_0000;
array[16350] <= 16'b0000_0000_0000_0000;
array[16351] <= 16'b0000_0000_0000_0000;
array[16352] <= 16'b0000_0000_0000_0000;
array[16353] <= 16'b0000_0000_0000_0000;
array[16354] <= 16'b0000_0000_0000_0000;
array[16355] <= 16'b0000_0000_0000_0000;
array[16356] <= 16'b0000_0000_0000_0000;
array[16357] <= 16'b0000_0000_0000_0000;
array[16358] <= 16'b0000_0000_0000_0000;
array[16359] <= 16'b0000_0000_0000_0000;
array[16360] <= 16'b0000_0000_0000_0000;
array[16361] <= 16'b0000_0000_0000_0000;
array[16362] <= 16'b0000_0000_0000_0000;
array[16363] <= 16'b0000_0000_0000_0000;
array[16364] <= 16'b0000_0000_0000_0000;
array[16365] <= 16'b0000_0000_0000_0000;
array[16366] <= 16'b0000_0000_0000_0000;
array[16367] <= 16'b0000_0000_0000_0000;
array[16368] <= 16'b0000_0000_0000_0000;
array[16369] <= 16'b0000_0000_0000_0000;
array[16370] <= 16'b0000_0000_0000_0000;
array[16371] <= 16'b0000_0000_0000_0000;
array[16372] <= 16'b0000_0000_0000_0000;
array[16373] <= 16'b0000_0000_0000_0000;
array[16374] <= 16'b0000_0000_0000_0000;
array[16375] <= 16'b0000_0000_0000_0000;
array[16376] <= 16'b0000_0000_0000_0000;
array[16377] <= 16'b0000_0000_0000_0000;
array[16378] <= 16'b0000_0000_0000_0000;
array[16379] <= 16'b0000_0000_0000_0000;
array[16380] <= 16'b0000_0000_0000_0000;
array[16381] <= 16'b0000_0000_0000_0000;
array[16382] <= 16'b0000_0000_0000_0000;
array[16383] <= 16'b0000_0000_0000_0000;
array[16384] <= 16'b0000_0000_0000_0000;
array[16385] <= 16'b0000_0000_0000_0000;
array[16386] <= 16'b0000_0000_0000_0000;
array[16387] <= 16'b0000_0000_0000_0000;
array[16388] <= 16'b0000_0000_0000_0000;
array[16389] <= 16'b0000_0000_0000_0000;
array[16390] <= 16'b0000_0000_0000_0000;
array[16391] <= 16'b0000_0000_0000_0000;
array[16392] <= 16'b0000_0000_0000_0000;
array[16393] <= 16'b0000_0000_0000_0000;
array[16394] <= 16'b0000_0000_0000_0000;
array[16395] <= 16'b0000_0000_0000_0000;
array[16396] <= 16'b0000_0000_0000_0000;
array[16397] <= 16'b0000_0000_0000_0000;
array[16398] <= 16'b0000_0000_0000_0000;
array[16399] <= 16'b0000_0000_0000_0000;
array[16400] <= 16'b0000_0000_0000_0000;
array[16401] <= 16'b0000_0000_0000_0000;
array[16402] <= 16'b0000_0000_0000_0000;
array[16403] <= 16'b0000_0000_0000_0000;
array[16404] <= 16'b0000_0000_0000_0000;
array[16405] <= 16'b0000_0000_0000_0000;
array[16406] <= 16'b0000_0000_0000_0000;
array[16407] <= 16'b0000_0000_0000_0000;
array[16408] <= 16'b0000_0000_0000_0000;
array[16409] <= 16'b0000_0000_0000_0000;
array[16410] <= 16'b0000_0000_0000_0000;
array[16411] <= 16'b0000_0000_0000_0000;
array[16412] <= 16'b0000_0000_0000_0000;
array[16413] <= 16'b0000_0000_0000_0000;
array[16414] <= 16'b0000_0000_0000_0000;
array[16415] <= 16'b0000_0000_0000_0000;
array[16416] <= 16'b0000_0000_0000_0000;
array[16417] <= 16'b0000_0000_0000_0000;
array[16418] <= 16'b0000_0000_0000_0000;
array[16419] <= 16'b0000_0000_0000_0000;
array[16420] <= 16'b0000_0000_0000_0000;
array[16421] <= 16'b0000_0000_0000_0000;
array[16422] <= 16'b0000_0000_0000_0000;
array[16423] <= 16'b0000_0000_0000_0000;
array[16424] <= 16'b0000_0000_0000_0000;
array[16425] <= 16'b0000_0000_0000_0000;
array[16426] <= 16'b0000_0000_0000_0000;
array[16427] <= 16'b0000_0000_0000_0000;
array[16428] <= 16'b0000_0000_0000_0000;
array[16429] <= 16'b0000_0000_0000_0000;
array[16430] <= 16'b0000_0000_0000_0000;
array[16431] <= 16'b0000_0000_0000_0000;
array[16432] <= 16'b0000_0000_0000_0000;
array[16433] <= 16'b0000_0000_0000_0000;
array[16434] <= 16'b0000_0000_0000_0000;
array[16435] <= 16'b0000_0000_0000_0000;
array[16436] <= 16'b0000_0000_0000_0000;
array[16437] <= 16'b0000_0000_0000_0000;
array[16438] <= 16'b0000_0000_0000_0000;
array[16439] <= 16'b0000_0000_0000_0000;
array[16440] <= 16'b0000_0000_0000_0000;
array[16441] <= 16'b0000_0000_0000_0000;
array[16442] <= 16'b0000_0000_0000_0000;
array[16443] <= 16'b0000_0000_0000_0000;
array[16444] <= 16'b0000_0000_0000_0000;
array[16445] <= 16'b0000_0000_0000_0000;
array[16446] <= 16'b0000_0000_0000_0000;
array[16447] <= 16'b0000_0000_0000_0000;
array[16448] <= 16'b0000_0000_0000_0000;
array[16449] <= 16'b0000_0000_0000_0000;
array[16450] <= 16'b0000_0000_0000_0000;
array[16451] <= 16'b0000_0000_0000_0000;
array[16452] <= 16'b0000_0000_0000_0000;
array[16453] <= 16'b0000_0000_0000_0000;
array[16454] <= 16'b0000_0000_0000_0000;
array[16455] <= 16'b0000_0000_0000_0000;
array[16456] <= 16'b0000_0000_0000_0000;
array[16457] <= 16'b0000_0000_0000_0000;
array[16458] <= 16'b0000_0000_0000_0000;
array[16459] <= 16'b0000_0000_0000_0000;
array[16460] <= 16'b0000_0000_0000_0000;
array[16461] <= 16'b0000_0000_0000_0000;
array[16462] <= 16'b0000_0000_0000_0000;
array[16463] <= 16'b0000_0000_0000_0000;
array[16464] <= 16'b0000_0000_0000_0000;
array[16465] <= 16'b0000_0000_0000_0000;
array[16466] <= 16'b0000_0000_0000_0000;
array[16467] <= 16'b0000_0000_0000_0000;
array[16468] <= 16'b0000_0000_0000_0000;
array[16469] <= 16'b0000_0000_0000_0000;
array[16470] <= 16'b0000_0000_0000_0000;
array[16471] <= 16'b0000_0000_0000_0000;
array[16472] <= 16'b0000_0000_0000_0000;
array[16473] <= 16'b0000_0000_0000_0000;
array[16474] <= 16'b0000_0000_0000_0000;
array[16475] <= 16'b0000_0000_0000_0000;
array[16476] <= 16'b0000_0000_0000_0000;
array[16477] <= 16'b0000_0000_0000_0000;
array[16478] <= 16'b0000_0000_0000_0000;
array[16479] <= 16'b0000_0000_0000_0000;
array[16480] <= 16'b0000_0000_0000_0000;
array[16481] <= 16'b0000_0000_0000_0000;
array[16482] <= 16'b0000_0000_0000_0000;
array[16483] <= 16'b0000_0000_0000_0000;
array[16484] <= 16'b0000_0000_0000_0000;
array[16485] <= 16'b0000_0000_0000_0000;
array[16486] <= 16'b0000_0000_0000_0000;
array[16487] <= 16'b0000_0000_0000_0000;
array[16488] <= 16'b0000_0000_0000_0000;
array[16489] <= 16'b0000_0000_0000_0000;
array[16490] <= 16'b0000_0000_0000_0000;
array[16491] <= 16'b0000_0000_0000_0000;
array[16492] <= 16'b0000_0000_0000_0000;
array[16493] <= 16'b0000_0000_0000_0000;
array[16494] <= 16'b0000_0000_0000_0000;
array[16495] <= 16'b0000_0000_0000_0000;
array[16496] <= 16'b0000_0000_0000_0000;
array[16497] <= 16'b0000_0000_0000_0000;
array[16498] <= 16'b0000_0000_0000_0000;
array[16499] <= 16'b0000_0000_0000_0000;
array[16500] <= 16'b0000_0000_0000_0000;
array[16501] <= 16'b0000_0000_0000_0000;
array[16502] <= 16'b0000_0000_0000_0000;
array[16503] <= 16'b0000_0000_0000_0000;
array[16504] <= 16'b0000_0000_0000_0000;
array[16505] <= 16'b0000_0000_0000_0000;
array[16506] <= 16'b0000_0000_0000_0000;
array[16507] <= 16'b0000_0000_0000_0000;
array[16508] <= 16'b0000_0000_0000_0000;
array[16509] <= 16'b0000_0000_0000_0000;
array[16510] <= 16'b0000_0000_0000_0000;
array[16511] <= 16'b0000_0000_0000_0000;
array[16512] <= 16'b0000_0000_0000_0000;
array[16513] <= 16'b0000_0000_0000_0000;
array[16514] <= 16'b0000_0000_0000_0000;
array[16515] <= 16'b0000_0000_0000_0000;
array[16516] <= 16'b0000_0000_0000_0000;
array[16517] <= 16'b0000_0000_0000_0000;
array[16518] <= 16'b0000_0000_0000_0000;
array[16519] <= 16'b0000_0000_0000_0000;
array[16520] <= 16'b0000_0000_0000_0000;
array[16521] <= 16'b0000_0000_0000_0000;
array[16522] <= 16'b0000_0000_0000_0000;
array[16523] <= 16'b0000_0000_0000_0000;
array[16524] <= 16'b0000_0000_0000_0000;
array[16525] <= 16'b0000_0000_0000_0000;
array[16526] <= 16'b0000_0000_0000_0000;
array[16527] <= 16'b0000_0000_0000_0000;
array[16528] <= 16'b0000_0000_0000_0000;
array[16529] <= 16'b0000_0000_0000_0000;
array[16530] <= 16'b0000_0000_0000_0000;
array[16531] <= 16'b0000_0000_0000_0000;
array[16532] <= 16'b0000_0000_0000_0000;
array[16533] <= 16'b0000_0000_0000_0000;
array[16534] <= 16'b0000_0000_0000_0000;
array[16535] <= 16'b0000_0000_0000_0000;
array[16536] <= 16'b0000_0000_0000_0000;
array[16537] <= 16'b0000_0000_0000_0000;
array[16538] <= 16'b0000_0000_0000_0000;
array[16539] <= 16'b0000_0000_0000_0000;
array[16540] <= 16'b0000_0000_0000_0000;
array[16541] <= 16'b0000_0000_0000_0000;
array[16542] <= 16'b0000_0000_0000_0000;
array[16543] <= 16'b0000_0000_0000_0000;
array[16544] <= 16'b0000_0000_0000_0000;
array[16545] <= 16'b0000_0000_0000_0000;
array[16546] <= 16'b0000_0000_0000_0000;
array[16547] <= 16'b0000_0000_0000_0000;
array[16548] <= 16'b0000_0000_0000_0000;
array[16549] <= 16'b0000_0000_0000_0000;
array[16550] <= 16'b0000_0000_0000_0000;
array[16551] <= 16'b0000_0000_0000_0000;
array[16552] <= 16'b0000_0000_0000_0000;
array[16553] <= 16'b0000_0000_0000_0000;
array[16554] <= 16'b0000_0000_0000_0000;
array[16555] <= 16'b0000_0000_0000_0000;
array[16556] <= 16'b0000_0000_0000_0000;
array[16557] <= 16'b0000_0000_0000_0000;
array[16558] <= 16'b0000_0000_0000_0000;
array[16559] <= 16'b0000_0000_0000_0000;
array[16560] <= 16'b0000_0000_0000_0000;
array[16561] <= 16'b0000_0000_0000_0000;
array[16562] <= 16'b0000_0000_0000_0000;
array[16563] <= 16'b0000_0000_0000_0000;
array[16564] <= 16'b0000_0000_0000_0000;
array[16565] <= 16'b0000_0000_0000_0000;
array[16566] <= 16'b0000_0000_0000_0000;
array[16567] <= 16'b0000_0000_0000_0000;
array[16568] <= 16'b0000_0000_0000_0000;
array[16569] <= 16'b0000_0000_0000_0000;
array[16570] <= 16'b0000_0000_0000_0000;
array[16571] <= 16'b0000_0000_0000_0000;
array[16572] <= 16'b0000_0000_0000_0000;
array[16573] <= 16'b0000_0000_0000_0000;
array[16574] <= 16'b0000_0000_0000_0000;
array[16575] <= 16'b0000_0000_0000_0000;
array[16576] <= 16'b0000_0000_0000_0000;
array[16577] <= 16'b0000_0000_0000_0000;
array[16578] <= 16'b0000_0000_0000_0000;
array[16579] <= 16'b0000_0000_0000_0000;
array[16580] <= 16'b0000_0000_0000_0000;
array[16581] <= 16'b0000_0000_0000_0000;
array[16582] <= 16'b0000_0000_0000_0000;
array[16583] <= 16'b0000_0000_0000_0000;
array[16584] <= 16'b0000_0000_0000_0000;
array[16585] <= 16'b0000_0000_0000_0000;
array[16586] <= 16'b0000_0000_0000_0000;
array[16587] <= 16'b0000_0000_0000_0000;
array[16588] <= 16'b0000_0000_0000_0000;
array[16589] <= 16'b0000_0000_0000_0000;
array[16590] <= 16'b0000_0000_0000_0000;
array[16591] <= 16'b0000_0000_0000_0000;
array[16592] <= 16'b0000_0000_0000_0000;
array[16593] <= 16'b0000_0000_0000_0000;
array[16594] <= 16'b0000_0000_0000_0000;
array[16595] <= 16'b0000_0000_0000_0000;
array[16596] <= 16'b0000_0000_0000_0000;
array[16597] <= 16'b0000_0000_0000_0000;
array[16598] <= 16'b0000_0000_0000_0000;
array[16599] <= 16'b0000_0000_0000_0000;
array[16600] <= 16'b0000_0000_0000_0000;
array[16601] <= 16'b0000_0000_0000_0000;
array[16602] <= 16'b0000_0000_0000_0000;
array[16603] <= 16'b0000_0000_0000_0000;
array[16604] <= 16'b0000_0000_0000_0000;
array[16605] <= 16'b0000_0000_0000_0000;
array[16606] <= 16'b0000_0000_0000_0000;
array[16607] <= 16'b0000_0000_0000_0000;
array[16608] <= 16'b0000_0000_0000_0000;
array[16609] <= 16'b0000_0000_0000_0000;
array[16610] <= 16'b0000_0000_0000_0000;
array[16611] <= 16'b0000_0000_0000_0000;
array[16612] <= 16'b0000_0000_0000_0000;
array[16613] <= 16'b0000_0000_0000_0000;
array[16614] <= 16'b0000_0000_0000_0000;
array[16615] <= 16'b0000_0000_0000_0000;
array[16616] <= 16'b0000_0000_0000_0000;
array[16617] <= 16'b0000_0000_0000_0000;
array[16618] <= 16'b0000_0000_0000_0000;
array[16619] <= 16'b0000_0000_0000_0000;
array[16620] <= 16'b0000_0000_0000_0000;
array[16621] <= 16'b0000_0000_0000_0000;
array[16622] <= 16'b0000_0000_0000_0000;
array[16623] <= 16'b0000_0000_0000_0000;
array[16624] <= 16'b0000_0000_0000_0000;
array[16625] <= 16'b0000_0000_0000_0000;
array[16626] <= 16'b0000_0000_0000_0000;
array[16627] <= 16'b0000_0000_0000_0000;
array[16628] <= 16'b0000_0000_0000_0000;
array[16629] <= 16'b0000_0000_0000_0000;
array[16630] <= 16'b0000_0000_0000_0000;
array[16631] <= 16'b0000_0000_0000_0000;
array[16632] <= 16'b0000_0000_0000_0000;
array[16633] <= 16'b0000_0000_0000_0000;
array[16634] <= 16'b0000_0000_0000_0000;
array[16635] <= 16'b0000_0000_0000_0000;
array[16636] <= 16'b0000_0000_0000_0000;
array[16637] <= 16'b0000_0000_0000_0000;
array[16638] <= 16'b0000_0000_0000_0000;
array[16639] <= 16'b0000_0000_0000_0000;
array[16640] <= 16'b0000_0000_0000_0000;
array[16641] <= 16'b0000_0000_0000_0000;
array[16642] <= 16'b0000_0000_0000_0000;
array[16643] <= 16'b0000_0000_0000_0000;
array[16644] <= 16'b0000_0000_0000_0000;
array[16645] <= 16'b0000_0000_0000_0000;
array[16646] <= 16'b0000_0000_0000_0000;
array[16647] <= 16'b0000_0000_0000_0000;
array[16648] <= 16'b0000_0000_0000_0000;
array[16649] <= 16'b0000_0000_0000_0000;
array[16650] <= 16'b0000_0000_0000_0000;
array[16651] <= 16'b0000_0000_0000_0000;
array[16652] <= 16'b0000_0000_0000_0000;
array[16653] <= 16'b0000_0000_0000_0000;
array[16654] <= 16'b0000_0000_0000_0000;
array[16655] <= 16'b0000_0000_0000_0000;
array[16656] <= 16'b0000_0000_0000_0000;
array[16657] <= 16'b0000_0000_0000_0000;
array[16658] <= 16'b0000_0000_0000_0000;
array[16659] <= 16'b0000_0000_0000_0000;
array[16660] <= 16'b0000_0000_0000_0000;
array[16661] <= 16'b0000_0000_0000_0000;
array[16662] <= 16'b0000_0000_0000_0000;
array[16663] <= 16'b0000_0000_0000_0000;
array[16664] <= 16'b0000_0000_0000_0000;
array[16665] <= 16'b0000_0000_0000_0000;
array[16666] <= 16'b0000_0000_0000_0000;
array[16667] <= 16'b0000_0000_0000_0000;
array[16668] <= 16'b0000_0000_0000_0000;
array[16669] <= 16'b0000_0000_0000_0000;
array[16670] <= 16'b0000_0000_0000_0000;
array[16671] <= 16'b0000_0000_0000_0000;
array[16672] <= 16'b0000_0000_0000_0000;
array[16673] <= 16'b0000_0000_0000_0000;
array[16674] <= 16'b0000_0000_0000_0000;
array[16675] <= 16'b0000_0000_0000_0000;
array[16676] <= 16'b0000_0000_0000_0000;
array[16677] <= 16'b0000_0000_0000_0000;
array[16678] <= 16'b0000_0000_0000_0000;
array[16679] <= 16'b0000_0000_0000_0000;
array[16680] <= 16'b0000_0000_0000_0000;
array[16681] <= 16'b0000_0000_0000_0000;
array[16682] <= 16'b0000_0000_0000_0000;
array[16683] <= 16'b0000_0000_0000_0000;
array[16684] <= 16'b0000_0000_0000_0000;
array[16685] <= 16'b0000_0000_0000_0000;
array[16686] <= 16'b0000_0000_0000_0000;
array[16687] <= 16'b0000_0000_0000_0000;
array[16688] <= 16'b0000_0000_0000_0000;
array[16689] <= 16'b0000_0000_0000_0000;
array[16690] <= 16'b0000_0000_0000_0000;
array[16691] <= 16'b0000_0000_0000_0000;
array[16692] <= 16'b0000_0000_0000_0000;
array[16693] <= 16'b0000_0000_0000_0000;
array[16694] <= 16'b0000_0000_0000_0000;
array[16695] <= 16'b0000_0000_0000_0000;
array[16696] <= 16'b0000_0000_0000_0000;
array[16697] <= 16'b0000_0000_0000_0000;
array[16698] <= 16'b0000_0000_0000_0000;
array[16699] <= 16'b0000_0000_0000_0000;
array[16700] <= 16'b0000_0000_0000_0000;
array[16701] <= 16'b0000_0000_0000_0000;
array[16702] <= 16'b0000_0000_0000_0000;
array[16703] <= 16'b0000_0000_0000_0000;
array[16704] <= 16'b0000_0000_0000_0000;
array[16705] <= 16'b0000_0000_0000_0000;
array[16706] <= 16'b0000_0000_0000_0000;
array[16707] <= 16'b0000_0000_0000_0000;
array[16708] <= 16'b0000_0000_0000_0000;
array[16709] <= 16'b0000_0000_0000_0000;
array[16710] <= 16'b0000_0000_0000_0000;
array[16711] <= 16'b0000_0000_0000_0000;
array[16712] <= 16'b0000_0000_0000_0000;
array[16713] <= 16'b0000_0000_0000_0000;
array[16714] <= 16'b0000_0000_0000_0000;
array[16715] <= 16'b0000_0000_0000_0000;
array[16716] <= 16'b0000_0000_0000_0000;
array[16717] <= 16'b0000_0000_0000_0000;
array[16718] <= 16'b0000_0000_0000_0000;
array[16719] <= 16'b0000_0000_0000_0000;
array[16720] <= 16'b0000_0000_0000_0000;
array[16721] <= 16'b0000_0000_0000_0000;
array[16722] <= 16'b0000_0000_0000_0000;
array[16723] <= 16'b0000_0000_0000_0000;
array[16724] <= 16'b0000_0000_0000_0000;
array[16725] <= 16'b0000_0000_0000_0000;
array[16726] <= 16'b0000_0000_0000_0000;
array[16727] <= 16'b0000_0000_0000_0000;
array[16728] <= 16'b0000_0000_0000_0000;
array[16729] <= 16'b0000_0000_0000_0000;
array[16730] <= 16'b0000_0000_0000_0000;
array[16731] <= 16'b0000_0000_0000_0000;
array[16732] <= 16'b0000_0000_0000_0000;
array[16733] <= 16'b0000_0000_0000_0000;
array[16734] <= 16'b0000_0000_0000_0000;
array[16735] <= 16'b0000_0000_0000_0000;
array[16736] <= 16'b0000_0000_0000_0000;
array[16737] <= 16'b0000_0000_0000_0000;
array[16738] <= 16'b0000_0000_0000_0000;
array[16739] <= 16'b0000_0000_0000_0000;
array[16740] <= 16'b0000_0000_0000_0000;
array[16741] <= 16'b0000_0000_0000_0000;
array[16742] <= 16'b0000_0000_0000_0000;
array[16743] <= 16'b0000_0000_0000_0000;
array[16744] <= 16'b0000_0000_0000_0000;
array[16745] <= 16'b0000_0000_0000_0000;
array[16746] <= 16'b0000_0000_0000_0000;
array[16747] <= 16'b0000_0000_0000_0000;
array[16748] <= 16'b0000_0000_0000_0000;
array[16749] <= 16'b0000_0000_0000_0000;
array[16750] <= 16'b0000_0000_0000_0000;
array[16751] <= 16'b0000_0000_0000_0000;
array[16752] <= 16'b0000_0000_0000_0000;
array[16753] <= 16'b0000_0000_0000_0000;
array[16754] <= 16'b0000_0000_0000_0000;
array[16755] <= 16'b0000_0000_0000_0000;
array[16756] <= 16'b0000_0000_0000_0000;
array[16757] <= 16'b0000_0000_0000_0000;
array[16758] <= 16'b0000_0000_0000_0000;
array[16759] <= 16'b0000_0000_0000_0000;
array[16760] <= 16'b0000_0000_0000_0000;
array[16761] <= 16'b0000_0000_0000_0000;
array[16762] <= 16'b0000_0000_0000_0000;
array[16763] <= 16'b0000_0000_0000_0000;
array[16764] <= 16'b0000_0000_0000_0000;
array[16765] <= 16'b0000_0000_0000_0000;
array[16766] <= 16'b0000_0000_0000_0000;
array[16767] <= 16'b0000_0000_0000_0000;
array[16768] <= 16'b0000_0000_0000_0000;
array[16769] <= 16'b0000_0000_0000_0000;
array[16770] <= 16'b0000_0000_0000_0000;
array[16771] <= 16'b0000_0000_0000_0000;
array[16772] <= 16'b0000_0000_0000_0000;
array[16773] <= 16'b0000_0000_0000_0000;
array[16774] <= 16'b0000_0000_0000_0000;
array[16775] <= 16'b0000_0000_0000_0000;
array[16776] <= 16'b0000_0000_0000_0000;
array[16777] <= 16'b0000_0000_0000_0000;
array[16778] <= 16'b0000_0000_0000_0000;
array[16779] <= 16'b0000_0000_0000_0000;
array[16780] <= 16'b0000_0000_0000_0000;
array[16781] <= 16'b0000_0000_0000_0000;
array[16782] <= 16'b0000_0000_0000_0000;
array[16783] <= 16'b0000_0000_0000_0000;
array[16784] <= 16'b0000_0000_0000_0000;
array[16785] <= 16'b0000_0000_0000_0000;
array[16786] <= 16'b0000_0000_0000_0000;
array[16787] <= 16'b0000_0000_0000_0000;
array[16788] <= 16'b0000_0000_0000_0000;
array[16789] <= 16'b0000_0000_0000_0000;
array[16790] <= 16'b0000_0000_0000_0000;
array[16791] <= 16'b0000_0000_0000_0000;
array[16792] <= 16'b0000_0000_0000_0000;
array[16793] <= 16'b0000_0000_0000_0000;
array[16794] <= 16'b0000_0000_0000_0000;
array[16795] <= 16'b0000_0000_0000_0000;
array[16796] <= 16'b0000_0000_0000_0000;
array[16797] <= 16'b0000_0000_0000_0000;
array[16798] <= 16'b0000_0000_0000_0000;
array[16799] <= 16'b0000_0000_0000_0000;
array[16800] <= 16'b0000_0000_0000_0000;
array[16801] <= 16'b0000_0000_0000_0000;
array[16802] <= 16'b0000_0000_0000_0000;
array[16803] <= 16'b0000_0000_0000_0000;
array[16804] <= 16'b0000_0000_0000_0000;
array[16805] <= 16'b0000_0000_0000_0000;
array[16806] <= 16'b0000_0000_0000_0000;
array[16807] <= 16'b0000_0000_0000_0000;
array[16808] <= 16'b0000_0000_0000_0000;
array[16809] <= 16'b0000_0000_0000_0000;
array[16810] <= 16'b0000_0000_0000_0000;
array[16811] <= 16'b0000_0000_0000_0000;
array[16812] <= 16'b0000_0000_0000_0000;
array[16813] <= 16'b0000_0000_0000_0000;
array[16814] <= 16'b0000_0000_0000_0000;
array[16815] <= 16'b0000_0000_0000_0000;
array[16816] <= 16'b0000_0000_0000_0000;
array[16817] <= 16'b0000_0000_0000_0000;
array[16818] <= 16'b0000_0000_0000_0000;
array[16819] <= 16'b0000_0000_0000_0000;
array[16820] <= 16'b0000_0000_0000_0000;
array[16821] <= 16'b0000_0000_0000_0000;
array[16822] <= 16'b0000_0000_0000_0000;
array[16823] <= 16'b0000_0000_0000_0000;
array[16824] <= 16'b0000_0000_0000_0000;
array[16825] <= 16'b0000_0000_0000_0000;
array[16826] <= 16'b0000_0000_0000_0000;
array[16827] <= 16'b0000_0000_0000_0000;
array[16828] <= 16'b0000_0000_0000_0000;
array[16829] <= 16'b0000_0000_0000_0000;
array[16830] <= 16'b0000_0000_0000_0000;
array[16831] <= 16'b0000_0000_0000_0000;
array[16832] <= 16'b0000_0000_0000_0000;
array[16833] <= 16'b0000_0000_0000_0000;
array[16834] <= 16'b0000_0000_0000_0000;
array[16835] <= 16'b0000_0000_0000_0000;
array[16836] <= 16'b0000_0000_0000_0000;
array[16837] <= 16'b0000_0000_0000_0000;
array[16838] <= 16'b0000_0000_0000_0000;
array[16839] <= 16'b0000_0000_0000_0000;
array[16840] <= 16'b0000_0000_0000_0000;
array[16841] <= 16'b0000_0000_0000_0000;
array[16842] <= 16'b0000_0000_0000_0000;
array[16843] <= 16'b0000_0000_0000_0000;
array[16844] <= 16'b0000_0000_0000_0000;
array[16845] <= 16'b0000_0000_0000_0000;
array[16846] <= 16'b0000_0000_0000_0000;
array[16847] <= 16'b0000_0000_0000_0000;
array[16848] <= 16'b0000_0000_0000_0000;
array[16849] <= 16'b0000_0000_0000_0000;
array[16850] <= 16'b0000_0000_0000_0000;
array[16851] <= 16'b0000_0000_0000_0000;
array[16852] <= 16'b0000_0000_0000_0000;
array[16853] <= 16'b0000_0000_0000_0000;
array[16854] <= 16'b0000_0000_0000_0000;
array[16855] <= 16'b0000_0000_0000_0000;
array[16856] <= 16'b0000_0000_0000_0000;
array[16857] <= 16'b0000_0000_0000_0000;
array[16858] <= 16'b0000_0000_0000_0000;
array[16859] <= 16'b0000_0000_0000_0000;
array[16860] <= 16'b0000_0000_0000_0000;
array[16861] <= 16'b0000_0000_0000_0000;
array[16862] <= 16'b0000_0000_0000_0000;
array[16863] <= 16'b0000_0000_0000_0000;
array[16864] <= 16'b0000_0000_0000_0000;
array[16865] <= 16'b0000_0000_0000_0000;
array[16866] <= 16'b0000_0000_0000_0000;
array[16867] <= 16'b0000_0000_0000_0000;
array[16868] <= 16'b0000_0000_0000_0000;
array[16869] <= 16'b0000_0000_0000_0000;
array[16870] <= 16'b0000_0000_0000_0000;
array[16871] <= 16'b0000_0000_0000_0000;
array[16872] <= 16'b0000_0000_0000_0000;
array[16873] <= 16'b0000_0000_0000_0000;
array[16874] <= 16'b0000_0000_0000_0000;
array[16875] <= 16'b0000_0000_0000_0000;
array[16876] <= 16'b0000_0000_0000_0000;
array[16877] <= 16'b0000_0000_0000_0000;
array[16878] <= 16'b0000_0000_0000_0000;
array[16879] <= 16'b0000_0000_0000_0000;
array[16880] <= 16'b0000_0000_0000_0000;
array[16881] <= 16'b0000_0000_0000_0000;
array[16882] <= 16'b0000_0000_0000_0000;
array[16883] <= 16'b0000_0000_0000_0000;
array[16884] <= 16'b0000_0000_0000_0000;
array[16885] <= 16'b0000_0000_0000_0000;
array[16886] <= 16'b0000_0000_0000_0000;
array[16887] <= 16'b0000_0000_0000_0000;
array[16888] <= 16'b0000_0000_0000_0000;
array[16889] <= 16'b0000_0000_0000_0000;
array[16890] <= 16'b0000_0000_0000_0000;
array[16891] <= 16'b0000_0000_0000_0000;
array[16892] <= 16'b0000_0000_0000_0000;
array[16893] <= 16'b0000_0000_0000_0000;
array[16894] <= 16'b0000_0000_0000_0000;
array[16895] <= 16'b0000_0000_0000_0000;
array[16896] <= 16'b0000_0000_0000_0000;
array[16897] <= 16'b0000_0000_0000_0000;
array[16898] <= 16'b0000_0000_0000_0000;
array[16899] <= 16'b0000_0000_0000_0000;
array[16900] <= 16'b0000_0000_0000_0000;
array[16901] <= 16'b0000_0000_0000_0000;
array[16902] <= 16'b0000_0000_0000_0000;
array[16903] <= 16'b0000_0000_0000_0000;
array[16904] <= 16'b0000_0000_0000_0000;
array[16905] <= 16'b0000_0000_0000_0000;
array[16906] <= 16'b0000_0000_0000_0000;
array[16907] <= 16'b0000_0000_0000_0000;
array[16908] <= 16'b0000_0000_0000_0000;
array[16909] <= 16'b0000_0000_0000_0000;
array[16910] <= 16'b0000_0000_0000_0000;
array[16911] <= 16'b0000_0000_0000_0000;
array[16912] <= 16'b0000_0000_0000_0000;
array[16913] <= 16'b0000_0000_0000_0000;
array[16914] <= 16'b0000_0000_0000_0000;
array[16915] <= 16'b0000_0000_0000_0000;
array[16916] <= 16'b0000_0000_0000_0000;
array[16917] <= 16'b0000_0000_0000_0000;
array[16918] <= 16'b0000_0000_0000_0000;
array[16919] <= 16'b0000_0000_0000_0000;
array[16920] <= 16'b0000_0000_0000_0000;
array[16921] <= 16'b0000_0000_0000_0000;
array[16922] <= 16'b0000_0000_0000_0000;
array[16923] <= 16'b0000_0000_0000_0000;
array[16924] <= 16'b0000_0000_0000_0000;
array[16925] <= 16'b0000_0000_0000_0000;
array[16926] <= 16'b0000_0000_0000_0000;
array[16927] <= 16'b0000_0000_0000_0000;
array[16928] <= 16'b0000_0000_0000_0000;
array[16929] <= 16'b0000_0000_0000_0000;
array[16930] <= 16'b0000_0000_0000_0000;
array[16931] <= 16'b0000_0000_0000_0000;
array[16932] <= 16'b0000_0000_0000_0000;
array[16933] <= 16'b0000_0000_0000_0000;
array[16934] <= 16'b0000_0000_0000_0000;
array[16935] <= 16'b0000_0000_0000_0000;
array[16936] <= 16'b0000_0000_0000_0000;
array[16937] <= 16'b0000_0000_0000_0000;
array[16938] <= 16'b0000_0000_0000_0000;
array[16939] <= 16'b0000_0000_0000_0000;
array[16940] <= 16'b0000_0000_0000_0000;
array[16941] <= 16'b0000_0000_0000_0000;
array[16942] <= 16'b0000_0000_0000_0000;
array[16943] <= 16'b0000_0000_0000_0000;
array[16944] <= 16'b0000_0000_0000_0000;
array[16945] <= 16'b0000_0000_0000_0000;
array[16946] <= 16'b0000_0000_0000_0000;
array[16947] <= 16'b0000_0000_0000_0000;
array[16948] <= 16'b0000_0000_0000_0000;
array[16949] <= 16'b0000_0000_0000_0000;
array[16950] <= 16'b0000_0000_0000_0000;
array[16951] <= 16'b0000_0000_0000_0000;
array[16952] <= 16'b0000_0000_0000_0000;
array[16953] <= 16'b0000_0000_0000_0000;
array[16954] <= 16'b0000_0000_0000_0000;
array[16955] <= 16'b0000_0000_0000_0000;
array[16956] <= 16'b0000_0000_0000_0000;
array[16957] <= 16'b0000_0000_0000_0000;
array[16958] <= 16'b0000_0000_0000_0000;
array[16959] <= 16'b0000_0000_0000_0000;
array[16960] <= 16'b0000_0000_0000_0000;
array[16961] <= 16'b0000_0000_0000_0000;
array[16962] <= 16'b0000_0000_0000_0000;
array[16963] <= 16'b0000_0000_0000_0000;
array[16964] <= 16'b0000_0000_0000_0000;
array[16965] <= 16'b0000_0000_0000_0000;
array[16966] <= 16'b0000_0000_0000_0000;
array[16967] <= 16'b0000_0000_0000_0000;
array[16968] <= 16'b0000_0000_0000_0000;
array[16969] <= 16'b0000_0000_0000_0000;
array[16970] <= 16'b0000_0000_0000_0000;
array[16971] <= 16'b0000_0000_0000_0000;
array[16972] <= 16'b0000_0000_0000_0000;
array[16973] <= 16'b0000_0000_0000_0000;
array[16974] <= 16'b0000_0000_0000_0000;
array[16975] <= 16'b0000_0000_0000_0000;
array[16976] <= 16'b0000_0000_0000_0000;
array[16977] <= 16'b0000_0000_0000_0000;
array[16978] <= 16'b0000_0000_0000_0000;
array[16979] <= 16'b0000_0000_0000_0000;
array[16980] <= 16'b0000_0000_0000_0000;
array[16981] <= 16'b0000_0000_0000_0000;
array[16982] <= 16'b0000_0000_0000_0000;
array[16983] <= 16'b0000_0000_0000_0000;
array[16984] <= 16'b0000_0000_0000_0000;
array[16985] <= 16'b0000_0000_0000_0000;
array[16986] <= 16'b0000_0000_0000_0000;
array[16987] <= 16'b0000_0000_0000_0000;
array[16988] <= 16'b0000_0000_0000_0000;
array[16989] <= 16'b0000_0000_0000_0000;
array[16990] <= 16'b0000_0000_0000_0000;
array[16991] <= 16'b0000_0000_0000_0000;
array[16992] <= 16'b0000_0000_0000_0000;
array[16993] <= 16'b0000_0000_0000_0000;
array[16994] <= 16'b0000_0000_0000_0000;
array[16995] <= 16'b0000_0000_0000_0000;
array[16996] <= 16'b0000_0000_0000_0000;
array[16997] <= 16'b0000_0000_0000_0000;
array[16998] <= 16'b0000_0000_0000_0000;
array[16999] <= 16'b0000_0000_0000_0000;
array[17000] <= 16'b0000_0000_0000_0000;
array[17001] <= 16'b0000_0000_0000_0000;
array[17002] <= 16'b0000_0000_0000_0000;
array[17003] <= 16'b0000_0000_0000_0000;
array[17004] <= 16'b0000_0000_0000_0000;
array[17005] <= 16'b0000_0000_0000_0000;
array[17006] <= 16'b0000_0000_0000_0000;
array[17007] <= 16'b0000_0000_0000_0000;
array[17008] <= 16'b0000_0000_0000_0000;
array[17009] <= 16'b0000_0000_0000_0000;
array[17010] <= 16'b0000_0000_0000_0000;
array[17011] <= 16'b0000_0000_0000_0000;
array[17012] <= 16'b0000_0000_0000_0000;
array[17013] <= 16'b0000_0000_0000_0000;
array[17014] <= 16'b0000_0000_0000_0000;
array[17015] <= 16'b0000_0000_0000_0000;
array[17016] <= 16'b0000_0000_0000_0000;
array[17017] <= 16'b0000_0000_0000_0000;
array[17018] <= 16'b0000_0000_0000_0000;
array[17019] <= 16'b0000_0000_0000_0000;
array[17020] <= 16'b0000_0000_0000_0000;
array[17021] <= 16'b0000_0000_0000_0000;
array[17022] <= 16'b0000_0000_0000_0000;
array[17023] <= 16'b0000_0000_0000_0000;
array[17024] <= 16'b0000_0000_0000_0000;
array[17025] <= 16'b0000_0000_0000_0000;
array[17026] <= 16'b0000_0000_0000_0000;
array[17027] <= 16'b0000_0000_0000_0000;
array[17028] <= 16'b0000_0000_0000_0000;
array[17029] <= 16'b0000_0000_0000_0000;
array[17030] <= 16'b0000_0000_0000_0000;
array[17031] <= 16'b0000_0000_0000_0000;
array[17032] <= 16'b0000_0000_0000_0000;
array[17033] <= 16'b0000_0000_0000_0000;
array[17034] <= 16'b0000_0000_0000_0000;
array[17035] <= 16'b0000_0000_0000_0000;
array[17036] <= 16'b0000_0000_0000_0000;
array[17037] <= 16'b0000_0000_0000_0000;
array[17038] <= 16'b0000_0000_0000_0000;
array[17039] <= 16'b0000_0000_0000_0000;
array[17040] <= 16'b0000_0000_0000_0000;
array[17041] <= 16'b0000_0000_0000_0000;
array[17042] <= 16'b0000_0000_0000_0000;
array[17043] <= 16'b0000_0000_0000_0000;
array[17044] <= 16'b0000_0000_0000_0000;
array[17045] <= 16'b0000_0000_0000_0000;
array[17046] <= 16'b0000_0000_0000_0000;
array[17047] <= 16'b0000_0000_0000_0000;
array[17048] <= 16'b0000_0000_0000_0000;
array[17049] <= 16'b0000_0000_0000_0000;
array[17050] <= 16'b0000_0000_0000_0000;
array[17051] <= 16'b0000_0000_0000_0000;
array[17052] <= 16'b0000_0000_0000_0000;
array[17053] <= 16'b0000_0000_0000_0000;
array[17054] <= 16'b0000_0000_0000_0000;
array[17055] <= 16'b0000_0000_0000_0000;
array[17056] <= 16'b0000_0000_0000_0000;
array[17057] <= 16'b0000_0000_0000_0000;
array[17058] <= 16'b0000_0000_0000_0000;
array[17059] <= 16'b0000_0000_0000_0000;
array[17060] <= 16'b0000_0000_0000_0000;
array[17061] <= 16'b0000_0000_0000_0000;
array[17062] <= 16'b0000_0000_0000_0000;
array[17063] <= 16'b0000_0000_0000_0000;
array[17064] <= 16'b0000_0000_0000_0000;
array[17065] <= 16'b0000_0000_0000_0000;
array[17066] <= 16'b0000_0000_0000_0000;
array[17067] <= 16'b0000_0000_0000_0000;
array[17068] <= 16'b0000_0000_0000_0000;
array[17069] <= 16'b0000_0000_0000_0000;
array[17070] <= 16'b0000_0000_0000_0000;
array[17071] <= 16'b0000_0000_0000_0000;
array[17072] <= 16'b0000_0000_0000_0000;
array[17073] <= 16'b0000_0000_0000_0000;
array[17074] <= 16'b0000_0000_0000_0000;
array[17075] <= 16'b0000_0000_0000_0000;
array[17076] <= 16'b0000_0000_0000_0000;
array[17077] <= 16'b0000_0000_0000_0000;
array[17078] <= 16'b0000_0000_0000_0000;
array[17079] <= 16'b0000_0000_0000_0000;
array[17080] <= 16'b0000_0000_0000_0000;
array[17081] <= 16'b0000_0000_0000_0000;
array[17082] <= 16'b0000_0000_0000_0000;
array[17083] <= 16'b0000_0000_0000_0000;
array[17084] <= 16'b0000_0000_0000_0000;
array[17085] <= 16'b0000_0000_0000_0000;
array[17086] <= 16'b0000_0000_0000_0000;
array[17087] <= 16'b0000_0000_0000_0000;
array[17088] <= 16'b0000_0000_0000_0000;
array[17089] <= 16'b0000_0000_0000_0000;
array[17090] <= 16'b0000_0000_0000_0000;
array[17091] <= 16'b0000_0000_0000_0000;
array[17092] <= 16'b0000_0000_0000_0000;
array[17093] <= 16'b0000_0000_0000_0000;
array[17094] <= 16'b0000_0000_0000_0000;
array[17095] <= 16'b0000_0000_0000_0000;
array[17096] <= 16'b0000_0000_0000_0000;
array[17097] <= 16'b0000_0000_0000_0000;
array[17098] <= 16'b0000_0000_0000_0000;
array[17099] <= 16'b0000_0000_0000_0000;
array[17100] <= 16'b0000_0000_0000_0000;
array[17101] <= 16'b0000_0000_0000_0000;
array[17102] <= 16'b0000_0000_0000_0000;
array[17103] <= 16'b0000_0000_0000_0000;
array[17104] <= 16'b0000_0000_0000_0000;
array[17105] <= 16'b0000_0000_0000_0000;
array[17106] <= 16'b0000_0000_0000_0000;
array[17107] <= 16'b0000_0000_0000_0000;
array[17108] <= 16'b0000_0000_0000_0000;
array[17109] <= 16'b0000_0000_0000_0000;
array[17110] <= 16'b0000_0000_0000_0000;
array[17111] <= 16'b0000_0000_0000_0000;
array[17112] <= 16'b0000_0000_0000_0000;
array[17113] <= 16'b0000_0000_0000_0000;
array[17114] <= 16'b0000_0000_0000_0000;
array[17115] <= 16'b0000_0000_0000_0000;
array[17116] <= 16'b0000_0000_0000_0000;
array[17117] <= 16'b0000_0000_0000_0000;
array[17118] <= 16'b0000_0000_0000_0000;
array[17119] <= 16'b0000_0000_0000_0000;
array[17120] <= 16'b0000_0000_0000_0000;
array[17121] <= 16'b0000_0000_0000_0000;
array[17122] <= 16'b0000_0000_0000_0000;
array[17123] <= 16'b0000_0000_0000_0000;
array[17124] <= 16'b0000_0000_0000_0000;
array[17125] <= 16'b0000_0000_0000_0000;
array[17126] <= 16'b0000_0000_0000_0000;
array[17127] <= 16'b0000_0000_0000_0000;
array[17128] <= 16'b0000_0000_0000_0000;
array[17129] <= 16'b0000_0000_0000_0000;
array[17130] <= 16'b0000_0000_0000_0000;
array[17131] <= 16'b0000_0000_0000_0000;
array[17132] <= 16'b0000_0000_0000_0000;
array[17133] <= 16'b0000_0000_0000_0000;
array[17134] <= 16'b0000_0000_0000_0000;
array[17135] <= 16'b0000_0000_0000_0000;
array[17136] <= 16'b0000_0000_0000_0000;
array[17137] <= 16'b0000_0000_0000_0000;
array[17138] <= 16'b0000_0000_0000_0000;
array[17139] <= 16'b0000_0000_0000_0000;
array[17140] <= 16'b0000_0000_0000_0000;
array[17141] <= 16'b0000_0000_0000_0000;
array[17142] <= 16'b0000_0000_0000_0000;
array[17143] <= 16'b0000_0000_0000_0000;
array[17144] <= 16'b0000_0000_0000_0000;
array[17145] <= 16'b0000_0000_0000_0000;
array[17146] <= 16'b0000_0000_0000_0000;
array[17147] <= 16'b0000_0000_0000_0000;
array[17148] <= 16'b0000_0000_0000_0000;
array[17149] <= 16'b0000_0000_0000_0000;
array[17150] <= 16'b0000_0000_0000_0000;
array[17151] <= 16'b0000_0000_0000_0000;
array[17152] <= 16'b0000_0000_0000_0000;
array[17153] <= 16'b0000_0000_0000_0000;
array[17154] <= 16'b0000_0000_0000_0000;
array[17155] <= 16'b0000_0000_0000_0000;
array[17156] <= 16'b0000_0000_0000_0000;
array[17157] <= 16'b0000_0000_0000_0000;
array[17158] <= 16'b0000_0000_0000_0000;
array[17159] <= 16'b0000_0000_0000_0000;
array[17160] <= 16'b0000_0000_0000_0000;
array[17161] <= 16'b0000_0000_0000_0000;
array[17162] <= 16'b0000_0000_0000_0000;
array[17163] <= 16'b0000_0000_0000_0000;
array[17164] <= 16'b0000_0000_0000_0000;
array[17165] <= 16'b0000_0000_0000_0000;
array[17166] <= 16'b0000_0000_0000_0000;
array[17167] <= 16'b0000_0000_0000_0000;
array[17168] <= 16'b0000_0000_0000_0000;
array[17169] <= 16'b0000_0000_0000_0000;
array[17170] <= 16'b0000_0000_0000_0000;
array[17171] <= 16'b0000_0000_0000_0000;
array[17172] <= 16'b0000_0000_0000_0000;
array[17173] <= 16'b0000_0000_0000_0000;
array[17174] <= 16'b0000_0000_0000_0000;
array[17175] <= 16'b0000_0000_0000_0000;
array[17176] <= 16'b0000_0000_0000_0000;
array[17177] <= 16'b0000_0000_0000_0000;
array[17178] <= 16'b0000_0000_0000_0000;
array[17179] <= 16'b0000_0000_0000_0000;
array[17180] <= 16'b0000_0000_0000_0000;
array[17181] <= 16'b0000_0000_0000_0000;
array[17182] <= 16'b0000_0000_0000_0000;
array[17183] <= 16'b0000_0000_0000_0000;
array[17184] <= 16'b0000_0000_0000_0000;
array[17185] <= 16'b0000_0000_0000_0000;
array[17186] <= 16'b0000_0000_0000_0000;
array[17187] <= 16'b0000_0000_0000_0000;
array[17188] <= 16'b0000_0000_0000_0000;
array[17189] <= 16'b0000_0000_0000_0000;
array[17190] <= 16'b0000_0000_0000_0000;
array[17191] <= 16'b0000_0000_0000_0000;
array[17192] <= 16'b0000_0000_0000_0000;
array[17193] <= 16'b0000_0000_0000_0000;
array[17194] <= 16'b0000_0000_0000_0000;
array[17195] <= 16'b0000_0000_0000_0000;
array[17196] <= 16'b0000_0000_0000_0000;
array[17197] <= 16'b0000_0000_0000_0000;
array[17198] <= 16'b0000_0000_0000_0000;
array[17199] <= 16'b0000_0000_0000_0000;
array[17200] <= 16'b0000_0000_0000_0000;
array[17201] <= 16'b0000_0000_0000_0000;
array[17202] <= 16'b0000_0000_0000_0000;
array[17203] <= 16'b0000_0000_0000_0000;
array[17204] <= 16'b0000_0000_0000_0000;
array[17205] <= 16'b0000_0000_0000_0000;
array[17206] <= 16'b0000_0000_0000_0000;
array[17207] <= 16'b0000_0000_0000_0000;
array[17208] <= 16'b0000_0000_0000_0000;
array[17209] <= 16'b0000_0000_0000_0000;
array[17210] <= 16'b0000_0000_0000_0000;
array[17211] <= 16'b0000_0000_0000_0000;
array[17212] <= 16'b0000_0000_0000_0000;
array[17213] <= 16'b0000_0000_0000_0000;
array[17214] <= 16'b0000_0000_0000_0000;
array[17215] <= 16'b0000_0000_0000_0000;
array[17216] <= 16'b0000_0000_0000_0000;
array[17217] <= 16'b0000_0000_0000_0000;
array[17218] <= 16'b0000_0000_0000_0000;
array[17219] <= 16'b0000_0000_0000_0000;
array[17220] <= 16'b0000_0000_0000_0000;
array[17221] <= 16'b0000_0000_0000_0000;
array[17222] <= 16'b0000_0000_0000_0000;
array[17223] <= 16'b0000_0000_0000_0000;
array[17224] <= 16'b0000_0000_0000_0000;
array[17225] <= 16'b0000_0000_0000_0000;
array[17226] <= 16'b0000_0000_0000_0000;
array[17227] <= 16'b0000_0000_0000_0000;
array[17228] <= 16'b0000_0000_0000_0000;
array[17229] <= 16'b0000_0000_0000_0000;
array[17230] <= 16'b0000_0000_0000_0000;
array[17231] <= 16'b0000_0000_0000_0000;
array[17232] <= 16'b0000_0000_0000_0000;
array[17233] <= 16'b0000_0000_0000_0000;
array[17234] <= 16'b0000_0000_0000_0000;
array[17235] <= 16'b0000_0000_0000_0000;
array[17236] <= 16'b0000_0000_0000_0000;
array[17237] <= 16'b0000_0000_0000_0000;
array[17238] <= 16'b0000_0000_0000_0000;
array[17239] <= 16'b0000_0000_0000_0000;
array[17240] <= 16'b0000_0000_0000_0000;
array[17241] <= 16'b0000_0000_0000_0000;
array[17242] <= 16'b0000_0000_0000_0000;
array[17243] <= 16'b0000_0000_0000_0000;
array[17244] <= 16'b0000_0000_0000_0000;
array[17245] <= 16'b0000_0000_0000_0000;
array[17246] <= 16'b0000_0000_0000_0000;
array[17247] <= 16'b0000_0000_0000_0000;
array[17248] <= 16'b0000_0000_0000_0000;
array[17249] <= 16'b0000_0000_0000_0000;
array[17250] <= 16'b0000_0000_0000_0000;
array[17251] <= 16'b0000_0000_0000_0000;
array[17252] <= 16'b0000_0000_0000_0000;
array[17253] <= 16'b0000_0000_0000_0000;
array[17254] <= 16'b0000_0000_0000_0000;
array[17255] <= 16'b0000_0000_0000_0000;
array[17256] <= 16'b0000_0000_0000_0000;
array[17257] <= 16'b0000_0000_0000_0000;
array[17258] <= 16'b0000_0000_0000_0000;
array[17259] <= 16'b0000_0000_0000_0000;
array[17260] <= 16'b0000_0000_0000_0000;
array[17261] <= 16'b0000_0000_0000_0000;
array[17262] <= 16'b0000_0000_0000_0000;
array[17263] <= 16'b0000_0000_0000_0000;
array[17264] <= 16'b0000_0000_0000_0000;
array[17265] <= 16'b0000_0000_0000_0000;
array[17266] <= 16'b0000_0000_0000_0000;
array[17267] <= 16'b0000_0000_0000_0000;
array[17268] <= 16'b0000_0000_0000_0000;
array[17269] <= 16'b0000_0000_0000_0000;
array[17270] <= 16'b0000_0000_0000_0000;
array[17271] <= 16'b0000_0000_0000_0000;
array[17272] <= 16'b0000_0000_0000_0000;
array[17273] <= 16'b0000_0000_0000_0000;
array[17274] <= 16'b0000_0000_0000_0000;
array[17275] <= 16'b0000_0000_0000_0000;
array[17276] <= 16'b0000_0000_0000_0000;
array[17277] <= 16'b0000_0000_0000_0000;
array[17278] <= 16'b0000_0000_0000_0000;
array[17279] <= 16'b0000_0000_0000_0000;
array[17280] <= 16'b0000_0000_0000_0000;
array[17281] <= 16'b0000_0000_0000_0000;
array[17282] <= 16'b0000_0000_0000_0000;
array[17283] <= 16'b0000_0000_0000_0000;
array[17284] <= 16'b0000_0000_0000_0000;
array[17285] <= 16'b0000_0000_0000_0000;
array[17286] <= 16'b0000_0000_0000_0000;
array[17287] <= 16'b0000_0000_0000_0000;
array[17288] <= 16'b0000_0000_0000_0000;
array[17289] <= 16'b0000_0000_0000_0000;
array[17290] <= 16'b0000_0000_0000_0000;
array[17291] <= 16'b0000_0000_0000_0000;
array[17292] <= 16'b0000_0000_0000_0000;
array[17293] <= 16'b0000_0000_0000_0000;
array[17294] <= 16'b0000_0000_0000_0000;
array[17295] <= 16'b0000_0000_0000_0000;
array[17296] <= 16'b0000_0000_0000_0000;
array[17297] <= 16'b0000_0000_0000_0000;
array[17298] <= 16'b0000_0000_0000_0000;
array[17299] <= 16'b0000_0000_0000_0000;
array[17300] <= 16'b0000_0000_0000_0000;
array[17301] <= 16'b0000_0000_0000_0000;
array[17302] <= 16'b0000_0000_0000_0000;
array[17303] <= 16'b0000_0000_0000_0000;
array[17304] <= 16'b0000_0000_0000_0000;
array[17305] <= 16'b0000_0000_0000_0000;
array[17306] <= 16'b0000_0000_0000_0000;
array[17307] <= 16'b0000_0000_0000_0000;
array[17308] <= 16'b0000_0000_0000_0000;
array[17309] <= 16'b0000_0000_0000_0000;
array[17310] <= 16'b0000_0000_0000_0000;
array[17311] <= 16'b0000_0000_0000_0000;
array[17312] <= 16'b0000_0000_0000_0000;
array[17313] <= 16'b0000_0000_0000_0000;
array[17314] <= 16'b0000_0000_0000_0000;
array[17315] <= 16'b0000_0000_0000_0000;
array[17316] <= 16'b0000_0000_0000_0000;
array[17317] <= 16'b0000_0000_0000_0000;
array[17318] <= 16'b0000_0000_0000_0000;
array[17319] <= 16'b0000_0000_0000_0000;
array[17320] <= 16'b0000_0000_0000_0000;
array[17321] <= 16'b0000_0000_0000_0000;
array[17322] <= 16'b0000_0000_0000_0000;
array[17323] <= 16'b0000_0000_0000_0000;
array[17324] <= 16'b0000_0000_0000_0000;
array[17325] <= 16'b0000_0000_0000_0000;
array[17326] <= 16'b0000_0000_0000_0000;
array[17327] <= 16'b0000_0000_0000_0000;
array[17328] <= 16'b0000_0000_0000_0000;
array[17329] <= 16'b0000_0000_0000_0000;
array[17330] <= 16'b0000_0000_0000_0000;
array[17331] <= 16'b0000_0000_0000_0000;
array[17332] <= 16'b0000_0000_0000_0000;
array[17333] <= 16'b0000_0000_0000_0000;
array[17334] <= 16'b0000_0000_0000_0000;
array[17335] <= 16'b0000_0000_0000_0000;
array[17336] <= 16'b0000_0000_0000_0000;
array[17337] <= 16'b0000_0000_0000_0000;
array[17338] <= 16'b0000_0000_0000_0000;
array[17339] <= 16'b0000_0000_0000_0000;
array[17340] <= 16'b0000_0000_0000_0000;
array[17341] <= 16'b0000_0000_0000_0000;
array[17342] <= 16'b0000_0000_0000_0000;
array[17343] <= 16'b0000_0000_0000_0000;
array[17344] <= 16'b0000_0000_0000_0000;
array[17345] <= 16'b0000_0000_0000_0000;
array[17346] <= 16'b0000_0000_0000_0000;
array[17347] <= 16'b0000_0000_0000_0000;
array[17348] <= 16'b0000_0000_0000_0000;
array[17349] <= 16'b0000_0000_0000_0000;
array[17350] <= 16'b0000_0000_0000_0000;
array[17351] <= 16'b0000_0000_0000_0000;
array[17352] <= 16'b0000_0000_0000_0000;
array[17353] <= 16'b0000_0000_0000_0000;
array[17354] <= 16'b0000_0000_0000_0000;
array[17355] <= 16'b0000_0000_0000_0000;
array[17356] <= 16'b0000_0000_0000_0000;
array[17357] <= 16'b0000_0000_0000_0000;
array[17358] <= 16'b0000_0000_0000_0000;
array[17359] <= 16'b0000_0000_0000_0000;
array[17360] <= 16'b0000_0000_0000_0000;
array[17361] <= 16'b0000_0000_0000_0000;
array[17362] <= 16'b0000_0000_0000_0000;
array[17363] <= 16'b0000_0000_0000_0000;
array[17364] <= 16'b0000_0000_0000_0000;
array[17365] <= 16'b0000_0000_0000_0000;
array[17366] <= 16'b0000_0000_0000_0000;
array[17367] <= 16'b0000_0000_0000_0000;
array[17368] <= 16'b0000_0000_0000_0000;
array[17369] <= 16'b0000_0000_0000_0000;
array[17370] <= 16'b0000_0000_0000_0000;
array[17371] <= 16'b0000_0000_0000_0000;
array[17372] <= 16'b0000_0000_0000_0000;
array[17373] <= 16'b0000_0000_0000_0000;
array[17374] <= 16'b0000_0000_0000_0000;
array[17375] <= 16'b0000_0000_0000_0000;
array[17376] <= 16'b0000_0000_0000_0000;
array[17377] <= 16'b0000_0000_0000_0000;
array[17378] <= 16'b0000_0000_0000_0000;
array[17379] <= 16'b0000_0000_0000_0000;
array[17380] <= 16'b0000_0000_0000_0000;
array[17381] <= 16'b0000_0000_0000_0000;
array[17382] <= 16'b0000_0000_0000_0000;
array[17383] <= 16'b0000_0000_0000_0000;
array[17384] <= 16'b0000_0000_0000_0000;
array[17385] <= 16'b0000_0000_0000_0000;
array[17386] <= 16'b0000_0000_0000_0000;
array[17387] <= 16'b0000_0000_0000_0000;
array[17388] <= 16'b0000_0000_0000_0000;
array[17389] <= 16'b0000_0000_0000_0000;
array[17390] <= 16'b0000_0000_0000_0000;
array[17391] <= 16'b0000_0000_0000_0000;
array[17392] <= 16'b0000_0000_0000_0000;
array[17393] <= 16'b0000_0000_0000_0000;
array[17394] <= 16'b0000_0000_0000_0000;
array[17395] <= 16'b0000_0000_0000_0000;
array[17396] <= 16'b0000_0000_0000_0000;
array[17397] <= 16'b0000_0000_0000_0000;
array[17398] <= 16'b0000_0000_0000_0000;
array[17399] <= 16'b0000_0000_0000_0000;
array[17400] <= 16'b0000_0000_0000_0000;
array[17401] <= 16'b0000_0000_0000_0000;
array[17402] <= 16'b0000_0000_0000_0000;
array[17403] <= 16'b0000_0000_0000_0000;
array[17404] <= 16'b0000_0000_0000_0000;
array[17405] <= 16'b0000_0000_0000_0000;
array[17406] <= 16'b0000_0000_0000_0000;
array[17407] <= 16'b0000_0000_0000_0000;
array[17408] <= 16'b0000_0000_0000_0000;
array[17409] <= 16'b0000_0000_0000_0000;
array[17410] <= 16'b0000_0000_0000_0000;
array[17411] <= 16'b0000_0000_0000_0000;
array[17412] <= 16'b0000_0000_0000_0000;
array[17413] <= 16'b0000_0000_0000_0000;
array[17414] <= 16'b0000_0000_0000_0000;
array[17415] <= 16'b0000_0000_0000_0000;
array[17416] <= 16'b0000_0000_0000_0000;
array[17417] <= 16'b0000_0000_0000_0000;
array[17418] <= 16'b0000_0000_0000_0000;
array[17419] <= 16'b0000_0000_0000_0000;
array[17420] <= 16'b0000_0000_0000_0000;
array[17421] <= 16'b0000_0000_0000_0000;
array[17422] <= 16'b0000_0000_0000_0000;
array[17423] <= 16'b0000_0000_0000_0000;
array[17424] <= 16'b0000_0000_0000_0000;
array[17425] <= 16'b0000_0000_0000_0000;
array[17426] <= 16'b0000_0000_0000_0000;
array[17427] <= 16'b0000_0000_0000_0000;
array[17428] <= 16'b0000_0000_0000_0000;
array[17429] <= 16'b0000_0000_0000_0000;
array[17430] <= 16'b0000_0000_0000_0000;
array[17431] <= 16'b0000_0000_0000_0000;
array[17432] <= 16'b0000_0000_0000_0000;
array[17433] <= 16'b0000_0000_0000_0000;
array[17434] <= 16'b0000_0000_0000_0000;
array[17435] <= 16'b0000_0000_0000_0000;
array[17436] <= 16'b0000_0000_0000_0000;
array[17437] <= 16'b0000_0000_0000_0000;
array[17438] <= 16'b0000_0000_0000_0000;
array[17439] <= 16'b0000_0000_0000_0000;
array[17440] <= 16'b0000_0000_0000_0000;
array[17441] <= 16'b0000_0000_0000_0000;
array[17442] <= 16'b0000_0000_0000_0000;
array[17443] <= 16'b0000_0000_0000_0000;
array[17444] <= 16'b0000_0000_0000_0000;
array[17445] <= 16'b0000_0000_0000_0000;
array[17446] <= 16'b0000_0000_0000_0000;
array[17447] <= 16'b0000_0000_0000_0000;
array[17448] <= 16'b0000_0000_0000_0000;
array[17449] <= 16'b0000_0000_0000_0000;
array[17450] <= 16'b0000_0000_0000_0000;
array[17451] <= 16'b0000_0000_0000_0000;
array[17452] <= 16'b0000_0000_0000_0000;
array[17453] <= 16'b0000_0000_0000_0000;
array[17454] <= 16'b0000_0000_0000_0000;
array[17455] <= 16'b0000_0000_0000_0000;
array[17456] <= 16'b0000_0000_0000_0000;
array[17457] <= 16'b0000_0000_0000_0000;
array[17458] <= 16'b0000_0000_0000_0000;
array[17459] <= 16'b0000_0000_0000_0000;
array[17460] <= 16'b0000_0000_0000_0000;
array[17461] <= 16'b0000_0000_0000_0000;
array[17462] <= 16'b0000_0000_0000_0000;
array[17463] <= 16'b0000_0000_0000_0000;
array[17464] <= 16'b0000_0000_0000_0000;
array[17465] <= 16'b0000_0000_0000_0000;
array[17466] <= 16'b0000_0000_0000_0000;
array[17467] <= 16'b0000_0000_0000_0000;
array[17468] <= 16'b0000_0000_0000_0000;
array[17469] <= 16'b0000_0000_0000_0000;
array[17470] <= 16'b0000_0000_0000_0000;
array[17471] <= 16'b0000_0000_0000_0000;
array[17472] <= 16'b0000_0000_0000_0000;
array[17473] <= 16'b0000_0000_0000_0000;
array[17474] <= 16'b0000_0000_0000_0000;
array[17475] <= 16'b0000_0000_0000_0000;
array[17476] <= 16'b0000_0000_0000_0000;
array[17477] <= 16'b0000_0000_0000_0000;
array[17478] <= 16'b0000_0000_0000_0000;
array[17479] <= 16'b0000_0000_0000_0000;
array[17480] <= 16'b0000_0000_0000_0000;
array[17481] <= 16'b0000_0000_0000_0000;
array[17482] <= 16'b0000_0000_0000_0000;
array[17483] <= 16'b0000_0000_0000_0000;
array[17484] <= 16'b0000_0000_0000_0000;
array[17485] <= 16'b0000_0000_0000_0000;
array[17486] <= 16'b0000_0000_0000_0000;
array[17487] <= 16'b0000_0000_0000_0000;
array[17488] <= 16'b0000_0000_0000_0000;
array[17489] <= 16'b0000_0000_0000_0000;
array[17490] <= 16'b0000_0000_0000_0000;
array[17491] <= 16'b0000_0000_0000_0000;
array[17492] <= 16'b0000_0000_0000_0000;
array[17493] <= 16'b0000_0000_0000_0000;
array[17494] <= 16'b0000_0000_0000_0000;
array[17495] <= 16'b0000_0000_0000_0000;
array[17496] <= 16'b0000_0000_0000_0000;
array[17497] <= 16'b0000_0000_0000_0000;
array[17498] <= 16'b0000_0000_0000_0000;
array[17499] <= 16'b0000_0000_0000_0000;
array[17500] <= 16'b0000_0000_0000_0000;
array[17501] <= 16'b0000_0000_0000_0000;
array[17502] <= 16'b0000_0000_0000_0000;
array[17503] <= 16'b0000_0000_0000_0000;
array[17504] <= 16'b0000_0000_0000_0000;
array[17505] <= 16'b0000_0000_0000_0000;
array[17506] <= 16'b0000_0000_0000_0000;
array[17507] <= 16'b0000_0000_0000_0000;
array[17508] <= 16'b0000_0000_0000_0000;
array[17509] <= 16'b0000_0000_0000_0000;
array[17510] <= 16'b0000_0000_0000_0000;
array[17511] <= 16'b0000_0000_0000_0000;
array[17512] <= 16'b0000_0000_0000_0000;
array[17513] <= 16'b0000_0000_0000_0000;
array[17514] <= 16'b0000_0000_0000_0000;
array[17515] <= 16'b0000_0000_0000_0000;
array[17516] <= 16'b0000_0000_0000_0000;
array[17517] <= 16'b0000_0000_0000_0000;
array[17518] <= 16'b0000_0000_0000_0000;
array[17519] <= 16'b0000_0000_0000_0000;
array[17520] <= 16'b0000_0000_0000_0000;
array[17521] <= 16'b0000_0000_0000_0000;
array[17522] <= 16'b0000_0000_0000_0000;
array[17523] <= 16'b0000_0000_0000_0000;
array[17524] <= 16'b0000_0000_0000_0000;
array[17525] <= 16'b0000_0000_0000_0000;
array[17526] <= 16'b0000_0000_0000_0000;
array[17527] <= 16'b0000_0000_0000_0000;
array[17528] <= 16'b0000_0000_0000_0000;
array[17529] <= 16'b0000_0000_0000_0000;
array[17530] <= 16'b0000_0000_0000_0000;
array[17531] <= 16'b0000_0000_0000_0000;
array[17532] <= 16'b0000_0000_0000_0000;
array[17533] <= 16'b0000_0000_0000_0000;
array[17534] <= 16'b0000_0000_0000_0000;
array[17535] <= 16'b0000_0000_0000_0000;
array[17536] <= 16'b0000_0000_0000_0000;
array[17537] <= 16'b0000_0000_0000_0000;
array[17538] <= 16'b0000_0000_0000_0000;
array[17539] <= 16'b0000_0000_0000_0000;
array[17540] <= 16'b0000_0000_0000_0000;
array[17541] <= 16'b0000_0000_0000_0000;
array[17542] <= 16'b0000_0000_0000_0000;
array[17543] <= 16'b0000_0000_0000_0000;
array[17544] <= 16'b0000_0000_0000_0000;
array[17545] <= 16'b0000_0000_0000_0000;
array[17546] <= 16'b0000_0000_0000_0000;
array[17547] <= 16'b0000_0000_0000_0000;
array[17548] <= 16'b0000_0000_0000_0000;
array[17549] <= 16'b0000_0000_0000_0000;
array[17550] <= 16'b0000_0000_0000_0000;
array[17551] <= 16'b0000_0000_0000_0000;
array[17552] <= 16'b0000_0000_0000_0000;
array[17553] <= 16'b0000_0000_0000_0000;
array[17554] <= 16'b0000_0000_0000_0000;
array[17555] <= 16'b0000_0000_0000_0000;
array[17556] <= 16'b0000_0000_0000_0000;
array[17557] <= 16'b0000_0000_0000_0000;
array[17558] <= 16'b0000_0000_0000_0000;
array[17559] <= 16'b0000_0000_0000_0000;
array[17560] <= 16'b0000_0000_0000_0000;
array[17561] <= 16'b0000_0000_0000_0000;
array[17562] <= 16'b0000_0000_0000_0000;
array[17563] <= 16'b0000_0000_0000_0000;
array[17564] <= 16'b0000_0000_0000_0000;
array[17565] <= 16'b0000_0000_0000_0000;
array[17566] <= 16'b0000_0000_0000_0000;
array[17567] <= 16'b0000_0000_0000_0000;
array[17568] <= 16'b0000_0000_0000_0000;
array[17569] <= 16'b0000_0000_0000_0000;
array[17570] <= 16'b0000_0000_0000_0000;
array[17571] <= 16'b0000_0000_0000_0000;
array[17572] <= 16'b0000_0000_0000_0000;
array[17573] <= 16'b0000_0000_0000_0000;
array[17574] <= 16'b0000_0000_0000_0000;
array[17575] <= 16'b0000_0000_0000_0000;
array[17576] <= 16'b0000_0000_0000_0000;
array[17577] <= 16'b0000_0000_0000_0000;
array[17578] <= 16'b0000_0000_0000_0000;
array[17579] <= 16'b0000_0000_0000_0000;
array[17580] <= 16'b0000_0000_0000_0000;
array[17581] <= 16'b0000_0000_0000_0000;
array[17582] <= 16'b0000_0000_0000_0000;
array[17583] <= 16'b0000_0000_0000_0000;
array[17584] <= 16'b0000_0000_0000_0000;
array[17585] <= 16'b0000_0000_0000_0000;
array[17586] <= 16'b0000_0000_0000_0000;
array[17587] <= 16'b0000_0000_0000_0000;
array[17588] <= 16'b0000_0000_0000_0000;
array[17589] <= 16'b0000_0000_0000_0000;
array[17590] <= 16'b0000_0000_0000_0000;
array[17591] <= 16'b0000_0000_0000_0000;
array[17592] <= 16'b0000_0000_0000_0000;
array[17593] <= 16'b0000_0000_0000_0000;
array[17594] <= 16'b0000_0000_0000_0000;
array[17595] <= 16'b0000_0000_0000_0000;
array[17596] <= 16'b0000_0000_0000_0000;
array[17597] <= 16'b0000_0000_0000_0000;
array[17598] <= 16'b0000_0000_0000_0000;
array[17599] <= 16'b0000_0000_0000_0000;
array[17600] <= 16'b0000_0000_0000_0000;
array[17601] <= 16'b0000_0000_0000_0000;
array[17602] <= 16'b0000_0000_0000_0000;
array[17603] <= 16'b0000_0000_0000_0000;
array[17604] <= 16'b0000_0000_0000_0000;
array[17605] <= 16'b0000_0000_0000_0000;
array[17606] <= 16'b0000_0000_0000_0000;
array[17607] <= 16'b0000_0000_0000_0000;
array[17608] <= 16'b0000_0000_0000_0000;
array[17609] <= 16'b0000_0000_0000_0000;
array[17610] <= 16'b0000_0000_0000_0000;
array[17611] <= 16'b0000_0000_0000_0000;
array[17612] <= 16'b0000_0000_0000_0000;
array[17613] <= 16'b0000_0000_0000_0000;
array[17614] <= 16'b0000_0000_0000_0000;
array[17615] <= 16'b0000_0000_0000_0000;
array[17616] <= 16'b0000_0000_0000_0000;
array[17617] <= 16'b0000_0000_0000_0000;
array[17618] <= 16'b0000_0000_0000_0000;
array[17619] <= 16'b0000_0000_0000_0000;
array[17620] <= 16'b0000_0000_0000_0000;
array[17621] <= 16'b0000_0000_0000_0000;
array[17622] <= 16'b0000_0000_0000_0000;
array[17623] <= 16'b0000_0000_0000_0000;
array[17624] <= 16'b0000_0000_0000_0000;
array[17625] <= 16'b0000_0000_0000_0000;
array[17626] <= 16'b0000_0000_0000_0000;
array[17627] <= 16'b0000_0000_0000_0000;
array[17628] <= 16'b0000_0000_0000_0000;
array[17629] <= 16'b0000_0000_0000_0000;
array[17630] <= 16'b0000_0000_0000_0000;
array[17631] <= 16'b0000_0000_0000_0000;
array[17632] <= 16'b0000_0000_0000_0000;
array[17633] <= 16'b0000_0000_0000_0000;
array[17634] <= 16'b0000_0000_0000_0000;
array[17635] <= 16'b0000_0000_0000_0000;
array[17636] <= 16'b0000_0000_0000_0000;
array[17637] <= 16'b0000_0000_0000_0000;
array[17638] <= 16'b0000_0000_0000_0000;
array[17639] <= 16'b0000_0000_0000_0000;
array[17640] <= 16'b0000_0000_0000_0000;
array[17641] <= 16'b0000_0000_0000_0000;
array[17642] <= 16'b0000_0000_0000_0000;
array[17643] <= 16'b0000_0000_0000_0000;
array[17644] <= 16'b0000_0000_0000_0000;
array[17645] <= 16'b0000_0000_0000_0000;
array[17646] <= 16'b0000_0000_0000_0000;
array[17647] <= 16'b0000_0000_0000_0000;
array[17648] <= 16'b0000_0000_0000_0000;
array[17649] <= 16'b0000_0000_0000_0000;
array[17650] <= 16'b0000_0000_0000_0000;
array[17651] <= 16'b0000_0000_0000_0000;
array[17652] <= 16'b0000_0000_0000_0000;
array[17653] <= 16'b0000_0000_0000_0000;
array[17654] <= 16'b0000_0000_0000_0000;
array[17655] <= 16'b0000_0000_0000_0000;
array[17656] <= 16'b0000_0000_0000_0000;
array[17657] <= 16'b0000_0000_0000_0000;
array[17658] <= 16'b0000_0000_0000_0000;
array[17659] <= 16'b0000_0000_0000_0000;
array[17660] <= 16'b0000_0000_0000_0000;
array[17661] <= 16'b0000_0000_0000_0000;
array[17662] <= 16'b0000_0000_0000_0000;
array[17663] <= 16'b0000_0000_0000_0000;
array[17664] <= 16'b0000_0000_0000_0000;
array[17665] <= 16'b0000_0000_0000_0000;
array[17666] <= 16'b0000_0000_0000_0000;
array[17667] <= 16'b0000_0000_0000_0000;
array[17668] <= 16'b0000_0000_0000_0000;
array[17669] <= 16'b0000_0000_0000_0000;
array[17670] <= 16'b0000_0000_0000_0000;
array[17671] <= 16'b0000_0000_0000_0000;
array[17672] <= 16'b0000_0000_0000_0000;
array[17673] <= 16'b0000_0000_0000_0000;
array[17674] <= 16'b0000_0000_0000_0000;
array[17675] <= 16'b0000_0000_0000_0000;
array[17676] <= 16'b0000_0000_0000_0000;
array[17677] <= 16'b0000_0000_0000_0000;
array[17678] <= 16'b0000_0000_0000_0000;
array[17679] <= 16'b0000_0000_0000_0000;
array[17680] <= 16'b0000_0000_0000_0000;
array[17681] <= 16'b0000_0000_0000_0000;
array[17682] <= 16'b0000_0000_0000_0000;
array[17683] <= 16'b0000_0000_0000_0000;
array[17684] <= 16'b0000_0000_0000_0000;
array[17685] <= 16'b0000_0000_0000_0000;
array[17686] <= 16'b0000_0000_0000_0000;
array[17687] <= 16'b0000_0000_0000_0000;
array[17688] <= 16'b0000_0000_0000_0000;
array[17689] <= 16'b0000_0000_0000_0000;
array[17690] <= 16'b0000_0000_0000_0000;
array[17691] <= 16'b0000_0000_0000_0000;
array[17692] <= 16'b0000_0000_0000_0000;
array[17693] <= 16'b0000_0000_0000_0000;
array[17694] <= 16'b0000_0000_0000_0000;
array[17695] <= 16'b0000_0000_0000_0000;
array[17696] <= 16'b0000_0000_0000_0000;
array[17697] <= 16'b0000_0000_0000_0000;
array[17698] <= 16'b0000_0000_0000_0000;
array[17699] <= 16'b0000_0000_0000_0000;
array[17700] <= 16'b0000_0000_0000_0000;
array[17701] <= 16'b0000_0000_0000_0000;
array[17702] <= 16'b0000_0000_0000_0000;
array[17703] <= 16'b0000_0000_0000_0000;
array[17704] <= 16'b0000_0000_0000_0000;
array[17705] <= 16'b0000_0000_0000_0000;
array[17706] <= 16'b0000_0000_0000_0000;
array[17707] <= 16'b0000_0000_0000_0000;
array[17708] <= 16'b0000_0000_0000_0000;
array[17709] <= 16'b0000_0000_0000_0000;
array[17710] <= 16'b0000_0000_0000_0000;
array[17711] <= 16'b0000_0000_0000_0000;
array[17712] <= 16'b0000_0000_0000_0000;
array[17713] <= 16'b0000_0000_0000_0000;
array[17714] <= 16'b0000_0000_0000_0000;
array[17715] <= 16'b0000_0000_0000_0000;
array[17716] <= 16'b0000_0000_0000_0000;
array[17717] <= 16'b0000_0000_0000_0000;
array[17718] <= 16'b0000_0000_0000_0000;
array[17719] <= 16'b0000_0000_0000_0000;
array[17720] <= 16'b0000_0000_0000_0000;
array[17721] <= 16'b0000_0000_0000_0000;
array[17722] <= 16'b0000_0000_0000_0000;
array[17723] <= 16'b0000_0000_0000_0000;
array[17724] <= 16'b0000_0000_0000_0000;
array[17725] <= 16'b0000_0000_0000_0000;
array[17726] <= 16'b0000_0000_0000_0000;
array[17727] <= 16'b0000_0000_0000_0000;
array[17728] <= 16'b0000_0000_0000_0000;
array[17729] <= 16'b0000_0000_0000_0000;
array[17730] <= 16'b0000_0000_0000_0000;
array[17731] <= 16'b0000_0000_0000_0000;
array[17732] <= 16'b0000_0000_0000_0000;
array[17733] <= 16'b0000_0000_0000_0000;
array[17734] <= 16'b0000_0000_0000_0000;
array[17735] <= 16'b0000_0000_0000_0000;
array[17736] <= 16'b0000_0000_0000_0000;
array[17737] <= 16'b0000_0000_0000_0000;
array[17738] <= 16'b0000_0000_0000_0000;
array[17739] <= 16'b0000_0000_0000_0000;
array[17740] <= 16'b0000_0000_0000_0000;
array[17741] <= 16'b0000_0000_0000_0000;
array[17742] <= 16'b0000_0000_0000_0000;
array[17743] <= 16'b0000_0000_0000_0000;
array[17744] <= 16'b0000_0000_0000_0000;
array[17745] <= 16'b0000_0000_0000_0000;
array[17746] <= 16'b0000_0000_0000_0000;
array[17747] <= 16'b0000_0000_0000_0000;
array[17748] <= 16'b0000_0000_0000_0000;
array[17749] <= 16'b0000_0000_0000_0000;
array[17750] <= 16'b0000_0000_0000_0000;
array[17751] <= 16'b0000_0000_0000_0000;
array[17752] <= 16'b0000_0000_0000_0000;
array[17753] <= 16'b0000_0000_0000_0000;
array[17754] <= 16'b0000_0000_0000_0000;
array[17755] <= 16'b0000_0000_0000_0000;
array[17756] <= 16'b0000_0000_0000_0000;
array[17757] <= 16'b0000_0000_0000_0000;
array[17758] <= 16'b0000_0000_0000_0000;
array[17759] <= 16'b0000_0000_0000_0000;
array[17760] <= 16'b0000_0000_0000_0000;
array[17761] <= 16'b0000_0000_0000_0000;
array[17762] <= 16'b0000_0000_0000_0000;
array[17763] <= 16'b0000_0000_0000_0000;
array[17764] <= 16'b0000_0000_0000_0000;
array[17765] <= 16'b0000_0000_0000_0000;
array[17766] <= 16'b0000_0000_0000_0000;
array[17767] <= 16'b0000_0000_0000_0000;
array[17768] <= 16'b0000_0000_0000_0000;
array[17769] <= 16'b0000_0000_0000_0000;
array[17770] <= 16'b0000_0000_0000_0000;
array[17771] <= 16'b0000_0000_0000_0000;
array[17772] <= 16'b0000_0000_0000_0000;
array[17773] <= 16'b0000_0000_0000_0000;
array[17774] <= 16'b0000_0000_0000_0000;
array[17775] <= 16'b0000_0000_0000_0000;
array[17776] <= 16'b0000_0000_0000_0000;
array[17777] <= 16'b0000_0000_0000_0000;
array[17778] <= 16'b0000_0000_0000_0000;
array[17779] <= 16'b0000_0000_0000_0000;
array[17780] <= 16'b0000_0000_0000_0000;
array[17781] <= 16'b0000_0000_0000_0000;
array[17782] <= 16'b0000_0000_0000_0000;
array[17783] <= 16'b0000_0000_0000_0000;
array[17784] <= 16'b0000_0000_0000_0000;
array[17785] <= 16'b0000_0000_0000_0000;
array[17786] <= 16'b0000_0000_0000_0000;
array[17787] <= 16'b0000_0000_0000_0000;
array[17788] <= 16'b0000_0000_0000_0000;
array[17789] <= 16'b0000_0000_0000_0000;
array[17790] <= 16'b0000_0000_0000_0000;
array[17791] <= 16'b0000_0000_0000_0000;
array[17792] <= 16'b0000_0000_0000_0000;
array[17793] <= 16'b0000_0000_0000_0000;
array[17794] <= 16'b0000_0000_0000_0000;
array[17795] <= 16'b0000_0000_0000_0000;
array[17796] <= 16'b0000_0000_0000_0000;
array[17797] <= 16'b0000_0000_0000_0000;
array[17798] <= 16'b0000_0000_0000_0000;
array[17799] <= 16'b0000_0000_0000_0000;
array[17800] <= 16'b0000_0000_0000_0000;
array[17801] <= 16'b0000_0000_0000_0000;
array[17802] <= 16'b0000_0000_0000_0000;
array[17803] <= 16'b0000_0000_0000_0000;
array[17804] <= 16'b0000_0000_0000_0000;
array[17805] <= 16'b0000_0000_0000_0000;
array[17806] <= 16'b0000_0000_0000_0000;
array[17807] <= 16'b0000_0000_0000_0000;
array[17808] <= 16'b0000_0000_0000_0000;
array[17809] <= 16'b0000_0000_0000_0000;
array[17810] <= 16'b0000_0000_0000_0000;
array[17811] <= 16'b0000_0000_0000_0000;
array[17812] <= 16'b0000_0000_0000_0000;
array[17813] <= 16'b0000_0000_0000_0000;
array[17814] <= 16'b0000_0000_0000_0000;
array[17815] <= 16'b0000_0000_0000_0000;
array[17816] <= 16'b0000_0000_0000_0000;
array[17817] <= 16'b0000_0000_0000_0000;
array[17818] <= 16'b0000_0000_0000_0000;
array[17819] <= 16'b0000_0000_0000_0000;
array[17820] <= 16'b0000_0000_0000_0000;
array[17821] <= 16'b0000_0000_0000_0000;
array[17822] <= 16'b0000_0000_0000_0000;
array[17823] <= 16'b0000_0000_0000_0000;
array[17824] <= 16'b0000_0000_0000_0000;
array[17825] <= 16'b0000_0000_0000_0000;
array[17826] <= 16'b0000_0000_0000_0000;
array[17827] <= 16'b0000_0000_0000_0000;
array[17828] <= 16'b0000_0000_0000_0000;
array[17829] <= 16'b0000_0000_0000_0000;
array[17830] <= 16'b0000_0000_0000_0000;
array[17831] <= 16'b0000_0000_0000_0000;
array[17832] <= 16'b0000_0000_0000_0000;
array[17833] <= 16'b0000_0000_0000_0000;
array[17834] <= 16'b0000_0000_0000_0000;
array[17835] <= 16'b0000_0000_0000_0000;
array[17836] <= 16'b0000_0000_0000_0000;
array[17837] <= 16'b0000_0000_0000_0000;
array[17838] <= 16'b0000_0000_0000_0000;
array[17839] <= 16'b0000_0000_0000_0000;
array[17840] <= 16'b0000_0000_0000_0000;
array[17841] <= 16'b0000_0000_0000_0000;
array[17842] <= 16'b0000_0000_0000_0000;
array[17843] <= 16'b0000_0000_0000_0000;
array[17844] <= 16'b0000_0000_0000_0000;
array[17845] <= 16'b0000_0000_0000_0000;
array[17846] <= 16'b0000_0000_0000_0000;
array[17847] <= 16'b0000_0000_0000_0000;
array[17848] <= 16'b0000_0000_0000_0000;
array[17849] <= 16'b0000_0000_0000_0000;
array[17850] <= 16'b0000_0000_0000_0000;
array[17851] <= 16'b0000_0000_0000_0000;
array[17852] <= 16'b0000_0000_0000_0000;
array[17853] <= 16'b0000_0000_0000_0000;
array[17854] <= 16'b0000_0000_0000_0000;
array[17855] <= 16'b0000_0000_0000_0000;
array[17856] <= 16'b0000_0000_0000_0000;
array[17857] <= 16'b0000_0000_0000_0000;
array[17858] <= 16'b0000_0000_0000_0000;
array[17859] <= 16'b0000_0000_0000_0000;
array[17860] <= 16'b0000_0000_0000_0000;
array[17861] <= 16'b0000_0000_0000_0000;
array[17862] <= 16'b0000_0000_0000_0000;
array[17863] <= 16'b0000_0000_0000_0000;
array[17864] <= 16'b0000_0000_0000_0000;
array[17865] <= 16'b0000_0000_0000_0000;
array[17866] <= 16'b0000_0000_0000_0000;
array[17867] <= 16'b0000_0000_0000_0000;
array[17868] <= 16'b0000_0000_0000_0000;
array[17869] <= 16'b0000_0000_0000_0000;
array[17870] <= 16'b0000_0000_0000_0000;
array[17871] <= 16'b0000_0000_0000_0000;
array[17872] <= 16'b0000_0000_0000_0000;
array[17873] <= 16'b0000_0000_0000_0000;
array[17874] <= 16'b0000_0000_0000_0000;
array[17875] <= 16'b0000_0000_0000_0000;
array[17876] <= 16'b0000_0000_0000_0000;
array[17877] <= 16'b0000_0000_0000_0000;
array[17878] <= 16'b0000_0000_0000_0000;
array[17879] <= 16'b0000_0000_0000_0000;
array[17880] <= 16'b0000_0000_0000_0000;
array[17881] <= 16'b0000_0000_0000_0000;
array[17882] <= 16'b0000_0000_0000_0000;
array[17883] <= 16'b0000_0000_0000_0000;
array[17884] <= 16'b0000_0000_0000_0000;
array[17885] <= 16'b0000_0000_0000_0000;
array[17886] <= 16'b0000_0000_0000_0000;
array[17887] <= 16'b0000_0000_0000_0000;
array[17888] <= 16'b0000_0000_0000_0000;
array[17889] <= 16'b0000_0000_0000_0000;
array[17890] <= 16'b0000_0000_0000_0000;
array[17891] <= 16'b0000_0000_0000_0000;
array[17892] <= 16'b0000_0000_0000_0000;
array[17893] <= 16'b0000_0000_0000_0000;
array[17894] <= 16'b0000_0000_0000_0000;
array[17895] <= 16'b0000_0000_0000_0000;
array[17896] <= 16'b0000_0000_0000_0000;
array[17897] <= 16'b0000_0000_0000_0000;
array[17898] <= 16'b0000_0000_0000_0000;
array[17899] <= 16'b0000_0000_0000_0000;
array[17900] <= 16'b0000_0000_0000_0000;
array[17901] <= 16'b0000_0000_0000_0000;
array[17902] <= 16'b0000_0000_0000_0000;
array[17903] <= 16'b0000_0000_0000_0000;
array[17904] <= 16'b0000_0000_0000_0000;
array[17905] <= 16'b0000_0000_0000_0000;
array[17906] <= 16'b0000_0000_0000_0000;
array[17907] <= 16'b0000_0000_0000_0000;
array[17908] <= 16'b0000_0000_0000_0000;
array[17909] <= 16'b0000_0000_0000_0000;
array[17910] <= 16'b0000_0000_0000_0000;
array[17911] <= 16'b0000_0000_0000_0000;
array[17912] <= 16'b0000_0000_0000_0000;
array[17913] <= 16'b0000_0000_0000_0000;
array[17914] <= 16'b0000_0000_0000_0000;
array[17915] <= 16'b0000_0000_0000_0000;
array[17916] <= 16'b0000_0000_0000_0000;
array[17917] <= 16'b0000_0000_0000_0000;
array[17918] <= 16'b0000_0000_0000_0000;
array[17919] <= 16'b0000_0000_0000_0000;
array[17920] <= 16'b0000_0000_0000_0000;
array[17921] <= 16'b0000_0000_0000_0000;
array[17922] <= 16'b0000_0000_0000_0000;
array[17923] <= 16'b0000_0000_0000_0000;
array[17924] <= 16'b0000_0000_0000_0000;
array[17925] <= 16'b0000_0000_0000_0000;
array[17926] <= 16'b0000_0000_0000_0000;
array[17927] <= 16'b0000_0000_0000_0000;
array[17928] <= 16'b0000_0000_0000_0000;
array[17929] <= 16'b0000_0000_0000_0000;
array[17930] <= 16'b0000_0000_0000_0000;
array[17931] <= 16'b0000_0000_0000_0000;
array[17932] <= 16'b0000_0000_0000_0000;
array[17933] <= 16'b0000_0000_0000_0000;
array[17934] <= 16'b0000_0000_0000_0000;
array[17935] <= 16'b0000_0000_0000_0000;
array[17936] <= 16'b0000_0000_0000_0000;
array[17937] <= 16'b0000_0000_0000_0000;
array[17938] <= 16'b0000_0000_0000_0000;
array[17939] <= 16'b0000_0000_0000_0000;
array[17940] <= 16'b0000_0000_0000_0000;
array[17941] <= 16'b0000_0000_0000_0000;
array[17942] <= 16'b0000_0000_0000_0000;
array[17943] <= 16'b0000_0000_0000_0000;
array[17944] <= 16'b0000_0000_0000_0000;
array[17945] <= 16'b0000_0000_0000_0000;
array[17946] <= 16'b0000_0000_0000_0000;
array[17947] <= 16'b0000_0000_0000_0000;
array[17948] <= 16'b0000_0000_0000_0000;
array[17949] <= 16'b0000_0000_0000_0000;
array[17950] <= 16'b0000_0000_0000_0000;
array[17951] <= 16'b0000_0000_0000_0000;
array[17952] <= 16'b0000_0000_0000_0000;
array[17953] <= 16'b0000_0000_0000_0000;
array[17954] <= 16'b0000_0000_0000_0000;
array[17955] <= 16'b0000_0000_0000_0000;
array[17956] <= 16'b0000_0000_0000_0000;
array[17957] <= 16'b0000_0000_0000_0000;
array[17958] <= 16'b0000_0000_0000_0000;
array[17959] <= 16'b0000_0000_0000_0000;
array[17960] <= 16'b0000_0000_0000_0000;
array[17961] <= 16'b0000_0000_0000_0000;
array[17962] <= 16'b0000_0000_0000_0000;
array[17963] <= 16'b0000_0000_0000_0000;
array[17964] <= 16'b0000_0000_0000_0000;
array[17965] <= 16'b0000_0000_0000_0000;
array[17966] <= 16'b0000_0000_0000_0000;
array[17967] <= 16'b0000_0000_0000_0000;
array[17968] <= 16'b0000_0000_0000_0000;
array[17969] <= 16'b0000_0000_0000_0000;
array[17970] <= 16'b0000_0000_0000_0000;
array[17971] <= 16'b0000_0000_0000_0000;
array[17972] <= 16'b0000_0000_0000_0000;
array[17973] <= 16'b0000_0000_0000_0000;
array[17974] <= 16'b0000_0000_0000_0000;
array[17975] <= 16'b0000_0000_0000_0000;
array[17976] <= 16'b0000_0000_0000_0000;
array[17977] <= 16'b0000_0000_0000_0000;
array[17978] <= 16'b0000_0000_0000_0000;
array[17979] <= 16'b0000_0000_0000_0000;
array[17980] <= 16'b0000_0000_0000_0000;
array[17981] <= 16'b0000_0000_0000_0000;
array[17982] <= 16'b0000_0000_0000_0000;
array[17983] <= 16'b0000_0000_0000_0000;
array[17984] <= 16'b0000_0000_0000_0000;
array[17985] <= 16'b0000_0000_0000_0000;
array[17986] <= 16'b0000_0000_0000_0000;
array[17987] <= 16'b0000_0000_0000_0000;
array[17988] <= 16'b0000_0000_0000_0000;
array[17989] <= 16'b0000_0000_0000_0000;
array[17990] <= 16'b0000_0000_0000_0000;
array[17991] <= 16'b0000_0000_0000_0000;
array[17992] <= 16'b0000_0000_0000_0000;
array[17993] <= 16'b0000_0000_0000_0000;
array[17994] <= 16'b0000_0000_0000_0000;
array[17995] <= 16'b0000_0000_0000_0000;
array[17996] <= 16'b0000_0000_0000_0000;
array[17997] <= 16'b0000_0000_0000_0000;
array[17998] <= 16'b0000_0000_0000_0000;
array[17999] <= 16'b0000_0000_0000_0000;
array[18000] <= 16'b0000_0000_0000_0000;
array[18001] <= 16'b0000_0000_0000_0000;
array[18002] <= 16'b0000_0000_0000_0000;
array[18003] <= 16'b0000_0000_0000_0000;
array[18004] <= 16'b0000_0000_0000_0000;
array[18005] <= 16'b0000_0000_0000_0000;
array[18006] <= 16'b0000_0000_0000_0000;
array[18007] <= 16'b0000_0000_0000_0000;
array[18008] <= 16'b0000_0000_0000_0000;
array[18009] <= 16'b0000_0000_0000_0000;
array[18010] <= 16'b0000_0000_0000_0000;
array[18011] <= 16'b0000_0000_0000_0000;
array[18012] <= 16'b0000_0000_0000_0000;
array[18013] <= 16'b0000_0000_0000_0000;
array[18014] <= 16'b0000_0000_0000_0000;
array[18015] <= 16'b0000_0000_0000_0000;
array[18016] <= 16'b0000_0000_0000_0000;
array[18017] <= 16'b0000_0000_0000_0000;
array[18018] <= 16'b0000_0000_0000_0000;
array[18019] <= 16'b0000_0000_0000_0000;
array[18020] <= 16'b0000_0000_0000_0000;
array[18021] <= 16'b0000_0000_0000_0000;
array[18022] <= 16'b0000_0000_0000_0000;
array[18023] <= 16'b0000_0000_0000_0000;
array[18024] <= 16'b0000_0000_0000_0000;
array[18025] <= 16'b0000_0000_0000_0000;
array[18026] <= 16'b0000_0000_0000_0000;
array[18027] <= 16'b0000_0000_0000_0000;
array[18028] <= 16'b0000_0000_0000_0000;
array[18029] <= 16'b0000_0000_0000_0000;
array[18030] <= 16'b0000_0000_0000_0000;
array[18031] <= 16'b0000_0000_0000_0000;
array[18032] <= 16'b0000_0000_0000_0000;
array[18033] <= 16'b0000_0000_0000_0000;
array[18034] <= 16'b0000_0000_0000_0000;
array[18035] <= 16'b0000_0000_0000_0000;
array[18036] <= 16'b0000_0000_0000_0000;
array[18037] <= 16'b0000_0000_0000_0000;
array[18038] <= 16'b0000_0000_0000_0000;
array[18039] <= 16'b0000_0000_0000_0000;
array[18040] <= 16'b0000_0000_0000_0000;
array[18041] <= 16'b0000_0000_0000_0000;
array[18042] <= 16'b0000_0000_0000_0000;
array[18043] <= 16'b0000_0000_0000_0000;
array[18044] <= 16'b0000_0000_0000_0000;
array[18045] <= 16'b0000_0000_0000_0000;
array[18046] <= 16'b0000_0000_0000_0000;
array[18047] <= 16'b0000_0000_0000_0000;
array[18048] <= 16'b0000_0000_0000_0000;
array[18049] <= 16'b0000_0000_0000_0000;
array[18050] <= 16'b0000_0000_0000_0000;
array[18051] <= 16'b0000_0000_0000_0000;
array[18052] <= 16'b0000_0000_0000_0000;
array[18053] <= 16'b0000_0000_0000_0000;
array[18054] <= 16'b0000_0000_0000_0000;
array[18055] <= 16'b0000_0000_0000_0000;
array[18056] <= 16'b0000_0000_0000_0000;
array[18057] <= 16'b0000_0000_0000_0000;
array[18058] <= 16'b0000_0000_0000_0000;
array[18059] <= 16'b0000_0000_0000_0000;
array[18060] <= 16'b0000_0000_0000_0000;
array[18061] <= 16'b0000_0000_0000_0000;
array[18062] <= 16'b0000_0000_0000_0000;
array[18063] <= 16'b0000_0000_0000_0000;
array[18064] <= 16'b0000_0000_0000_0000;
array[18065] <= 16'b0000_0000_0000_0000;
array[18066] <= 16'b0000_0000_0000_0000;
array[18067] <= 16'b0000_0000_0000_0000;
array[18068] <= 16'b0000_0000_0000_0000;
array[18069] <= 16'b0000_0000_0000_0000;
array[18070] <= 16'b0000_0000_0000_0000;
array[18071] <= 16'b0000_0000_0000_0000;
array[18072] <= 16'b0000_0000_0000_0000;
array[18073] <= 16'b0000_0000_0000_0000;
array[18074] <= 16'b0000_0000_0000_0000;
array[18075] <= 16'b0000_0000_0000_0000;
array[18076] <= 16'b0000_0000_0000_0000;
array[18077] <= 16'b0000_0000_0000_0000;
array[18078] <= 16'b0000_0000_0000_0000;
array[18079] <= 16'b0000_0000_0000_0000;
array[18080] <= 16'b0000_0000_0000_0000;
array[18081] <= 16'b0000_0000_0000_0000;
array[18082] <= 16'b0000_0000_0000_0000;
array[18083] <= 16'b0000_0000_0000_0000;
array[18084] <= 16'b0000_0000_0000_0000;
array[18085] <= 16'b0000_0000_0000_0000;
array[18086] <= 16'b0000_0000_0000_0000;
array[18087] <= 16'b0000_0000_0000_0000;
array[18088] <= 16'b0000_0000_0000_0000;
array[18089] <= 16'b0000_0000_0000_0000;
array[18090] <= 16'b0000_0000_0000_0000;
array[18091] <= 16'b0000_0000_0000_0000;
array[18092] <= 16'b0000_0000_0000_0000;
array[18093] <= 16'b0000_0000_0000_0000;
array[18094] <= 16'b0000_0000_0000_0000;
array[18095] <= 16'b0000_0000_0000_0000;
array[18096] <= 16'b0000_0000_0000_0000;
array[18097] <= 16'b0000_0000_0000_0000;
array[18098] <= 16'b0000_0000_0000_0000;
array[18099] <= 16'b0000_0000_0000_0000;
array[18100] <= 16'b0000_0000_0000_0000;
array[18101] <= 16'b0000_0000_0000_0000;
array[18102] <= 16'b0000_0000_0000_0000;
array[18103] <= 16'b0000_0000_0000_0000;
array[18104] <= 16'b0000_0000_0000_0000;
array[18105] <= 16'b0000_0000_0000_0000;
array[18106] <= 16'b0000_0000_0000_0000;
array[18107] <= 16'b0000_0000_0000_0000;
array[18108] <= 16'b0000_0000_0000_0000;
array[18109] <= 16'b0000_0000_0000_0000;
array[18110] <= 16'b0000_0000_0000_0000;
array[18111] <= 16'b0000_0000_0000_0000;
array[18112] <= 16'b0000_0000_0000_0000;
array[18113] <= 16'b0000_0000_0000_0000;
array[18114] <= 16'b0000_0000_0000_0000;
array[18115] <= 16'b0000_0000_0000_0000;
array[18116] <= 16'b0000_0000_0000_0000;
array[18117] <= 16'b0000_0000_0000_0000;
array[18118] <= 16'b0000_0000_0000_0000;
array[18119] <= 16'b0000_0000_0000_0000;
array[18120] <= 16'b0000_0000_0000_0000;
array[18121] <= 16'b0000_0000_0000_0000;
array[18122] <= 16'b0000_0000_0000_0000;
array[18123] <= 16'b0000_0000_0000_0000;
array[18124] <= 16'b0000_0000_0000_0000;
array[18125] <= 16'b0000_0000_0000_0000;
array[18126] <= 16'b0000_0000_0000_0000;
array[18127] <= 16'b0000_0000_0000_0000;
array[18128] <= 16'b0000_0000_0000_0000;
array[18129] <= 16'b0000_0000_0000_0000;
array[18130] <= 16'b0000_0000_0000_0000;
array[18131] <= 16'b0000_0000_0000_0000;
array[18132] <= 16'b0000_0000_0000_0000;
array[18133] <= 16'b0000_0000_0000_0000;
array[18134] <= 16'b0000_0000_0000_0000;
array[18135] <= 16'b0000_0000_0000_0000;
array[18136] <= 16'b0000_0000_0000_0000;
array[18137] <= 16'b0000_0000_0000_0000;
array[18138] <= 16'b0000_0000_0000_0000;
array[18139] <= 16'b0000_0000_0000_0000;
array[18140] <= 16'b0000_0000_0000_0000;
array[18141] <= 16'b0000_0000_0000_0000;
array[18142] <= 16'b0000_0000_0000_0000;
array[18143] <= 16'b0000_0000_0000_0000;
array[18144] <= 16'b0000_0000_0000_0000;
array[18145] <= 16'b0000_0000_0000_0000;
array[18146] <= 16'b0000_0000_0000_0000;
array[18147] <= 16'b0000_0000_0000_0000;
array[18148] <= 16'b0000_0000_0000_0000;
array[18149] <= 16'b0000_0000_0000_0000;
array[18150] <= 16'b0000_0000_0000_0000;
array[18151] <= 16'b0000_0000_0000_0000;
array[18152] <= 16'b0000_0000_0000_0000;
array[18153] <= 16'b0000_0000_0000_0000;
array[18154] <= 16'b0000_0000_0000_0000;
array[18155] <= 16'b0000_0000_0000_0000;
array[18156] <= 16'b0000_0000_0000_0000;
array[18157] <= 16'b0000_0000_0000_0000;
array[18158] <= 16'b0000_0000_0000_0000;
array[18159] <= 16'b0000_0000_0000_0000;
array[18160] <= 16'b0000_0000_0000_0000;
array[18161] <= 16'b0000_0000_0000_0000;
array[18162] <= 16'b0000_0000_0000_0000;
array[18163] <= 16'b0000_0000_0000_0000;
array[18164] <= 16'b0000_0000_0000_0000;
array[18165] <= 16'b0000_0000_0000_0000;
array[18166] <= 16'b0000_0000_0000_0000;
array[18167] <= 16'b0000_0000_0000_0000;
array[18168] <= 16'b0000_0000_0000_0000;
array[18169] <= 16'b0000_0000_0000_0000;
array[18170] <= 16'b0000_0000_0000_0000;
array[18171] <= 16'b0000_0000_0000_0000;
array[18172] <= 16'b0000_0000_0000_0000;
array[18173] <= 16'b0000_0000_0000_0000;
array[18174] <= 16'b0000_0000_0000_0000;
array[18175] <= 16'b0000_0000_0000_0000;
array[18176] <= 16'b0000_0000_0000_0000;
array[18177] <= 16'b0000_0000_0000_0000;
array[18178] <= 16'b0000_0000_0000_0000;
array[18179] <= 16'b0000_0000_0000_0000;
array[18180] <= 16'b0000_0000_0000_0000;
array[18181] <= 16'b0000_0000_0000_0000;
array[18182] <= 16'b0000_0000_0000_0000;
array[18183] <= 16'b0000_0000_0000_0000;
array[18184] <= 16'b0000_0000_0000_0000;
array[18185] <= 16'b0000_0000_0000_0000;
array[18186] <= 16'b0000_0000_0000_0000;
array[18187] <= 16'b0000_0000_0000_0000;
array[18188] <= 16'b0000_0000_0000_0000;
array[18189] <= 16'b0000_0000_0000_0000;
array[18190] <= 16'b0000_0000_0000_0000;
array[18191] <= 16'b0000_0000_0000_0000;
array[18192] <= 16'b0000_0000_0000_0000;
array[18193] <= 16'b0000_0000_0000_0000;
array[18194] <= 16'b0000_0000_0000_0000;
array[18195] <= 16'b0000_0000_0000_0000;
array[18196] <= 16'b0000_0000_0000_0000;
array[18197] <= 16'b0000_0000_0000_0000;
array[18198] <= 16'b0000_0000_0000_0000;
array[18199] <= 16'b0000_0000_0000_0000;
array[18200] <= 16'b0000_0000_0000_0000;
array[18201] <= 16'b0000_0000_0000_0000;
array[18202] <= 16'b0000_0000_0000_0000;
array[18203] <= 16'b0000_0000_0000_0000;
array[18204] <= 16'b0000_0000_0000_0000;
array[18205] <= 16'b0000_0000_0000_0000;
array[18206] <= 16'b0000_0000_0000_0000;
array[18207] <= 16'b0000_0000_0000_0000;
array[18208] <= 16'b0000_0000_0000_0000;
array[18209] <= 16'b0000_0000_0000_0000;
array[18210] <= 16'b0000_0000_0000_0000;
array[18211] <= 16'b0000_0000_0000_0000;
array[18212] <= 16'b0000_0000_0000_0000;
array[18213] <= 16'b0000_0000_0000_0000;
array[18214] <= 16'b0000_0000_0000_0000;
array[18215] <= 16'b0000_0000_0000_0000;
array[18216] <= 16'b0000_0000_0000_0000;
array[18217] <= 16'b0000_0000_0000_0000;
array[18218] <= 16'b0000_0000_0000_0000;
array[18219] <= 16'b0000_0000_0000_0000;
array[18220] <= 16'b0000_0000_0000_0000;
array[18221] <= 16'b0000_0000_0000_0000;
array[18222] <= 16'b0000_0000_0000_0000;
array[18223] <= 16'b0000_0000_0000_0000;
array[18224] <= 16'b0000_0000_0000_0000;
array[18225] <= 16'b0000_0000_0000_0000;
array[18226] <= 16'b0000_0000_0000_0000;
array[18227] <= 16'b0000_0000_0000_0000;
array[18228] <= 16'b0000_0000_0000_0000;
array[18229] <= 16'b0000_0000_0000_0000;
array[18230] <= 16'b0000_0000_0000_0000;
array[18231] <= 16'b0000_0000_0000_0000;
array[18232] <= 16'b0000_0000_0000_0000;
array[18233] <= 16'b0000_0000_0000_0000;
array[18234] <= 16'b0000_0000_0000_0000;
array[18235] <= 16'b0000_0000_0000_0000;
array[18236] <= 16'b0000_0000_0000_0000;
array[18237] <= 16'b0000_0000_0000_0000;
array[18238] <= 16'b0000_0000_0000_0000;
array[18239] <= 16'b0000_0000_0000_0000;
array[18240] <= 16'b0000_0000_0000_0000;
array[18241] <= 16'b0000_0000_0000_0000;
array[18242] <= 16'b0000_0000_0000_0000;
array[18243] <= 16'b0000_0000_0000_0000;
array[18244] <= 16'b0000_0000_0000_0000;
array[18245] <= 16'b0000_0000_0000_0000;
array[18246] <= 16'b0000_0000_0000_0000;
array[18247] <= 16'b0000_0000_0000_0000;
array[18248] <= 16'b0000_0000_0000_0000;
array[18249] <= 16'b0000_0000_0000_0000;
array[18250] <= 16'b0000_0000_0000_0000;
array[18251] <= 16'b0000_0000_0000_0000;
array[18252] <= 16'b0000_0000_0000_0000;
array[18253] <= 16'b0000_0000_0000_0000;
array[18254] <= 16'b0000_0000_0000_0000;
array[18255] <= 16'b0000_0000_0000_0000;
array[18256] <= 16'b0000_0000_0000_0000;
array[18257] <= 16'b0000_0000_0000_0000;
array[18258] <= 16'b0000_0000_0000_0000;
array[18259] <= 16'b0000_0000_0000_0000;
array[18260] <= 16'b0000_0000_0000_0000;
array[18261] <= 16'b0000_0000_0000_0000;
array[18262] <= 16'b0000_0000_0000_0000;
array[18263] <= 16'b0000_0000_0000_0000;
array[18264] <= 16'b0000_0000_0000_0000;
array[18265] <= 16'b0000_0000_0000_0000;
array[18266] <= 16'b0000_0000_0000_0000;
array[18267] <= 16'b0000_0000_0000_0000;
array[18268] <= 16'b0000_0000_0000_0000;
array[18269] <= 16'b0000_0000_0000_0000;
array[18270] <= 16'b0000_0000_0000_0000;
array[18271] <= 16'b0000_0000_0000_0000;
array[18272] <= 16'b0000_0000_0000_0000;
array[18273] <= 16'b0000_0000_0000_0000;
array[18274] <= 16'b0000_0000_0000_0000;
array[18275] <= 16'b0000_0000_0000_0000;
array[18276] <= 16'b0000_0000_0000_0000;
array[18277] <= 16'b0000_0000_0000_0000;
array[18278] <= 16'b0000_0000_0000_0000;
array[18279] <= 16'b0000_0000_0000_0000;
array[18280] <= 16'b0000_0000_0000_0000;
array[18281] <= 16'b0000_0000_0000_0000;
array[18282] <= 16'b0000_0000_0000_0000;
array[18283] <= 16'b0000_0000_0000_0000;
array[18284] <= 16'b0000_0000_0000_0000;
array[18285] <= 16'b0000_0000_0000_0000;
array[18286] <= 16'b0000_0000_0000_0000;
array[18287] <= 16'b0000_0000_0000_0000;
array[18288] <= 16'b0000_0000_0000_0000;
array[18289] <= 16'b0000_0000_0000_0000;
array[18290] <= 16'b0000_0000_0000_0000;
array[18291] <= 16'b0000_0000_0000_0000;
array[18292] <= 16'b0000_0000_0000_0000;
array[18293] <= 16'b0000_0000_0000_0000;
array[18294] <= 16'b0000_0000_0000_0000;
array[18295] <= 16'b0000_0000_0000_0000;
array[18296] <= 16'b0000_0000_0000_0000;
array[18297] <= 16'b0000_0000_0000_0000;
array[18298] <= 16'b0000_0000_0000_0000;
array[18299] <= 16'b0000_0000_0000_0000;
array[18300] <= 16'b0000_0000_0000_0000;
array[18301] <= 16'b0000_0000_0000_0000;
array[18302] <= 16'b0000_0000_0000_0000;
array[18303] <= 16'b0000_0000_0000_0000;
array[18304] <= 16'b0000_0000_0000_0000;
array[18305] <= 16'b0000_0000_0000_0000;
array[18306] <= 16'b0000_0000_0000_0000;
array[18307] <= 16'b0000_0000_0000_0000;
array[18308] <= 16'b0000_0000_0000_0000;
array[18309] <= 16'b0000_0000_0000_0000;
array[18310] <= 16'b0000_0000_0000_0000;
array[18311] <= 16'b0000_0000_0000_0000;
array[18312] <= 16'b0000_0000_0000_0000;
array[18313] <= 16'b0000_0000_0000_0000;
array[18314] <= 16'b0000_0000_0000_0000;
array[18315] <= 16'b0000_0000_0000_0000;
array[18316] <= 16'b0000_0000_0000_0000;
array[18317] <= 16'b0000_0000_0000_0000;
array[18318] <= 16'b0000_0000_0000_0000;
array[18319] <= 16'b0000_0000_0000_0000;
array[18320] <= 16'b0000_0000_0000_0000;
array[18321] <= 16'b0000_0000_0000_0000;
array[18322] <= 16'b0000_0000_0000_0000;
array[18323] <= 16'b0000_0000_0000_0000;
array[18324] <= 16'b0000_0000_0000_0000;
array[18325] <= 16'b0000_0000_0000_0000;
array[18326] <= 16'b0000_0000_0000_0000;
array[18327] <= 16'b0000_0000_0000_0000;
array[18328] <= 16'b0000_0000_0000_0000;
array[18329] <= 16'b0000_0000_0000_0000;
array[18330] <= 16'b0000_0000_0000_0000;
array[18331] <= 16'b0000_0000_0000_0000;
array[18332] <= 16'b0000_0000_0000_0000;
array[18333] <= 16'b0000_0000_0000_0000;
array[18334] <= 16'b0000_0000_0000_0000;
array[18335] <= 16'b0000_0000_0000_0000;
array[18336] <= 16'b0000_0000_0000_0000;
array[18337] <= 16'b0000_0000_0000_0000;
array[18338] <= 16'b0000_0000_0000_0000;
array[18339] <= 16'b0000_0000_0000_0000;
array[18340] <= 16'b0000_0000_0000_0000;
array[18341] <= 16'b0000_0000_0000_0000;
array[18342] <= 16'b0000_0000_0000_0000;
array[18343] <= 16'b0000_0000_0000_0000;
array[18344] <= 16'b0000_0000_0000_0000;
array[18345] <= 16'b0000_0000_0000_0000;
array[18346] <= 16'b0000_0000_0000_0000;
array[18347] <= 16'b0000_0000_0000_0000;
array[18348] <= 16'b0000_0000_0000_0000;
array[18349] <= 16'b0000_0000_0000_0000;
array[18350] <= 16'b0000_0000_0000_0000;
array[18351] <= 16'b0000_0000_0000_0000;
array[18352] <= 16'b0000_0000_0000_0000;
array[18353] <= 16'b0000_0000_0000_0000;
array[18354] <= 16'b0000_0000_0000_0000;
array[18355] <= 16'b0000_0000_0000_0000;
array[18356] <= 16'b0000_0000_0000_0000;
array[18357] <= 16'b0000_0000_0000_0000;
array[18358] <= 16'b0000_0000_0000_0000;
array[18359] <= 16'b0000_0000_0000_0000;
array[18360] <= 16'b0000_0000_0000_0000;
array[18361] <= 16'b0000_0000_0000_0000;
array[18362] <= 16'b0000_0000_0000_0000;
array[18363] <= 16'b0000_0000_0000_0000;
array[18364] <= 16'b0000_0000_0000_0000;
array[18365] <= 16'b0000_0000_0000_0000;
array[18366] <= 16'b0000_0000_0000_0000;
array[18367] <= 16'b0000_0000_0000_0000;
array[18368] <= 16'b0000_0000_0000_0000;
array[18369] <= 16'b0000_0000_0000_0000;
array[18370] <= 16'b0000_0000_0000_0000;
array[18371] <= 16'b0000_0000_0000_0000;
array[18372] <= 16'b0000_0000_0000_0000;
array[18373] <= 16'b0000_0000_0000_0000;
array[18374] <= 16'b0000_0000_0000_0000;
array[18375] <= 16'b0000_0000_0000_0000;
array[18376] <= 16'b0000_0000_0000_0000;
array[18377] <= 16'b0000_0000_0000_0000;
array[18378] <= 16'b0000_0000_0000_0000;
array[18379] <= 16'b0000_0000_0000_0000;
array[18380] <= 16'b0000_0000_0000_0000;
array[18381] <= 16'b0000_0000_0000_0000;
array[18382] <= 16'b0000_0000_0000_0000;
array[18383] <= 16'b0000_0000_0000_0000;
array[18384] <= 16'b0000_0000_0000_0000;
array[18385] <= 16'b0000_0000_0000_0000;
array[18386] <= 16'b0000_0000_0000_0000;
array[18387] <= 16'b0000_0000_0000_0000;
array[18388] <= 16'b0000_0000_0000_0000;
array[18389] <= 16'b0000_0000_0000_0000;
array[18390] <= 16'b0000_0000_0000_0000;
array[18391] <= 16'b0000_0000_0000_0000;
array[18392] <= 16'b0000_0000_0000_0000;
array[18393] <= 16'b0000_0000_0000_0000;
array[18394] <= 16'b0000_0000_0000_0000;
array[18395] <= 16'b0000_0000_0000_0000;
array[18396] <= 16'b0000_0000_0000_0000;
array[18397] <= 16'b0000_0000_0000_0000;
array[18398] <= 16'b0000_0000_0000_0000;
array[18399] <= 16'b0000_0000_0000_0000;
array[18400] <= 16'b0000_0000_0000_0000;
array[18401] <= 16'b0000_0000_0000_0000;
array[18402] <= 16'b0000_0000_0000_0000;
array[18403] <= 16'b0000_0000_0000_0000;
array[18404] <= 16'b0000_0000_0000_0000;
array[18405] <= 16'b0000_0000_0000_0000;
array[18406] <= 16'b0000_0000_0000_0000;
array[18407] <= 16'b0000_0000_0000_0000;
array[18408] <= 16'b0000_0000_0000_0000;
array[18409] <= 16'b0000_0000_0000_0000;
array[18410] <= 16'b0000_0000_0000_0000;
array[18411] <= 16'b0000_0000_0000_0000;
array[18412] <= 16'b0000_0000_0000_0000;
array[18413] <= 16'b0000_0000_0000_0000;
array[18414] <= 16'b0000_0000_0000_0000;
array[18415] <= 16'b0000_0000_0000_0000;
array[18416] <= 16'b0000_0000_0000_0000;
array[18417] <= 16'b0000_0000_0000_0000;
array[18418] <= 16'b0000_0000_0000_0000;
array[18419] <= 16'b0000_0000_0000_0000;
array[18420] <= 16'b0000_0000_0000_0000;
array[18421] <= 16'b0000_0000_0000_0000;
array[18422] <= 16'b0000_0000_0000_0000;
array[18423] <= 16'b0000_0000_0000_0000;
array[18424] <= 16'b0000_0000_0000_0000;
array[18425] <= 16'b0000_0000_0000_0000;
array[18426] <= 16'b0000_0000_0000_0000;
array[18427] <= 16'b0000_0000_0000_0000;
array[18428] <= 16'b0000_0000_0000_0000;
array[18429] <= 16'b0000_0000_0000_0000;
array[18430] <= 16'b0000_0000_0000_0000;
array[18431] <= 16'b0000_0000_0000_0000;
array[18432] <= 16'b0000_0000_0000_0000;
array[18433] <= 16'b0000_0000_0000_0000;
array[18434] <= 16'b0000_0000_0000_0000;
array[18435] <= 16'b0000_0000_0000_0000;
array[18436] <= 16'b0000_0000_0000_0000;
array[18437] <= 16'b0000_0000_0000_0000;
array[18438] <= 16'b0000_0000_0000_0000;
array[18439] <= 16'b0000_0000_0000_0000;
array[18440] <= 16'b0000_0000_0000_0000;
array[18441] <= 16'b0000_0000_0000_0000;
array[18442] <= 16'b0000_0000_0000_0000;
array[18443] <= 16'b0000_0000_0000_0000;
array[18444] <= 16'b0000_0000_0000_0000;
array[18445] <= 16'b0000_0000_0000_0000;
array[18446] <= 16'b0000_0000_0000_0000;
array[18447] <= 16'b0000_0000_0000_0000;
array[18448] <= 16'b0000_0000_0000_0000;
array[18449] <= 16'b0000_0000_0000_0000;
array[18450] <= 16'b0000_0000_0000_0000;
array[18451] <= 16'b0000_0000_0000_0000;
array[18452] <= 16'b0000_0000_0000_0000;
array[18453] <= 16'b0000_0000_0000_0000;
array[18454] <= 16'b0000_0000_0000_0000;
array[18455] <= 16'b0000_0000_0000_0000;
array[18456] <= 16'b0000_0000_0000_0000;
array[18457] <= 16'b0000_0000_0000_0000;
array[18458] <= 16'b0000_0000_0000_0000;
array[18459] <= 16'b0000_0000_0000_0000;
array[18460] <= 16'b0000_0000_0000_0000;
array[18461] <= 16'b0000_0000_0000_0000;
array[18462] <= 16'b0000_0000_0000_0000;
array[18463] <= 16'b0000_0000_0000_0000;
array[18464] <= 16'b0000_0000_0000_0000;
array[18465] <= 16'b0000_0000_0000_0000;
array[18466] <= 16'b0000_0000_0000_0000;
array[18467] <= 16'b0000_0000_0000_0000;
array[18468] <= 16'b0000_0000_0000_0000;
array[18469] <= 16'b0000_0000_0000_0000;
array[18470] <= 16'b0000_0000_0000_0000;
array[18471] <= 16'b0000_0000_0000_0000;
array[18472] <= 16'b0000_0000_0000_0000;
array[18473] <= 16'b0000_0000_0000_0000;
array[18474] <= 16'b0000_0000_0000_0000;
array[18475] <= 16'b0000_0000_0000_0000;
array[18476] <= 16'b0000_0000_0000_0000;
array[18477] <= 16'b0000_0000_0000_0000;
array[18478] <= 16'b0000_0000_0000_0000;
array[18479] <= 16'b0000_0000_0000_0000;
array[18480] <= 16'b0000_0000_0000_0000;
array[18481] <= 16'b0000_0000_0000_0000;
array[18482] <= 16'b0000_0000_0000_0000;
array[18483] <= 16'b0000_0000_0000_0000;
array[18484] <= 16'b0000_0000_0000_0000;
array[18485] <= 16'b0000_0000_0000_0000;
array[18486] <= 16'b0000_0000_0000_0000;
array[18487] <= 16'b0000_0000_0000_0000;
array[18488] <= 16'b0000_0000_0000_0000;
array[18489] <= 16'b0000_0000_0000_0000;
array[18490] <= 16'b0000_0000_0000_0000;
array[18491] <= 16'b0000_0000_0000_0000;
array[18492] <= 16'b0000_0000_0000_0000;
array[18493] <= 16'b0000_0000_0000_0000;
array[18494] <= 16'b0000_0000_0000_0000;
array[18495] <= 16'b0000_0000_0000_0000;
array[18496] <= 16'b0000_0000_0000_0000;
array[18497] <= 16'b0000_0000_0000_0000;
array[18498] <= 16'b0000_0000_0000_0000;
array[18499] <= 16'b0000_0000_0000_0000;
array[18500] <= 16'b0000_0000_0000_0000;
array[18501] <= 16'b0000_0000_0000_0000;
array[18502] <= 16'b0000_0000_0000_0000;
array[18503] <= 16'b0000_0000_0000_0000;
array[18504] <= 16'b0000_0000_0000_0000;
array[18505] <= 16'b0000_0000_0000_0000;
array[18506] <= 16'b0000_0000_0000_0000;
array[18507] <= 16'b0000_0000_0000_0000;
array[18508] <= 16'b0000_0000_0000_0000;
array[18509] <= 16'b0000_0000_0000_0000;
array[18510] <= 16'b0000_0000_0000_0000;
array[18511] <= 16'b0000_0000_0000_0000;
array[18512] <= 16'b0000_0000_0000_0000;
array[18513] <= 16'b0000_0000_0000_0000;
array[18514] <= 16'b0000_0000_0000_0000;
array[18515] <= 16'b0000_0000_0000_0000;
array[18516] <= 16'b0000_0000_0000_0000;
array[18517] <= 16'b0000_0000_0000_0000;
array[18518] <= 16'b0000_0000_0000_0000;
array[18519] <= 16'b0000_0000_0000_0000;
array[18520] <= 16'b0000_0000_0000_0000;
array[18521] <= 16'b0000_0000_0000_0000;
array[18522] <= 16'b0000_0000_0000_0000;
array[18523] <= 16'b0000_0000_0000_0000;
array[18524] <= 16'b0000_0000_0000_0000;
array[18525] <= 16'b0000_0000_0000_0000;
array[18526] <= 16'b0000_0000_0000_0000;
array[18527] <= 16'b0000_0000_0000_0000;
array[18528] <= 16'b0000_0000_0000_0000;
array[18529] <= 16'b0000_0000_0000_0000;
array[18530] <= 16'b0000_0000_0000_0000;
array[18531] <= 16'b0000_0000_0000_0000;
array[18532] <= 16'b0000_0000_0000_0000;
array[18533] <= 16'b0000_0000_0000_0000;
array[18534] <= 16'b0000_0000_0000_0000;
array[18535] <= 16'b0000_0000_0000_0000;
array[18536] <= 16'b0000_0000_0000_0000;
array[18537] <= 16'b0000_0000_0000_0000;
array[18538] <= 16'b0000_0000_0000_0000;
array[18539] <= 16'b0000_0000_0000_0000;
array[18540] <= 16'b0000_0000_0000_0000;
array[18541] <= 16'b0000_0000_0000_0000;
array[18542] <= 16'b0000_0000_0000_0000;
array[18543] <= 16'b0000_0000_0000_0000;
array[18544] <= 16'b0000_0000_0000_0000;
array[18545] <= 16'b0000_0000_0000_0000;
array[18546] <= 16'b0000_0000_0000_0000;
array[18547] <= 16'b0000_0000_0000_0000;
array[18548] <= 16'b0000_0000_0000_0000;
array[18549] <= 16'b0000_0000_0000_0000;
array[18550] <= 16'b0000_0000_0000_0000;
array[18551] <= 16'b0000_0000_0000_0000;
array[18552] <= 16'b0000_0000_0000_0000;
array[18553] <= 16'b0000_0000_0000_0000;
array[18554] <= 16'b0000_0000_0000_0000;
array[18555] <= 16'b0000_0000_0000_0000;
array[18556] <= 16'b0000_0000_0000_0000;
array[18557] <= 16'b0000_0000_0000_0000;
array[18558] <= 16'b0000_0000_0000_0000;
array[18559] <= 16'b0000_0000_0000_0000;
array[18560] <= 16'b0000_0000_0000_0000;
array[18561] <= 16'b0000_0000_0000_0000;
array[18562] <= 16'b0000_0000_0000_0000;
array[18563] <= 16'b0000_0000_0000_0000;
array[18564] <= 16'b0000_0000_0000_0000;
array[18565] <= 16'b0000_0000_0000_0000;
array[18566] <= 16'b0000_0000_0000_0000;
array[18567] <= 16'b0000_0000_0000_0000;
array[18568] <= 16'b0000_0000_0000_0000;
array[18569] <= 16'b0000_0000_0000_0000;
array[18570] <= 16'b0000_0000_0000_0000;
array[18571] <= 16'b0000_0000_0000_0000;
array[18572] <= 16'b0000_0000_0000_0000;
array[18573] <= 16'b0000_0000_0000_0000;
array[18574] <= 16'b0000_0000_0000_0000;
array[18575] <= 16'b0000_0000_0000_0000;
array[18576] <= 16'b0000_0000_0000_0000;
array[18577] <= 16'b0000_0000_0000_0000;
array[18578] <= 16'b0000_0000_0000_0000;
array[18579] <= 16'b0000_0000_0000_0000;
array[18580] <= 16'b0000_0000_0000_0000;
array[18581] <= 16'b0000_0000_0000_0000;
array[18582] <= 16'b0000_0000_0000_0000;
array[18583] <= 16'b0000_0000_0000_0000;
array[18584] <= 16'b0000_0000_0000_0000;
array[18585] <= 16'b0000_0000_0000_0000;
array[18586] <= 16'b0000_0000_0000_0000;
array[18587] <= 16'b0000_0000_0000_0000;
array[18588] <= 16'b0000_0000_0000_0000;
array[18589] <= 16'b0000_0000_0000_0000;
array[18590] <= 16'b0000_0000_0000_0000;
array[18591] <= 16'b0000_0000_0000_0000;
array[18592] <= 16'b0000_0000_0000_0000;
array[18593] <= 16'b0000_0000_0000_0000;
array[18594] <= 16'b0000_0000_0000_0000;
array[18595] <= 16'b0000_0000_0000_0000;
array[18596] <= 16'b0000_0000_0000_0000;
array[18597] <= 16'b0000_0000_0000_0000;
array[18598] <= 16'b0000_0000_0000_0000;
array[18599] <= 16'b0000_0000_0000_0000;
array[18600] <= 16'b0000_0000_0000_0000;
array[18601] <= 16'b0000_0000_0000_0000;
array[18602] <= 16'b0000_0000_0000_0000;
array[18603] <= 16'b0000_0000_0000_0000;
array[18604] <= 16'b0000_0000_0000_0000;
array[18605] <= 16'b0000_0000_0000_0000;
array[18606] <= 16'b0000_0000_0000_0000;
array[18607] <= 16'b0000_0000_0000_0000;
array[18608] <= 16'b0000_0000_0000_0000;
array[18609] <= 16'b0000_0000_0000_0000;
array[18610] <= 16'b0000_0000_0000_0000;
array[18611] <= 16'b0000_0000_0000_0000;
array[18612] <= 16'b0000_0000_0000_0000;
array[18613] <= 16'b0000_0000_0000_0000;
array[18614] <= 16'b0000_0000_0000_0000;
array[18615] <= 16'b0000_0000_0000_0000;
array[18616] <= 16'b0000_0000_0000_0000;
array[18617] <= 16'b0000_0000_0000_0000;
array[18618] <= 16'b0000_0000_0000_0000;
array[18619] <= 16'b0000_0000_0000_0000;
array[18620] <= 16'b0000_0000_0000_0000;
array[18621] <= 16'b0000_0000_0000_0000;
array[18622] <= 16'b0000_0000_0000_0000;
array[18623] <= 16'b0000_0000_0000_0000;
array[18624] <= 16'b0000_0000_0000_0000;
array[18625] <= 16'b0000_0000_0000_0000;
array[18626] <= 16'b0000_0000_0000_0000;
array[18627] <= 16'b0000_0000_0000_0000;
array[18628] <= 16'b0000_0000_0000_0000;
array[18629] <= 16'b0000_0000_0000_0000;
array[18630] <= 16'b0000_0000_0000_0000;
array[18631] <= 16'b0000_0000_0000_0000;
array[18632] <= 16'b0000_0000_0000_0000;
array[18633] <= 16'b0000_0000_0000_0000;
array[18634] <= 16'b0000_0000_0000_0000;
array[18635] <= 16'b0000_0000_0000_0000;
array[18636] <= 16'b0000_0000_0000_0000;
array[18637] <= 16'b0000_0000_0000_0000;
array[18638] <= 16'b0000_0000_0000_0000;
array[18639] <= 16'b0000_0000_0000_0000;
array[18640] <= 16'b0000_0000_0000_0000;
array[18641] <= 16'b0000_0000_0000_0000;
array[18642] <= 16'b0000_0000_0000_0000;
array[18643] <= 16'b0000_0000_0000_0000;
array[18644] <= 16'b0000_0000_0000_0000;
array[18645] <= 16'b0000_0000_0000_0000;
array[18646] <= 16'b0000_0000_0000_0000;
array[18647] <= 16'b0000_0000_0000_0000;
array[18648] <= 16'b0000_0000_0000_0000;
array[18649] <= 16'b0000_0000_0000_0000;
array[18650] <= 16'b0000_0000_0000_0000;
array[18651] <= 16'b0000_0000_0000_0000;
array[18652] <= 16'b0000_0000_0000_0000;
array[18653] <= 16'b0000_0000_0000_0000;
array[18654] <= 16'b0000_0000_0000_0000;
array[18655] <= 16'b0000_0000_0000_0000;
array[18656] <= 16'b0000_0000_0000_0000;
array[18657] <= 16'b0000_0000_0000_0000;
array[18658] <= 16'b0000_0000_0000_0000;
array[18659] <= 16'b0000_0000_0000_0000;
array[18660] <= 16'b0000_0000_0000_0000;
array[18661] <= 16'b0000_0000_0000_0000;
array[18662] <= 16'b0000_0000_0000_0000;
array[18663] <= 16'b0000_0000_0000_0000;
array[18664] <= 16'b0000_0000_0000_0000;
array[18665] <= 16'b0000_0000_0000_0000;
array[18666] <= 16'b0000_0000_0000_0000;
array[18667] <= 16'b0000_0000_0000_0000;
array[18668] <= 16'b0000_0000_0000_0000;
array[18669] <= 16'b0000_0000_0000_0000;
array[18670] <= 16'b0000_0000_0000_0000;
array[18671] <= 16'b0000_0000_0000_0000;
array[18672] <= 16'b0000_0000_0000_0000;
array[18673] <= 16'b0000_0000_0000_0000;
array[18674] <= 16'b0000_0000_0000_0000;
array[18675] <= 16'b0000_0000_0000_0000;
array[18676] <= 16'b0000_0000_0000_0000;
array[18677] <= 16'b0000_0000_0000_0000;
array[18678] <= 16'b0000_0000_0000_0000;
array[18679] <= 16'b0000_0000_0000_0000;
array[18680] <= 16'b0000_0000_0000_0000;
array[18681] <= 16'b0000_0000_0000_0000;
array[18682] <= 16'b0000_0000_0000_0000;
array[18683] <= 16'b0000_0000_0000_0000;
array[18684] <= 16'b0000_0000_0000_0000;
array[18685] <= 16'b0000_0000_0000_0000;
array[18686] <= 16'b0000_0000_0000_0000;
array[18687] <= 16'b0000_0000_0000_0000;
array[18688] <= 16'b0000_0000_0000_0000;
array[18689] <= 16'b0000_0000_0000_0000;
array[18690] <= 16'b0000_0000_0000_0000;
array[18691] <= 16'b0000_0000_0000_0000;
array[18692] <= 16'b0000_0000_0000_0000;
array[18693] <= 16'b0000_0000_0000_0000;
array[18694] <= 16'b0000_0000_0000_0000;
array[18695] <= 16'b0000_0000_0000_0000;
array[18696] <= 16'b0000_0000_0000_0000;
array[18697] <= 16'b0000_0000_0000_0000;
array[18698] <= 16'b0000_0000_0000_0000;
array[18699] <= 16'b0000_0000_0000_0000;
array[18700] <= 16'b0000_0000_0000_0000;
array[18701] <= 16'b0000_0000_0000_0000;
array[18702] <= 16'b0000_0000_0000_0000;
array[18703] <= 16'b0000_0000_0000_0000;
array[18704] <= 16'b0000_0000_0000_0000;
array[18705] <= 16'b0000_0000_0000_0000;
array[18706] <= 16'b0000_0000_0000_0000;
array[18707] <= 16'b0000_0000_0000_0000;
array[18708] <= 16'b0000_0000_0000_0000;
array[18709] <= 16'b0000_0000_0000_0000;
array[18710] <= 16'b0000_0000_0000_0000;
array[18711] <= 16'b0000_0000_0000_0000;
array[18712] <= 16'b0000_0000_0000_0000;
array[18713] <= 16'b0000_0000_0000_0000;
array[18714] <= 16'b0000_0000_0000_0000;
array[18715] <= 16'b0000_0000_0000_0000;
array[18716] <= 16'b0000_0000_0000_0000;
array[18717] <= 16'b0000_0000_0000_0000;
array[18718] <= 16'b0000_0000_0000_0000;
array[18719] <= 16'b0000_0000_0000_0000;
array[18720] <= 16'b0000_0000_0000_0000;
array[18721] <= 16'b0000_0000_0000_0000;
array[18722] <= 16'b0000_0000_0000_0000;
array[18723] <= 16'b0000_0000_0000_0000;
array[18724] <= 16'b0000_0000_0000_0000;
array[18725] <= 16'b0000_0000_0000_0000;
array[18726] <= 16'b0000_0000_0000_0000;
array[18727] <= 16'b0000_0000_0000_0000;
array[18728] <= 16'b0000_0000_0000_0000;
array[18729] <= 16'b0000_0000_0000_0000;
array[18730] <= 16'b0000_0000_0000_0000;
array[18731] <= 16'b0000_0000_0000_0000;
array[18732] <= 16'b0000_0000_0000_0000;
array[18733] <= 16'b0000_0000_0000_0000;
array[18734] <= 16'b0000_0000_0000_0000;
array[18735] <= 16'b0000_0000_0000_0000;
array[18736] <= 16'b0000_0000_0000_0000;
array[18737] <= 16'b0000_0000_0000_0000;
array[18738] <= 16'b0000_0000_0000_0000;
array[18739] <= 16'b0000_0000_0000_0000;
array[18740] <= 16'b0000_0000_0000_0000;
array[18741] <= 16'b0000_0000_0000_0000;
array[18742] <= 16'b0000_0000_0000_0000;
array[18743] <= 16'b0000_0000_0000_0000;
array[18744] <= 16'b0000_0000_0000_0000;
array[18745] <= 16'b0000_0000_0000_0000;
array[18746] <= 16'b0000_0000_0000_0000;
array[18747] <= 16'b0000_0000_0000_0000;
array[18748] <= 16'b0000_0000_0000_0000;
array[18749] <= 16'b0000_0000_0000_0000;
array[18750] <= 16'b0000_0000_0000_0000;
array[18751] <= 16'b0000_0000_0000_0000;
array[18752] <= 16'b0000_0000_0000_0000;
array[18753] <= 16'b0000_0000_0000_0000;
array[18754] <= 16'b0000_0000_0000_0000;
array[18755] <= 16'b0000_0000_0000_0000;
array[18756] <= 16'b0000_0000_0000_0000;
array[18757] <= 16'b0000_0000_0000_0000;
array[18758] <= 16'b0000_0000_0000_0000;
array[18759] <= 16'b0000_0000_0000_0000;
array[18760] <= 16'b0000_0000_0000_0000;
array[18761] <= 16'b0000_0000_0000_0000;
array[18762] <= 16'b0000_0000_0000_0000;
array[18763] <= 16'b0000_0000_0000_0000;
array[18764] <= 16'b0000_0000_0000_0000;
array[18765] <= 16'b0000_0000_0000_0000;
array[18766] <= 16'b0000_0000_0000_0000;
array[18767] <= 16'b0000_0000_0000_0000;
array[18768] <= 16'b0000_0000_0000_0000;
array[18769] <= 16'b0000_0000_0000_0000;
array[18770] <= 16'b0000_0000_0000_0000;
array[18771] <= 16'b0000_0000_0000_0000;
array[18772] <= 16'b0000_0000_0000_0000;
array[18773] <= 16'b0000_0000_0000_0000;
array[18774] <= 16'b0000_0000_0000_0000;
array[18775] <= 16'b0000_0000_0000_0000;
array[18776] <= 16'b0000_0000_0000_0000;
array[18777] <= 16'b0000_0000_0000_0000;
array[18778] <= 16'b0000_0000_0000_0000;
array[18779] <= 16'b0000_0000_0000_0000;
array[18780] <= 16'b0000_0000_0000_0000;
array[18781] <= 16'b0000_0000_0000_0000;
array[18782] <= 16'b0000_0000_0000_0000;
array[18783] <= 16'b0000_0000_0000_0000;
array[18784] <= 16'b0000_0000_0000_0000;
array[18785] <= 16'b0000_0000_0000_0000;
array[18786] <= 16'b0000_0000_0000_0000;
array[18787] <= 16'b0000_0000_0000_0000;
array[18788] <= 16'b0000_0000_0000_0000;
array[18789] <= 16'b0000_0000_0000_0000;
array[18790] <= 16'b0000_0000_0000_0000;
array[18791] <= 16'b0000_0000_0000_0000;
array[18792] <= 16'b0000_0000_0000_0000;
array[18793] <= 16'b0000_0000_0000_0000;
array[18794] <= 16'b0000_0000_0000_0000;
array[18795] <= 16'b0000_0000_0000_0000;
array[18796] <= 16'b0000_0000_0000_0000;
array[18797] <= 16'b0000_0000_0000_0000;
array[18798] <= 16'b0000_0000_0000_0000;
array[18799] <= 16'b0000_0000_0000_0000;
array[18800] <= 16'b0000_0000_0000_0000;
array[18801] <= 16'b0000_0000_0000_0000;
array[18802] <= 16'b0000_0000_0000_0000;
array[18803] <= 16'b0000_0000_0000_0000;
array[18804] <= 16'b0000_0000_0000_0000;
array[18805] <= 16'b0000_0000_0000_0000;
array[18806] <= 16'b0000_0000_0000_0000;
array[18807] <= 16'b0000_0000_0000_0000;
array[18808] <= 16'b0000_0000_0000_0000;
array[18809] <= 16'b0000_0000_0000_0000;
array[18810] <= 16'b0000_0000_0000_0000;
array[18811] <= 16'b0000_0000_0000_0000;
array[18812] <= 16'b0000_0000_0000_0000;
array[18813] <= 16'b0000_0000_0000_0000;
array[18814] <= 16'b0000_0000_0000_0000;
array[18815] <= 16'b0000_0000_0000_0000;
array[18816] <= 16'b0000_0000_0000_0000;
array[18817] <= 16'b0000_0000_0000_0000;
array[18818] <= 16'b0000_0000_0000_0000;
array[18819] <= 16'b0000_0000_0000_0000;
array[18820] <= 16'b0000_0000_0000_0000;
array[18821] <= 16'b0000_0000_0000_0000;
array[18822] <= 16'b0000_0000_0000_0000;
array[18823] <= 16'b0000_0000_0000_0000;
array[18824] <= 16'b0000_0000_0000_0000;
array[18825] <= 16'b0000_0000_0000_0000;
array[18826] <= 16'b0000_0000_0000_0000;
array[18827] <= 16'b0000_0000_0000_0000;
array[18828] <= 16'b0000_0000_0000_0000;
array[18829] <= 16'b0000_0000_0000_0000;
array[18830] <= 16'b0000_0000_0000_0000;
array[18831] <= 16'b0000_0000_0000_0000;
array[18832] <= 16'b0000_0000_0000_0000;
array[18833] <= 16'b0000_0000_0000_0000;
array[18834] <= 16'b0000_0000_0000_0000;
array[18835] <= 16'b0000_0000_0000_0000;
array[18836] <= 16'b0000_0000_0000_0000;
array[18837] <= 16'b0000_0000_0000_0000;
array[18838] <= 16'b0000_0000_0000_0000;
array[18839] <= 16'b0000_0000_0000_0000;
array[18840] <= 16'b0000_0000_0000_0000;
array[18841] <= 16'b0000_0000_0000_0000;
array[18842] <= 16'b0000_0000_0000_0000;
array[18843] <= 16'b0000_0000_0000_0000;
array[18844] <= 16'b0000_0000_0000_0000;
array[18845] <= 16'b0000_0000_0000_0000;
array[18846] <= 16'b0000_0000_0000_0000;
array[18847] <= 16'b0000_0000_0000_0000;
array[18848] <= 16'b0000_0000_0000_0000;
array[18849] <= 16'b0000_0000_0000_0000;
array[18850] <= 16'b0000_0000_0000_0000;
array[18851] <= 16'b0000_0000_0000_0000;
array[18852] <= 16'b0000_0000_0000_0000;
array[18853] <= 16'b0000_0000_0000_0000;
array[18854] <= 16'b0000_0000_0000_0000;
array[18855] <= 16'b0000_0000_0000_0000;
array[18856] <= 16'b0000_0000_0000_0000;
array[18857] <= 16'b0000_0000_0000_0000;
array[18858] <= 16'b0000_0000_0000_0000;
array[18859] <= 16'b0000_0000_0000_0000;
array[18860] <= 16'b0000_0000_0000_0000;
array[18861] <= 16'b0000_0000_0000_0000;
array[18862] <= 16'b0000_0000_0000_0000;
array[18863] <= 16'b0000_0000_0000_0000;
array[18864] <= 16'b0000_0000_0000_0000;
array[18865] <= 16'b0000_0000_0000_0000;
array[18866] <= 16'b0000_0000_0000_0000;
array[18867] <= 16'b0000_0000_0000_0000;
array[18868] <= 16'b0000_0000_0000_0000;
array[18869] <= 16'b0000_0000_0000_0000;
array[18870] <= 16'b0000_0000_0000_0000;
array[18871] <= 16'b0000_0000_0000_0000;
array[18872] <= 16'b0000_0000_0000_0000;
array[18873] <= 16'b0000_0000_0000_0000;
array[18874] <= 16'b0000_0000_0000_0000;
array[18875] <= 16'b0000_0000_0000_0000;
array[18876] <= 16'b0000_0000_0000_0000;
array[18877] <= 16'b0000_0000_0000_0000;
array[18878] <= 16'b0000_0000_0000_0000;
array[18879] <= 16'b0000_0000_0000_0000;
array[18880] <= 16'b0000_0000_0000_0000;
array[18881] <= 16'b0000_0000_0000_0000;
array[18882] <= 16'b0000_0000_0000_0000;
array[18883] <= 16'b0000_0000_0000_0000;
array[18884] <= 16'b0000_0000_0000_0000;
array[18885] <= 16'b0000_0000_0000_0000;
array[18886] <= 16'b0000_0000_0000_0000;
array[18887] <= 16'b0000_0000_0000_0000;
array[18888] <= 16'b0000_0000_0000_0000;
array[18889] <= 16'b0000_0000_0000_0000;
array[18890] <= 16'b0000_0000_0000_0000;
array[18891] <= 16'b0000_0000_0000_0000;
array[18892] <= 16'b0000_0000_0000_0000;
array[18893] <= 16'b0000_0000_0000_0000;
array[18894] <= 16'b0000_0000_0000_0000;
array[18895] <= 16'b0000_0000_0000_0000;
array[18896] <= 16'b0000_0000_0000_0000;
array[18897] <= 16'b0000_0000_0000_0000;
array[18898] <= 16'b0000_0000_0000_0000;
array[18899] <= 16'b0000_0000_0000_0000;
array[18900] <= 16'b0000_0000_0000_0000;
array[18901] <= 16'b0000_0000_0000_0000;
array[18902] <= 16'b0000_0000_0000_0000;
array[18903] <= 16'b0000_0000_0000_0000;
array[18904] <= 16'b0000_0000_0000_0000;
array[18905] <= 16'b0000_0000_0000_0000;
array[18906] <= 16'b0000_0000_0000_0000;
array[18907] <= 16'b0000_0000_0000_0000;
array[18908] <= 16'b0000_0000_0000_0000;
array[18909] <= 16'b0000_0000_0000_0000;
array[18910] <= 16'b0000_0000_0000_0000;
array[18911] <= 16'b0000_0000_0000_0000;
array[18912] <= 16'b0000_0000_0000_0000;
array[18913] <= 16'b0000_0000_0000_0000;
array[18914] <= 16'b0000_0000_0000_0000;
array[18915] <= 16'b0000_0000_0000_0000;
array[18916] <= 16'b0000_0000_0000_0000;
array[18917] <= 16'b0000_0000_0000_0000;
array[18918] <= 16'b0000_0000_0000_0000;
array[18919] <= 16'b0000_0000_0000_0000;
array[18920] <= 16'b0000_0000_0000_0000;
array[18921] <= 16'b0000_0000_0000_0000;
array[18922] <= 16'b0000_0000_0000_0000;
array[18923] <= 16'b0000_0000_0000_0000;
array[18924] <= 16'b0000_0000_0000_0000;
array[18925] <= 16'b0000_0000_0000_0000;
array[18926] <= 16'b0000_0000_0000_0000;
array[18927] <= 16'b0000_0000_0000_0000;
array[18928] <= 16'b0000_0000_0000_0000;
array[18929] <= 16'b0000_0000_0000_0000;
array[18930] <= 16'b0000_0000_0000_0000;
array[18931] <= 16'b0000_0000_0000_0000;
array[18932] <= 16'b0000_0000_0000_0000;
array[18933] <= 16'b0000_0000_0000_0000;
array[18934] <= 16'b0000_0000_0000_0000;
array[18935] <= 16'b0000_0000_0000_0000;
array[18936] <= 16'b0000_0000_0000_0000;
array[18937] <= 16'b0000_0000_0000_0000;
array[18938] <= 16'b0000_0000_0000_0000;
array[18939] <= 16'b0000_0000_0000_0000;
array[18940] <= 16'b0000_0000_0000_0000;
array[18941] <= 16'b0000_0000_0000_0000;
array[18942] <= 16'b0000_0000_0000_0000;
array[18943] <= 16'b0000_0000_0000_0000;
array[18944] <= 16'b0000_0000_0000_0000;
array[18945] <= 16'b0000_0000_0000_0000;
array[18946] <= 16'b0000_0000_0000_0000;
array[18947] <= 16'b0000_0000_0000_0000;
array[18948] <= 16'b0000_0000_0000_0000;
array[18949] <= 16'b0000_0000_0000_0000;
array[18950] <= 16'b0000_0000_0000_0000;
array[18951] <= 16'b0000_0000_0000_0000;
array[18952] <= 16'b0000_0000_0000_0000;
array[18953] <= 16'b0000_0000_0000_0000;
array[18954] <= 16'b0000_0000_0000_0000;
array[18955] <= 16'b0000_0000_0000_0000;
array[18956] <= 16'b0000_0000_0000_0000;
array[18957] <= 16'b0000_0000_0000_0000;
array[18958] <= 16'b0000_0000_0000_0000;
array[18959] <= 16'b0000_0000_0000_0000;
array[18960] <= 16'b0000_0000_0000_0000;
array[18961] <= 16'b0000_0000_0000_0000;
array[18962] <= 16'b0000_0000_0000_0000;
array[18963] <= 16'b0000_0000_0000_0000;
array[18964] <= 16'b0000_0000_0000_0000;
array[18965] <= 16'b0000_0000_0000_0000;
array[18966] <= 16'b0000_0000_0000_0000;
array[18967] <= 16'b0000_0000_0000_0000;
array[18968] <= 16'b0000_0000_0000_0000;
array[18969] <= 16'b0000_0000_0000_0000;
array[18970] <= 16'b0000_0000_0000_0000;
array[18971] <= 16'b0000_0000_0000_0000;
array[18972] <= 16'b0000_0000_0000_0000;
array[18973] <= 16'b0000_0000_0000_0000;
array[18974] <= 16'b0000_0000_0000_0000;
array[18975] <= 16'b0000_0000_0000_0000;
array[18976] <= 16'b0000_0000_0000_0000;
array[18977] <= 16'b0000_0000_0000_0000;
array[18978] <= 16'b0000_0000_0000_0000;
array[18979] <= 16'b0000_0000_0000_0000;
array[18980] <= 16'b0000_0000_0000_0000;
array[18981] <= 16'b0000_0000_0000_0000;
array[18982] <= 16'b0000_0000_0000_0000;
array[18983] <= 16'b0000_0000_0000_0000;
array[18984] <= 16'b0000_0000_0000_0000;
array[18985] <= 16'b0000_0000_0000_0000;
array[18986] <= 16'b0000_0000_0000_0000;
array[18987] <= 16'b0000_0000_0000_0000;
array[18988] <= 16'b0000_0000_0000_0000;
array[18989] <= 16'b0000_0000_0000_0000;
array[18990] <= 16'b0000_0000_0000_0000;
array[18991] <= 16'b0000_0000_0000_0000;
array[18992] <= 16'b0000_0000_0000_0000;
array[18993] <= 16'b0000_0000_0000_0000;
array[18994] <= 16'b0000_0000_0000_0000;
array[18995] <= 16'b0000_0000_0000_0000;
array[18996] <= 16'b0000_0000_0000_0000;
array[18997] <= 16'b0000_0000_0000_0000;
array[18998] <= 16'b0000_0000_0000_0000;
array[18999] <= 16'b0000_0000_0000_0000;
array[19000] <= 16'b0000_0000_0000_0000;
array[19001] <= 16'b0000_0000_0000_0000;
array[19002] <= 16'b0000_0000_0000_0000;
array[19003] <= 16'b0000_0000_0000_0000;
array[19004] <= 16'b0000_0000_0000_0000;
array[19005] <= 16'b0000_0000_0000_0000;
array[19006] <= 16'b0000_0000_0000_0000;
array[19007] <= 16'b0000_0000_0000_0000;
array[19008] <= 16'b0000_0000_0000_0000;
array[19009] <= 16'b0000_0000_0000_0000;
array[19010] <= 16'b0000_0000_0000_0000;
array[19011] <= 16'b0000_0000_0000_0000;
array[19012] <= 16'b0000_0000_0000_0000;
array[19013] <= 16'b0000_0000_0000_0000;
array[19014] <= 16'b0000_0000_0000_0000;
array[19015] <= 16'b0000_0000_0000_0000;
array[19016] <= 16'b0000_0000_0000_0000;
array[19017] <= 16'b0000_0000_0000_0000;
array[19018] <= 16'b0000_0000_0000_0000;
array[19019] <= 16'b0000_0000_0000_0000;
array[19020] <= 16'b0000_0000_0000_0000;
array[19021] <= 16'b0000_0000_0000_0000;
array[19022] <= 16'b0000_0000_0000_0000;
array[19023] <= 16'b0000_0000_0000_0000;
array[19024] <= 16'b0000_0000_0000_0000;
array[19025] <= 16'b0000_0000_0000_0000;
array[19026] <= 16'b0000_0000_0000_0000;
array[19027] <= 16'b0000_0000_0000_0000;
array[19028] <= 16'b0000_0000_0000_0000;
array[19029] <= 16'b0000_0000_0000_0000;
array[19030] <= 16'b0000_0000_0000_0000;
array[19031] <= 16'b0000_0000_0000_0000;
array[19032] <= 16'b0000_0000_0000_0000;
array[19033] <= 16'b0000_0000_0000_0000;
array[19034] <= 16'b0000_0000_0000_0000;
array[19035] <= 16'b0000_0000_0000_0000;
array[19036] <= 16'b0000_0000_0000_0000;
array[19037] <= 16'b0000_0000_0000_0000;
array[19038] <= 16'b0000_0000_0000_0000;
array[19039] <= 16'b0000_0000_0000_0000;
array[19040] <= 16'b0000_0000_0000_0000;
array[19041] <= 16'b0000_0000_0000_0000;
array[19042] <= 16'b0000_0000_0000_0000;
array[19043] <= 16'b0000_0000_0000_0000;
array[19044] <= 16'b0000_0000_0000_0000;
array[19045] <= 16'b0000_0000_0000_0000;
array[19046] <= 16'b0000_0000_0000_0000;
array[19047] <= 16'b0000_0000_0000_0000;
array[19048] <= 16'b0000_0000_0000_0000;
array[19049] <= 16'b0000_0000_0000_0000;
array[19050] <= 16'b0000_0000_0000_0000;
array[19051] <= 16'b0000_0000_0000_0000;
array[19052] <= 16'b0000_0000_0000_0000;
array[19053] <= 16'b0000_0000_0000_0000;
array[19054] <= 16'b0000_0000_0000_0000;
array[19055] <= 16'b0000_0000_0000_0000;
array[19056] <= 16'b0000_0000_0000_0000;
array[19057] <= 16'b0000_0000_0000_0000;
array[19058] <= 16'b0000_0000_0000_0000;
array[19059] <= 16'b0000_0000_0000_0000;
array[19060] <= 16'b0000_0000_0000_0000;
array[19061] <= 16'b0000_0000_0000_0000;
array[19062] <= 16'b0000_0000_0000_0000;
array[19063] <= 16'b0000_0000_0000_0000;
array[19064] <= 16'b0000_0000_0000_0000;
array[19065] <= 16'b0000_0000_0000_0000;
array[19066] <= 16'b0000_0000_0000_0000;
array[19067] <= 16'b0000_0000_0000_0000;
array[19068] <= 16'b0000_0000_0000_0000;
array[19069] <= 16'b0000_0000_0000_0000;
array[19070] <= 16'b0000_0000_0000_0000;
array[19071] <= 16'b0000_0000_0000_0000;
array[19072] <= 16'b0000_0000_0000_0000;
array[19073] <= 16'b0000_0000_0000_0000;
array[19074] <= 16'b0000_0000_0000_0000;
array[19075] <= 16'b0000_0000_0000_0000;
array[19076] <= 16'b0000_0000_0000_0000;
array[19077] <= 16'b0000_0000_0000_0000;
array[19078] <= 16'b0000_0000_0000_0000;
array[19079] <= 16'b0000_0000_0000_0000;
array[19080] <= 16'b0000_0000_0000_0000;
array[19081] <= 16'b0000_0000_0000_0000;
array[19082] <= 16'b0000_0000_0000_0000;
array[19083] <= 16'b0000_0000_0000_0000;
array[19084] <= 16'b0000_0000_0000_0000;
array[19085] <= 16'b0000_0000_0000_0000;
array[19086] <= 16'b0000_0000_0000_0000;
array[19087] <= 16'b0000_0000_0000_0000;
array[19088] <= 16'b0000_0000_0000_0000;
array[19089] <= 16'b0000_0000_0000_0000;
array[19090] <= 16'b0000_0000_0000_0000;
array[19091] <= 16'b0000_0000_0000_0000;
array[19092] <= 16'b0000_0000_0000_0000;
array[19093] <= 16'b0000_0000_0000_0000;
array[19094] <= 16'b0000_0000_0000_0000;
array[19095] <= 16'b0000_0000_0000_0000;
array[19096] <= 16'b0000_0000_0000_0000;
array[19097] <= 16'b0000_0000_0000_0000;
array[19098] <= 16'b0000_0000_0000_0000;
array[19099] <= 16'b0000_0000_0000_0000;
array[19100] <= 16'b0000_0000_0000_0000;
array[19101] <= 16'b0000_0000_0000_0000;
array[19102] <= 16'b0000_0000_0000_0000;
array[19103] <= 16'b0000_0000_0000_0000;
array[19104] <= 16'b0000_0000_0000_0000;
array[19105] <= 16'b0000_0000_0000_0000;
array[19106] <= 16'b0000_0000_0000_0000;
array[19107] <= 16'b0000_0000_0000_0000;
array[19108] <= 16'b0000_0000_0000_0000;
array[19109] <= 16'b0000_0000_0000_0000;
array[19110] <= 16'b0000_0000_0000_0000;
array[19111] <= 16'b0000_0000_0000_0000;
array[19112] <= 16'b0000_0000_0000_0000;
array[19113] <= 16'b0000_0000_0000_0000;
array[19114] <= 16'b0000_0000_0000_0000;
array[19115] <= 16'b0000_0000_0000_0000;
array[19116] <= 16'b0000_0000_0000_0000;
array[19117] <= 16'b0000_0000_0000_0000;
array[19118] <= 16'b0000_0000_0000_0000;
array[19119] <= 16'b0000_0000_0000_0000;
array[19120] <= 16'b0000_0000_0000_0000;
array[19121] <= 16'b0000_0000_0000_0000;
array[19122] <= 16'b0000_0000_0000_0000;
array[19123] <= 16'b0000_0000_0000_0000;
array[19124] <= 16'b0000_0000_0000_0000;
array[19125] <= 16'b0000_0000_0000_0000;
array[19126] <= 16'b0000_0000_0000_0000;
array[19127] <= 16'b0000_0000_0000_0000;
array[19128] <= 16'b0000_0000_0000_0000;
array[19129] <= 16'b0000_0000_0000_0000;
array[19130] <= 16'b0000_0000_0000_0000;
array[19131] <= 16'b0000_0000_0000_0000;
array[19132] <= 16'b0000_0000_0000_0000;
array[19133] <= 16'b0000_0000_0000_0000;
array[19134] <= 16'b0000_0000_0000_0000;
array[19135] <= 16'b0000_0000_0000_0000;
array[19136] <= 16'b0000_0000_0000_0000;
array[19137] <= 16'b0000_0000_0000_0000;
array[19138] <= 16'b0000_0000_0000_0000;
array[19139] <= 16'b0000_0000_0000_0000;
array[19140] <= 16'b0000_0000_0000_0000;
array[19141] <= 16'b0000_0000_0000_0000;
array[19142] <= 16'b0000_0000_0000_0000;
array[19143] <= 16'b0000_0000_0000_0000;
array[19144] <= 16'b0000_0000_0000_0000;
array[19145] <= 16'b0000_0000_0000_0000;
array[19146] <= 16'b0000_0000_0000_0000;
array[19147] <= 16'b0000_0000_0000_0000;
array[19148] <= 16'b0000_0000_0000_0000;
array[19149] <= 16'b0000_0000_0000_0000;
array[19150] <= 16'b0000_0000_0000_0000;
array[19151] <= 16'b0000_0000_0000_0000;
array[19152] <= 16'b0000_0000_0000_0000;
array[19153] <= 16'b0000_0000_0000_0000;
array[19154] <= 16'b0000_0000_0000_0000;
array[19155] <= 16'b0000_0000_0000_0000;
array[19156] <= 16'b0000_0000_0000_0000;
array[19157] <= 16'b0000_0000_0000_0000;
array[19158] <= 16'b0000_0000_0000_0000;
array[19159] <= 16'b0000_0000_0000_0000;
array[19160] <= 16'b0000_0000_0000_0000;
array[19161] <= 16'b0000_0000_0000_0000;
array[19162] <= 16'b0000_0000_0000_0000;
array[19163] <= 16'b0000_0000_0000_0000;
array[19164] <= 16'b0000_0000_0000_0000;
array[19165] <= 16'b0000_0000_0000_0000;
array[19166] <= 16'b0000_0000_0000_0000;
array[19167] <= 16'b0000_0000_0000_0000;
array[19168] <= 16'b0000_0000_0000_0000;
array[19169] <= 16'b0000_0000_0000_0000;
array[19170] <= 16'b0000_0000_0000_0000;
array[19171] <= 16'b0000_0000_0000_0000;
array[19172] <= 16'b0000_0000_0000_0000;
array[19173] <= 16'b0000_0000_0000_0000;
array[19174] <= 16'b0000_0000_0000_0000;
array[19175] <= 16'b0000_0000_0000_0000;
array[19176] <= 16'b0000_0000_0000_0000;
array[19177] <= 16'b0000_0000_0000_0000;
array[19178] <= 16'b0000_0000_0000_0000;
array[19179] <= 16'b0000_0000_0000_0000;
array[19180] <= 16'b0000_0000_0000_0000;
array[19181] <= 16'b0000_0000_0000_0000;
array[19182] <= 16'b0000_0000_0000_0000;
array[19183] <= 16'b0000_0000_0000_0000;
array[19184] <= 16'b0000_0000_0000_0000;
array[19185] <= 16'b0000_0000_0000_0000;
array[19186] <= 16'b0000_0000_0000_0000;
array[19187] <= 16'b0000_0000_0000_0000;
array[19188] <= 16'b0000_0000_0000_0000;
array[19189] <= 16'b0000_0000_0000_0000;
array[19190] <= 16'b0000_0000_0000_0000;
array[19191] <= 16'b0000_0000_0000_0000;
array[19192] <= 16'b0000_0000_0000_0000;
array[19193] <= 16'b0000_0000_0000_0000;
array[19194] <= 16'b0000_0000_0000_0000;
array[19195] <= 16'b0000_0000_0000_0000;
array[19196] <= 16'b0000_0000_0000_0000;
array[19197] <= 16'b0000_0000_0000_0000;
array[19198] <= 16'b0000_0000_0000_0000;
array[19199] <= 16'b0000_0000_0000_0000;
array[19200] <= 16'b0000_0000_0000_0000;
array[19201] <= 16'b0000_0000_0000_0000;
array[19202] <= 16'b0000_0000_0000_0000;
array[19203] <= 16'b0000_0000_0000_0000;
array[19204] <= 16'b0000_0000_0000_0000;
array[19205] <= 16'b0000_0000_0000_0000;
array[19206] <= 16'b0000_0000_0000_0000;
array[19207] <= 16'b0000_0000_0000_0000;
array[19208] <= 16'b0000_0000_0000_0000;
array[19209] <= 16'b0000_0000_0000_0000;
array[19210] <= 16'b0000_0000_0000_0000;
array[19211] <= 16'b0000_0000_0000_0000;
array[19212] <= 16'b0000_0000_0000_0000;
array[19213] <= 16'b0000_0000_0000_0000;
array[19214] <= 16'b0000_0000_0000_0000;
array[19215] <= 16'b0000_0000_0000_0000;
array[19216] <= 16'b0000_0000_0000_0000;
array[19217] <= 16'b0000_0000_0000_0000;
array[19218] <= 16'b0000_0000_0000_0000;
array[19219] <= 16'b0000_0000_0000_0000;
array[19220] <= 16'b0000_0000_0000_0000;
array[19221] <= 16'b0000_0000_0000_0000;
array[19222] <= 16'b0000_0000_0000_0000;
array[19223] <= 16'b0000_0000_0000_0000;
array[19224] <= 16'b0000_0000_0000_0000;
array[19225] <= 16'b0000_0000_0000_0000;
array[19226] <= 16'b0000_0000_0000_0000;
array[19227] <= 16'b0000_0000_0000_0000;
array[19228] <= 16'b0000_0000_0000_0000;
array[19229] <= 16'b0000_0000_0000_0000;
array[19230] <= 16'b0000_0000_0000_0000;
array[19231] <= 16'b0000_0000_0000_0000;
array[19232] <= 16'b0000_0000_0000_0000;
array[19233] <= 16'b0000_0000_0000_0000;
array[19234] <= 16'b0000_0000_0000_0000;
array[19235] <= 16'b0000_0000_0000_0000;
array[19236] <= 16'b0000_0000_0000_0000;
array[19237] <= 16'b0000_0000_0000_0000;
array[19238] <= 16'b0000_0000_0000_0000;
array[19239] <= 16'b0000_0000_0000_0000;
array[19240] <= 16'b0000_0000_0000_0000;
array[19241] <= 16'b0000_0000_0000_0000;
array[19242] <= 16'b0000_0000_0000_0000;
array[19243] <= 16'b0000_0000_0000_0000;
array[19244] <= 16'b0000_0000_0000_0000;
array[19245] <= 16'b0000_0000_0000_0000;
array[19246] <= 16'b0000_0000_0000_0000;
array[19247] <= 16'b0000_0000_0000_0000;
array[19248] <= 16'b0000_0000_0000_0000;
array[19249] <= 16'b0000_0000_0000_0000;
array[19250] <= 16'b0000_0000_0000_0000;
array[19251] <= 16'b0000_0000_0000_0000;
array[19252] <= 16'b0000_0000_0000_0000;
array[19253] <= 16'b0000_0000_0000_0000;
array[19254] <= 16'b0000_0000_0000_0000;
array[19255] <= 16'b0000_0000_0000_0000;
array[19256] <= 16'b0000_0000_0000_0000;
array[19257] <= 16'b0000_0000_0000_0000;
array[19258] <= 16'b0000_0000_0000_0000;
array[19259] <= 16'b0000_0000_0000_0000;
array[19260] <= 16'b0000_0000_0000_0000;
array[19261] <= 16'b0000_0000_0000_0000;
array[19262] <= 16'b0000_0000_0000_0000;
array[19263] <= 16'b0000_0000_0000_0000;
array[19264] <= 16'b0000_0000_0000_0000;
array[19265] <= 16'b0000_0000_0000_0000;
array[19266] <= 16'b0000_0000_0000_0000;
array[19267] <= 16'b0000_0000_0000_0000;
array[19268] <= 16'b0000_0000_0000_0000;
array[19269] <= 16'b0000_0000_0000_0000;
array[19270] <= 16'b0000_0000_0000_0000;
array[19271] <= 16'b0000_0000_0000_0000;
array[19272] <= 16'b0000_0000_0000_0000;
array[19273] <= 16'b0000_0000_0000_0000;
array[19274] <= 16'b0000_0000_0000_0000;
array[19275] <= 16'b0000_0000_0000_0000;
array[19276] <= 16'b0000_0000_0000_0000;
array[19277] <= 16'b0000_0000_0000_0000;
array[19278] <= 16'b0000_0000_0000_0000;
array[19279] <= 16'b0000_0000_0000_0000;
array[19280] <= 16'b0000_0000_0000_0000;
array[19281] <= 16'b0000_0000_0000_0000;
array[19282] <= 16'b0000_0000_0000_0000;
array[19283] <= 16'b0000_0000_0000_0000;
array[19284] <= 16'b0000_0000_0000_0000;
array[19285] <= 16'b0000_0000_0000_0000;
array[19286] <= 16'b0000_0000_0000_0000;
array[19287] <= 16'b0000_0000_0000_0000;
array[19288] <= 16'b0000_0000_0000_0000;
array[19289] <= 16'b0000_0000_0000_0000;
array[19290] <= 16'b0000_0000_0000_0000;
array[19291] <= 16'b0000_0000_0000_0000;
array[19292] <= 16'b0000_0000_0000_0000;
array[19293] <= 16'b0000_0000_0000_0000;
array[19294] <= 16'b0000_0000_0000_0000;
array[19295] <= 16'b0000_0000_0000_0000;
array[19296] <= 16'b0000_0000_0000_0000;
array[19297] <= 16'b0000_0000_0000_0000;
array[19298] <= 16'b0000_0000_0000_0000;
array[19299] <= 16'b0000_0000_0000_0000;
array[19300] <= 16'b0000_0000_0000_0000;
array[19301] <= 16'b0000_0000_0000_0000;
array[19302] <= 16'b0000_0000_0000_0000;
array[19303] <= 16'b0000_0000_0000_0000;
array[19304] <= 16'b0000_0000_0000_0000;
array[19305] <= 16'b0000_0000_0000_0000;
array[19306] <= 16'b0000_0000_0000_0000;
array[19307] <= 16'b0000_0000_0000_0000;
array[19308] <= 16'b0000_0000_0000_0000;
array[19309] <= 16'b0000_0000_0000_0000;
array[19310] <= 16'b0000_0000_0000_0000;
array[19311] <= 16'b0000_0000_0000_0000;
array[19312] <= 16'b0000_0000_0000_0000;
array[19313] <= 16'b0000_0000_0000_0000;
array[19314] <= 16'b0000_0000_0000_0000;
array[19315] <= 16'b0000_0000_0000_0000;
array[19316] <= 16'b0000_0000_0000_0000;
array[19317] <= 16'b0000_0000_0000_0000;
array[19318] <= 16'b0000_0000_0000_0000;
array[19319] <= 16'b0000_0000_0000_0000;
array[19320] <= 16'b0000_0000_0000_0000;
array[19321] <= 16'b0000_0000_0000_0000;
array[19322] <= 16'b0000_0000_0000_0000;
array[19323] <= 16'b0000_0000_0000_0000;
array[19324] <= 16'b0000_0000_0000_0000;
array[19325] <= 16'b0000_0000_0000_0000;
array[19326] <= 16'b0000_0000_0000_0000;
array[19327] <= 16'b0000_0000_0000_0000;
array[19328] <= 16'b0000_0000_0000_0000;
array[19329] <= 16'b0000_0000_0000_0000;
array[19330] <= 16'b0000_0000_0000_0000;
array[19331] <= 16'b0000_0000_0000_0000;
array[19332] <= 16'b0000_0000_0000_0000;
array[19333] <= 16'b0000_0000_0000_0000;
array[19334] <= 16'b0000_0000_0000_0000;
array[19335] <= 16'b0000_0000_0000_0000;
array[19336] <= 16'b0000_0000_0000_0000;
array[19337] <= 16'b0000_0000_0000_0000;
array[19338] <= 16'b0000_0000_0000_0000;
array[19339] <= 16'b0000_0000_0000_0000;
array[19340] <= 16'b0000_0000_0000_0000;
array[19341] <= 16'b0000_0000_0000_0000;
array[19342] <= 16'b0000_0000_0000_0000;
array[19343] <= 16'b0000_0000_0000_0000;
array[19344] <= 16'b0000_0000_0000_0000;
array[19345] <= 16'b0000_0000_0000_0000;
array[19346] <= 16'b0000_0000_0000_0000;
array[19347] <= 16'b0000_0000_0000_0000;
array[19348] <= 16'b0000_0000_0000_0000;
array[19349] <= 16'b0000_0000_0000_0000;
array[19350] <= 16'b0000_0000_0000_0000;
array[19351] <= 16'b0000_0000_0000_0000;
array[19352] <= 16'b0000_0000_0000_0000;
array[19353] <= 16'b0000_0000_0000_0000;
array[19354] <= 16'b0000_0000_0000_0000;
array[19355] <= 16'b0000_0000_0000_0000;
array[19356] <= 16'b0000_0000_0000_0000;
array[19357] <= 16'b0000_0000_0000_0000;
array[19358] <= 16'b0000_0000_0000_0000;
array[19359] <= 16'b0000_0000_0000_0000;
array[19360] <= 16'b0000_0000_0000_0000;
array[19361] <= 16'b0000_0000_0000_0000;
array[19362] <= 16'b0000_0000_0000_0000;
array[19363] <= 16'b0000_0000_0000_0000;
array[19364] <= 16'b0000_0000_0000_0000;
array[19365] <= 16'b0000_0000_0000_0000;
array[19366] <= 16'b0000_0000_0000_0000;
array[19367] <= 16'b0000_0000_0000_0000;
array[19368] <= 16'b0000_0000_0000_0000;
array[19369] <= 16'b0000_0000_0000_0000;
array[19370] <= 16'b0000_0000_0000_0000;
array[19371] <= 16'b0000_0000_0000_0000;
array[19372] <= 16'b0000_0000_0000_0000;
array[19373] <= 16'b0000_0000_0000_0000;
array[19374] <= 16'b0000_0000_0000_0000;
array[19375] <= 16'b0000_0000_0000_0000;
array[19376] <= 16'b0000_0000_0000_0000;
array[19377] <= 16'b0000_0000_0000_0000;
array[19378] <= 16'b0000_0000_0000_0000;
array[19379] <= 16'b0000_0000_0000_0000;
array[19380] <= 16'b0000_0000_0000_0000;
array[19381] <= 16'b0000_0000_0000_0000;
array[19382] <= 16'b0000_0000_0000_0000;
array[19383] <= 16'b0000_0000_0000_0000;
array[19384] <= 16'b0000_0000_0000_0000;
array[19385] <= 16'b0000_0000_0000_0000;
array[19386] <= 16'b0000_0000_0000_0000;
array[19387] <= 16'b0000_0000_0000_0000;
array[19388] <= 16'b0000_0000_0000_0000;
array[19389] <= 16'b0000_0000_0000_0000;
array[19390] <= 16'b0000_0000_0000_0000;
array[19391] <= 16'b0000_0000_0000_0000;
array[19392] <= 16'b0000_0000_0000_0000;
array[19393] <= 16'b0000_0000_0000_0000;
array[19394] <= 16'b0000_0000_0000_0000;
array[19395] <= 16'b0000_0000_0000_0000;
array[19396] <= 16'b0000_0000_0000_0000;
array[19397] <= 16'b0000_0000_0000_0000;
array[19398] <= 16'b0000_0000_0000_0000;
array[19399] <= 16'b0000_0000_0000_0000;
array[19400] <= 16'b0000_0000_0000_0000;
array[19401] <= 16'b0000_0000_0000_0000;
array[19402] <= 16'b0000_0000_0000_0000;
array[19403] <= 16'b0000_0000_0000_0000;
array[19404] <= 16'b0000_0000_0000_0000;
array[19405] <= 16'b0000_0000_0000_0000;
array[19406] <= 16'b0000_0000_0000_0000;
array[19407] <= 16'b0000_0000_0000_0000;
array[19408] <= 16'b0000_0000_0000_0000;
array[19409] <= 16'b0000_0000_0000_0000;
array[19410] <= 16'b0000_0000_0000_0000;
array[19411] <= 16'b0000_0000_0000_0000;
array[19412] <= 16'b0000_0000_0000_0000;
array[19413] <= 16'b0000_0000_0000_0000;
array[19414] <= 16'b0000_0000_0000_0000;
array[19415] <= 16'b0000_0000_0000_0000;
array[19416] <= 16'b0000_0000_0000_0000;
array[19417] <= 16'b0000_0000_0000_0000;
array[19418] <= 16'b0000_0000_0000_0000;
array[19419] <= 16'b0000_0000_0000_0000;
array[19420] <= 16'b0000_0000_0000_0000;
array[19421] <= 16'b0000_0000_0000_0000;
array[19422] <= 16'b0000_0000_0000_0000;
array[19423] <= 16'b0000_0000_0000_0000;
array[19424] <= 16'b0000_0000_0000_0000;
array[19425] <= 16'b0000_0000_0000_0000;
array[19426] <= 16'b0000_0000_0000_0000;
array[19427] <= 16'b0000_0000_0000_0000;
array[19428] <= 16'b0000_0000_0000_0000;
array[19429] <= 16'b0000_0000_0000_0000;
array[19430] <= 16'b0000_0000_0000_0000;
array[19431] <= 16'b0000_0000_0000_0000;
array[19432] <= 16'b0000_0000_0000_0000;
array[19433] <= 16'b0000_0000_0000_0000;
array[19434] <= 16'b0000_0000_0000_0000;
array[19435] <= 16'b0000_0000_0000_0000;
array[19436] <= 16'b0000_0000_0000_0000;
array[19437] <= 16'b0000_0000_0000_0000;
array[19438] <= 16'b0000_0000_0000_0000;
array[19439] <= 16'b0000_0000_0000_0000;
array[19440] <= 16'b0000_0000_0000_0000;
array[19441] <= 16'b0000_0000_0000_0000;
array[19442] <= 16'b0000_0000_0000_0000;
array[19443] <= 16'b0000_0000_0000_0000;
array[19444] <= 16'b0000_0000_0000_0000;
array[19445] <= 16'b0000_0000_0000_0000;
array[19446] <= 16'b0000_0000_0000_0000;
array[19447] <= 16'b0000_0000_0000_0000;
array[19448] <= 16'b0000_0000_0000_0000;
array[19449] <= 16'b0000_0000_0000_0000;
array[19450] <= 16'b0000_0000_0000_0000;
array[19451] <= 16'b0000_0000_0000_0000;
array[19452] <= 16'b0000_0000_0000_0000;
array[19453] <= 16'b0000_0000_0000_0000;
array[19454] <= 16'b0000_0000_0000_0000;
array[19455] <= 16'b0000_0000_0000_0000;
array[19456] <= 16'b0000_0000_0000_0000;
array[19457] <= 16'b0000_0000_0000_0000;
array[19458] <= 16'b0000_0000_0000_0000;
array[19459] <= 16'b0000_0000_0000_0000;
array[19460] <= 16'b0000_0000_0000_0000;
array[19461] <= 16'b0000_0000_0000_0000;
array[19462] <= 16'b0000_0000_0000_0000;
array[19463] <= 16'b0000_0000_0000_0000;
array[19464] <= 16'b0000_0000_0000_0000;
array[19465] <= 16'b0000_0000_0000_0000;
array[19466] <= 16'b0000_0000_0000_0000;
array[19467] <= 16'b0000_0000_0000_0000;
array[19468] <= 16'b0000_0000_0000_0000;
array[19469] <= 16'b0000_0000_0000_0000;
array[19470] <= 16'b0000_0000_0000_0000;
array[19471] <= 16'b0000_0000_0000_0000;
array[19472] <= 16'b0000_0000_0000_0000;
array[19473] <= 16'b0000_0000_0000_0000;
array[19474] <= 16'b0000_0000_0000_0000;
array[19475] <= 16'b0000_0000_0000_0000;
array[19476] <= 16'b0000_0000_0000_0000;
array[19477] <= 16'b0000_0000_0000_0000;
array[19478] <= 16'b0000_0000_0000_0000;
array[19479] <= 16'b0000_0000_0000_0000;
array[19480] <= 16'b0000_0000_0000_0000;
array[19481] <= 16'b0000_0000_0000_0000;
array[19482] <= 16'b0000_0000_0000_0000;
array[19483] <= 16'b0000_0000_0000_0000;
array[19484] <= 16'b0000_0000_0000_0000;
array[19485] <= 16'b0000_0000_0000_0000;
array[19486] <= 16'b0000_0000_0000_0000;
array[19487] <= 16'b0000_0000_0000_0000;
array[19488] <= 16'b0000_0000_0000_0000;
array[19489] <= 16'b0000_0000_0000_0000;
array[19490] <= 16'b0000_0000_0000_0000;
array[19491] <= 16'b0000_0000_0000_0000;
array[19492] <= 16'b0000_0000_0000_0000;
array[19493] <= 16'b0000_0000_0000_0000;
array[19494] <= 16'b0000_0000_0000_0000;
array[19495] <= 16'b0000_0000_0000_0000;
array[19496] <= 16'b0000_0000_0000_0000;
array[19497] <= 16'b0000_0000_0000_0000;
array[19498] <= 16'b0000_0000_0000_0000;
array[19499] <= 16'b0000_0000_0000_0000;
array[19500] <= 16'b0000_0000_0000_0000;
array[19501] <= 16'b0000_0000_0000_0000;
array[19502] <= 16'b0000_0000_0000_0000;
array[19503] <= 16'b0000_0000_0000_0000;
array[19504] <= 16'b0000_0000_0000_0000;
array[19505] <= 16'b0000_0000_0000_0000;
array[19506] <= 16'b0000_0000_0000_0000;
array[19507] <= 16'b0000_0000_0000_0000;
array[19508] <= 16'b0000_0000_0000_0000;
array[19509] <= 16'b0000_0000_0000_0000;
array[19510] <= 16'b0000_0000_0000_0000;
array[19511] <= 16'b0000_0000_0000_0000;
array[19512] <= 16'b0000_0000_0000_0000;
array[19513] <= 16'b0000_0000_0000_0000;
array[19514] <= 16'b0000_0000_0000_0000;
array[19515] <= 16'b0000_0000_0000_0000;
array[19516] <= 16'b0000_0000_0000_0000;
array[19517] <= 16'b0000_0000_0000_0000;
array[19518] <= 16'b0000_0000_0000_0000;
array[19519] <= 16'b0000_0000_0000_0000;
array[19520] <= 16'b0000_0000_0000_0000;
array[19521] <= 16'b0000_0000_0000_0000;
array[19522] <= 16'b0000_0000_0000_0000;
array[19523] <= 16'b0000_0000_0000_0000;
array[19524] <= 16'b0000_0000_0000_0000;
array[19525] <= 16'b0000_0000_0000_0000;
array[19526] <= 16'b0000_0000_0000_0000;
array[19527] <= 16'b0000_0000_0000_0000;
array[19528] <= 16'b0000_0000_0000_0000;
array[19529] <= 16'b0000_0000_0000_0000;
array[19530] <= 16'b0000_0000_0000_0000;
array[19531] <= 16'b0000_0000_0000_0000;
array[19532] <= 16'b0000_0000_0000_0000;
array[19533] <= 16'b0000_0000_0000_0000;
array[19534] <= 16'b0000_0000_0000_0000;
array[19535] <= 16'b0000_0000_0000_0000;
array[19536] <= 16'b0000_0000_0000_0000;
array[19537] <= 16'b0000_0000_0000_0000;
array[19538] <= 16'b0000_0000_0000_0000;
array[19539] <= 16'b0000_0000_0000_0000;
array[19540] <= 16'b0000_0000_0000_0000;
array[19541] <= 16'b0000_0000_0000_0000;
array[19542] <= 16'b0000_0000_0000_0000;
array[19543] <= 16'b0000_0000_0000_0000;
array[19544] <= 16'b0000_0000_0000_0000;
array[19545] <= 16'b0000_0000_0000_0000;
array[19546] <= 16'b0000_0000_0000_0000;
array[19547] <= 16'b0000_0000_0000_0000;
array[19548] <= 16'b0000_0000_0000_0000;
array[19549] <= 16'b0000_0000_0000_0000;
array[19550] <= 16'b0000_0000_0000_0000;
array[19551] <= 16'b0000_0000_0000_0000;
array[19552] <= 16'b0000_0000_0000_0000;
array[19553] <= 16'b0000_0000_0000_0000;
array[19554] <= 16'b0000_0000_0000_0000;
array[19555] <= 16'b0000_0000_0000_0000;
array[19556] <= 16'b0000_0000_0000_0000;
array[19557] <= 16'b0000_0000_0000_0000;
array[19558] <= 16'b0000_0000_0000_0000;
array[19559] <= 16'b0000_0000_0000_0000;
array[19560] <= 16'b0000_0000_0000_0000;
array[19561] <= 16'b0000_0000_0000_0000;
array[19562] <= 16'b0000_0000_0000_0000;
array[19563] <= 16'b0000_0000_0000_0000;
array[19564] <= 16'b0000_0000_0000_0000;
array[19565] <= 16'b0000_0000_0000_0000;
array[19566] <= 16'b0000_0000_0000_0000;
array[19567] <= 16'b0000_0000_0000_0000;
array[19568] <= 16'b0000_0000_0000_0000;
array[19569] <= 16'b0000_0000_0000_0000;
array[19570] <= 16'b0000_0000_0000_0000;
array[19571] <= 16'b0000_0000_0000_0000;
array[19572] <= 16'b0000_0000_0000_0000;
array[19573] <= 16'b0000_0000_0000_0000;
array[19574] <= 16'b0000_0000_0000_0000;
array[19575] <= 16'b0000_0000_0000_0000;
array[19576] <= 16'b0000_0000_0000_0000;
array[19577] <= 16'b0000_0000_0000_0000;
array[19578] <= 16'b0000_0000_0000_0000;
array[19579] <= 16'b0000_0000_0000_0000;
array[19580] <= 16'b0000_0000_0000_0000;
array[19581] <= 16'b0000_0000_0000_0000;
array[19582] <= 16'b0000_0000_0000_0000;
array[19583] <= 16'b0000_0000_0000_0000;
array[19584] <= 16'b0000_0000_0000_0000;
array[19585] <= 16'b0000_0000_0000_0000;
array[19586] <= 16'b0000_0000_0000_0000;
array[19587] <= 16'b0000_0000_0000_0000;
array[19588] <= 16'b0000_0000_0000_0000;
array[19589] <= 16'b0000_0000_0000_0000;
array[19590] <= 16'b0000_0000_0000_0000;
array[19591] <= 16'b0000_0000_0000_0000;
array[19592] <= 16'b0000_0000_0000_0000;
array[19593] <= 16'b0000_0000_0000_0000;
array[19594] <= 16'b0000_0000_0000_0000;
array[19595] <= 16'b0000_0000_0000_0000;
array[19596] <= 16'b0000_0000_0000_0000;
array[19597] <= 16'b0000_0000_0000_0000;
array[19598] <= 16'b0000_0000_0000_0000;
array[19599] <= 16'b0000_0000_0000_0000;
array[19600] <= 16'b0000_0000_0000_0000;
array[19601] <= 16'b0000_0000_0000_0000;
array[19602] <= 16'b0000_0000_0000_0000;
array[19603] <= 16'b0000_0000_0000_0000;
array[19604] <= 16'b0000_0000_0000_0000;
array[19605] <= 16'b0000_0000_0000_0000;
array[19606] <= 16'b0000_0000_0000_0000;
array[19607] <= 16'b0000_0000_0000_0000;
array[19608] <= 16'b0000_0000_0000_0000;
array[19609] <= 16'b0000_0000_0000_0000;
array[19610] <= 16'b0000_0000_0000_0000;
array[19611] <= 16'b0000_0000_0000_0000;
array[19612] <= 16'b0000_0000_0000_0000;
array[19613] <= 16'b0000_0000_0000_0000;
array[19614] <= 16'b0000_0000_0000_0000;
array[19615] <= 16'b0000_0000_0000_0000;
array[19616] <= 16'b0000_0000_0000_0000;
array[19617] <= 16'b0000_0000_0000_0000;
array[19618] <= 16'b0000_0000_0000_0000;
array[19619] <= 16'b0000_0000_0000_0000;
array[19620] <= 16'b0000_0000_0000_0000;
array[19621] <= 16'b0000_0000_0000_0000;
array[19622] <= 16'b0000_0000_0000_0000;
array[19623] <= 16'b0000_0000_0000_0000;
array[19624] <= 16'b0000_0000_0000_0000;
array[19625] <= 16'b0000_0000_0000_0000;
array[19626] <= 16'b0000_0000_0000_0000;
array[19627] <= 16'b0000_0000_0000_0000;
array[19628] <= 16'b0000_0000_0000_0000;
array[19629] <= 16'b0000_0000_0000_0000;
array[19630] <= 16'b0000_0000_0000_0000;
array[19631] <= 16'b0000_0000_0000_0000;
array[19632] <= 16'b0000_0000_0000_0000;
array[19633] <= 16'b0000_0000_0000_0000;
array[19634] <= 16'b0000_0000_0000_0000;
array[19635] <= 16'b0000_0000_0000_0000;
array[19636] <= 16'b0000_0000_0000_0000;
array[19637] <= 16'b0000_0000_0000_0000;
array[19638] <= 16'b0000_0000_0000_0000;
array[19639] <= 16'b0000_0000_0000_0000;
array[19640] <= 16'b0000_0000_0000_0000;
array[19641] <= 16'b0000_0000_0000_0000;
array[19642] <= 16'b0000_0000_0000_0000;
array[19643] <= 16'b0000_0000_0000_0000;
array[19644] <= 16'b0000_0000_0000_0000;
array[19645] <= 16'b0000_0000_0000_0000;
array[19646] <= 16'b0000_0000_0000_0000;
array[19647] <= 16'b0000_0000_0000_0000;
array[19648] <= 16'b0000_0000_0000_0000;
array[19649] <= 16'b0000_0000_0000_0000;
array[19650] <= 16'b0000_0000_0000_0000;
array[19651] <= 16'b0000_0000_0000_0000;
array[19652] <= 16'b0000_0000_0000_0000;
array[19653] <= 16'b0000_0000_0000_0000;
array[19654] <= 16'b0000_0000_0000_0000;
array[19655] <= 16'b0000_0000_0000_0000;
array[19656] <= 16'b0000_0000_0000_0000;
array[19657] <= 16'b0000_0000_0000_0000;
array[19658] <= 16'b0000_0000_0000_0000;
array[19659] <= 16'b0000_0000_0000_0000;
array[19660] <= 16'b0000_0000_0000_0000;
array[19661] <= 16'b0000_0000_0000_0000;
array[19662] <= 16'b0000_0000_0000_0000;
array[19663] <= 16'b0000_0000_0000_0000;
array[19664] <= 16'b0000_0000_0000_0000;
array[19665] <= 16'b0000_0000_0000_0000;
array[19666] <= 16'b0000_0000_0000_0000;
array[19667] <= 16'b0000_0000_0000_0000;
array[19668] <= 16'b0000_0000_0000_0000;
array[19669] <= 16'b0000_0000_0000_0000;
array[19670] <= 16'b0000_0000_0000_0000;
array[19671] <= 16'b0000_0000_0000_0000;
array[19672] <= 16'b0000_0000_0000_0000;
array[19673] <= 16'b0000_0000_0000_0000;
array[19674] <= 16'b0000_0000_0000_0000;
array[19675] <= 16'b0000_0000_0000_0000;
array[19676] <= 16'b0000_0000_0000_0000;
array[19677] <= 16'b0000_0000_0000_0000;
array[19678] <= 16'b0000_0000_0000_0000;
array[19679] <= 16'b0000_0000_0000_0000;
array[19680] <= 16'b0000_0000_0000_0000;
array[19681] <= 16'b0000_0000_0000_0000;
array[19682] <= 16'b0000_0000_0000_0000;
array[19683] <= 16'b0000_0000_0000_0000;
array[19684] <= 16'b0000_0000_0000_0000;
array[19685] <= 16'b0000_0000_0000_0000;
array[19686] <= 16'b0000_0000_0000_0000;
array[19687] <= 16'b0000_0000_0000_0000;
array[19688] <= 16'b0000_0000_0000_0000;
array[19689] <= 16'b0000_0000_0000_0000;
array[19690] <= 16'b0000_0000_0000_0000;
array[19691] <= 16'b0000_0000_0000_0000;
array[19692] <= 16'b0000_0000_0000_0000;
array[19693] <= 16'b0000_0000_0000_0000;
array[19694] <= 16'b0000_0000_0000_0000;
array[19695] <= 16'b0000_0000_0000_0000;
array[19696] <= 16'b0000_0000_0000_0000;
array[19697] <= 16'b0000_0000_0000_0000;
array[19698] <= 16'b0000_0000_0000_0000;
array[19699] <= 16'b0000_0000_0000_0000;
array[19700] <= 16'b0000_0000_0000_0000;
array[19701] <= 16'b0000_0000_0000_0000;
array[19702] <= 16'b0000_0000_0000_0000;
array[19703] <= 16'b0000_0000_0000_0000;
array[19704] <= 16'b0000_0000_0000_0000;
array[19705] <= 16'b0000_0000_0000_0000;
array[19706] <= 16'b0000_0000_0000_0000;
array[19707] <= 16'b0000_0000_0000_0000;
array[19708] <= 16'b0000_0000_0000_0000;
array[19709] <= 16'b0000_0000_0000_0000;
array[19710] <= 16'b0000_0000_0000_0000;
array[19711] <= 16'b0000_0000_0000_0000;
array[19712] <= 16'b0000_0000_0000_0000;
array[19713] <= 16'b0000_0000_0000_0000;
array[19714] <= 16'b0000_0000_0000_0000;
array[19715] <= 16'b0000_0000_0000_0000;
array[19716] <= 16'b0000_0000_0000_0000;
array[19717] <= 16'b0000_0000_0000_0000;
array[19718] <= 16'b0000_0000_0000_0000;
array[19719] <= 16'b0000_0000_0000_0000;
array[19720] <= 16'b0000_0000_0000_0000;
array[19721] <= 16'b0000_0000_0000_0000;
array[19722] <= 16'b0000_0000_0000_0000;
array[19723] <= 16'b0000_0000_0000_0000;
array[19724] <= 16'b0000_0000_0000_0000;
array[19725] <= 16'b0000_0000_0000_0000;
array[19726] <= 16'b0000_0000_0000_0000;
array[19727] <= 16'b0000_0000_0000_0000;
array[19728] <= 16'b0000_0000_0000_0000;
array[19729] <= 16'b0000_0000_0000_0000;
array[19730] <= 16'b0000_0000_0000_0000;
array[19731] <= 16'b0000_0000_0000_0000;
array[19732] <= 16'b0000_0000_0000_0000;
array[19733] <= 16'b0000_0000_0000_0000;
array[19734] <= 16'b0000_0000_0000_0000;
array[19735] <= 16'b0000_0000_0000_0000;
array[19736] <= 16'b0000_0000_0000_0000;
array[19737] <= 16'b0000_0000_0000_0000;
array[19738] <= 16'b0000_0000_0000_0000;
array[19739] <= 16'b0000_0000_0000_0000;
array[19740] <= 16'b0000_0000_0000_0000;
array[19741] <= 16'b0000_0000_0000_0000;
array[19742] <= 16'b0000_0000_0000_0000;
array[19743] <= 16'b0000_0000_0000_0000;
array[19744] <= 16'b0000_0000_0000_0000;
array[19745] <= 16'b0000_0000_0000_0000;
array[19746] <= 16'b0000_0000_0000_0000;
array[19747] <= 16'b0000_0000_0000_0000;
array[19748] <= 16'b0000_0000_0000_0000;
array[19749] <= 16'b0000_0000_0000_0000;
array[19750] <= 16'b0000_0000_0000_0000;
array[19751] <= 16'b0000_0000_0000_0000;
array[19752] <= 16'b0000_0000_0000_0000;
array[19753] <= 16'b0000_0000_0000_0000;
array[19754] <= 16'b0000_0000_0000_0000;
array[19755] <= 16'b0000_0000_0000_0000;
array[19756] <= 16'b0000_0000_0000_0000;
array[19757] <= 16'b0000_0000_0000_0000;
array[19758] <= 16'b0000_0000_0000_0000;
array[19759] <= 16'b0000_0000_0000_0000;
array[19760] <= 16'b0000_0000_0000_0000;
array[19761] <= 16'b0000_0000_0000_0000;
array[19762] <= 16'b0000_0000_0000_0000;
array[19763] <= 16'b0000_0000_0000_0000;
array[19764] <= 16'b0000_0000_0000_0000;
array[19765] <= 16'b0000_0000_0000_0000;
array[19766] <= 16'b0000_0000_0000_0000;
array[19767] <= 16'b0000_0000_0000_0000;
array[19768] <= 16'b0000_0000_0000_0000;
array[19769] <= 16'b0000_0000_0000_0000;
array[19770] <= 16'b0000_0000_0000_0000;
array[19771] <= 16'b0000_0000_0000_0000;
array[19772] <= 16'b0000_0000_0000_0000;
array[19773] <= 16'b0000_0000_0000_0000;
array[19774] <= 16'b0000_0000_0000_0000;
array[19775] <= 16'b0000_0000_0000_0000;
array[19776] <= 16'b0000_0000_0000_0000;
array[19777] <= 16'b0000_0000_0000_0000;
array[19778] <= 16'b0000_0000_0000_0000;
array[19779] <= 16'b0000_0000_0000_0000;
array[19780] <= 16'b0000_0000_0000_0000;
array[19781] <= 16'b0000_0000_0000_0000;
array[19782] <= 16'b0000_0000_0000_0000;
array[19783] <= 16'b0000_0000_0000_0000;
array[19784] <= 16'b0000_0000_0000_0000;
array[19785] <= 16'b0000_0000_0000_0000;
array[19786] <= 16'b0000_0000_0000_0000;
array[19787] <= 16'b0000_0000_0000_0000;
array[19788] <= 16'b0000_0000_0000_0000;
array[19789] <= 16'b0000_0000_0000_0000;
array[19790] <= 16'b0000_0000_0000_0000;
array[19791] <= 16'b0000_0000_0000_0000;
array[19792] <= 16'b0000_0000_0000_0000;
array[19793] <= 16'b0000_0000_0000_0000;
array[19794] <= 16'b0000_0000_0000_0000;
array[19795] <= 16'b0000_0000_0000_0000;
array[19796] <= 16'b0000_0000_0000_0000;
array[19797] <= 16'b0000_0000_0000_0000;
array[19798] <= 16'b0000_0000_0000_0000;
array[19799] <= 16'b0000_0000_0000_0000;
array[19800] <= 16'b0000_0000_0000_0000;
array[19801] <= 16'b0000_0000_0000_0000;
array[19802] <= 16'b0000_0000_0000_0000;
array[19803] <= 16'b0000_0000_0000_0000;
array[19804] <= 16'b0000_0000_0000_0000;
array[19805] <= 16'b0000_0000_0000_0000;
array[19806] <= 16'b0000_0000_0000_0000;
array[19807] <= 16'b0000_0000_0000_0000;
array[19808] <= 16'b0000_0000_0000_0000;
array[19809] <= 16'b0000_0000_0000_0000;
array[19810] <= 16'b0000_0000_0000_0000;
array[19811] <= 16'b0000_0000_0000_0000;
array[19812] <= 16'b0000_0000_0000_0000;
array[19813] <= 16'b0000_0000_0000_0000;
array[19814] <= 16'b0000_0000_0000_0000;
array[19815] <= 16'b0000_0000_0000_0000;
array[19816] <= 16'b0000_0000_0000_0000;
array[19817] <= 16'b0000_0000_0000_0000;
array[19818] <= 16'b0000_0000_0000_0000;
array[19819] <= 16'b0000_0000_0000_0000;
array[19820] <= 16'b0000_0000_0000_0000;
array[19821] <= 16'b0000_0000_0000_0000;
array[19822] <= 16'b0000_0000_0000_0000;
array[19823] <= 16'b0000_0000_0000_0000;
array[19824] <= 16'b0000_0000_0000_0000;
array[19825] <= 16'b0000_0000_0000_0000;
array[19826] <= 16'b0000_0000_0000_0000;
array[19827] <= 16'b0000_0000_0000_0000;
array[19828] <= 16'b0000_0000_0000_0000;
array[19829] <= 16'b0000_0000_0000_0000;
array[19830] <= 16'b0000_0000_0000_0000;
array[19831] <= 16'b0000_0000_0000_0000;
array[19832] <= 16'b0000_0000_0000_0000;
array[19833] <= 16'b0000_0000_0000_0000;
array[19834] <= 16'b0000_0000_0000_0000;
array[19835] <= 16'b0000_0000_0000_0000;
array[19836] <= 16'b0000_0000_0000_0000;
array[19837] <= 16'b0000_0000_0000_0000;
array[19838] <= 16'b0000_0000_0000_0000;
array[19839] <= 16'b0000_0000_0000_0000;
array[19840] <= 16'b0000_0000_0000_0000;
array[19841] <= 16'b0000_0000_0000_0000;
array[19842] <= 16'b0000_0000_0000_0000;
array[19843] <= 16'b0000_0000_0000_0000;
array[19844] <= 16'b0000_0000_0000_0000;
array[19845] <= 16'b0000_0000_0000_0000;
array[19846] <= 16'b0000_0000_0000_0000;
array[19847] <= 16'b0000_0000_0000_0000;
array[19848] <= 16'b0000_0000_0000_0000;
array[19849] <= 16'b0000_0000_0000_0000;
array[19850] <= 16'b0000_0000_0000_0000;
array[19851] <= 16'b0000_0000_0000_0000;
array[19852] <= 16'b0000_0000_0000_0000;
array[19853] <= 16'b0000_0000_0000_0000;
array[19854] <= 16'b0000_0000_0000_0000;
array[19855] <= 16'b0000_0000_0000_0000;
array[19856] <= 16'b0000_0000_0000_0000;
array[19857] <= 16'b0000_0000_0000_0000;
array[19858] <= 16'b0000_0000_0000_0000;
array[19859] <= 16'b0000_0000_0000_0000;
array[19860] <= 16'b0000_0000_0000_0000;
array[19861] <= 16'b0000_0000_0000_0000;
array[19862] <= 16'b0000_0000_0000_0000;
array[19863] <= 16'b0000_0000_0000_0000;
array[19864] <= 16'b0000_0000_0000_0000;
array[19865] <= 16'b0000_0000_0000_0000;
array[19866] <= 16'b0000_0000_0000_0000;
array[19867] <= 16'b0000_0000_0000_0000;
array[19868] <= 16'b0000_0000_0000_0000;
array[19869] <= 16'b0000_0000_0000_0000;
array[19870] <= 16'b0000_0000_0000_0000;
array[19871] <= 16'b0000_0000_0000_0000;
array[19872] <= 16'b0000_0000_0000_0000;
array[19873] <= 16'b0000_0000_0000_0000;
array[19874] <= 16'b0000_0000_0000_0000;
array[19875] <= 16'b0000_0000_0000_0000;
array[19876] <= 16'b0000_0000_0000_0000;
array[19877] <= 16'b0000_0000_0000_0000;
array[19878] <= 16'b0000_0000_0000_0000;
array[19879] <= 16'b0000_0000_0000_0000;
array[19880] <= 16'b0000_0000_0000_0000;
array[19881] <= 16'b0000_0000_0000_0000;
array[19882] <= 16'b0000_0000_0000_0000;
array[19883] <= 16'b0000_0000_0000_0000;
array[19884] <= 16'b0000_0000_0000_0000;
array[19885] <= 16'b0000_0000_0000_0000;
array[19886] <= 16'b0000_0000_0000_0000;
array[19887] <= 16'b0000_0000_0000_0000;
array[19888] <= 16'b0000_0000_0000_0000;
array[19889] <= 16'b0000_0000_0000_0000;
array[19890] <= 16'b0000_0000_0000_0000;
array[19891] <= 16'b0000_0000_0000_0000;
array[19892] <= 16'b0000_0000_0000_0000;
array[19893] <= 16'b0000_0000_0000_0000;
array[19894] <= 16'b0000_0000_0000_0000;
array[19895] <= 16'b0000_0000_0000_0000;
array[19896] <= 16'b0000_0000_0000_0000;
array[19897] <= 16'b0000_0000_0000_0000;
array[19898] <= 16'b0000_0000_0000_0000;
array[19899] <= 16'b0000_0000_0000_0000;
array[19900] <= 16'b0000_0000_0000_0000;
array[19901] <= 16'b0000_0000_0000_0000;
array[19902] <= 16'b0000_0000_0000_0000;
array[19903] <= 16'b0000_0000_0000_0000;
array[19904] <= 16'b0000_0000_0000_0000;
array[19905] <= 16'b0000_0000_0000_0000;
array[19906] <= 16'b0000_0000_0000_0000;
array[19907] <= 16'b0000_0000_0000_0000;
array[19908] <= 16'b0000_0000_0000_0000;
array[19909] <= 16'b0000_0000_0000_0000;
array[19910] <= 16'b0000_0000_0000_0000;
array[19911] <= 16'b0000_0000_0000_0000;
array[19912] <= 16'b0000_0000_0000_0000;
array[19913] <= 16'b0000_0000_0000_0000;
array[19914] <= 16'b0000_0000_0000_0000;
array[19915] <= 16'b0000_0000_0000_0000;
array[19916] <= 16'b0000_0000_0000_0000;
array[19917] <= 16'b0000_0000_0000_0000;
array[19918] <= 16'b0000_0000_0000_0000;
array[19919] <= 16'b0000_0000_0000_0000;
array[19920] <= 16'b0000_0000_0000_0000;
array[19921] <= 16'b0000_0000_0000_0000;
array[19922] <= 16'b0000_0000_0000_0000;
array[19923] <= 16'b0000_0000_0000_0000;
array[19924] <= 16'b0000_0000_0000_0000;
array[19925] <= 16'b0000_0000_0000_0000;
array[19926] <= 16'b0000_0000_0000_0000;
array[19927] <= 16'b0000_0000_0000_0000;
array[19928] <= 16'b0000_0000_0000_0000;
array[19929] <= 16'b0000_0000_0000_0000;
array[19930] <= 16'b0000_0000_0000_0000;
array[19931] <= 16'b0000_0000_0000_0000;
array[19932] <= 16'b0000_0000_0000_0000;
array[19933] <= 16'b0000_0000_0000_0000;
array[19934] <= 16'b0000_0000_0000_0000;
array[19935] <= 16'b0000_0000_0000_0000;
array[19936] <= 16'b0000_0000_0000_0000;
array[19937] <= 16'b0000_0000_0000_0000;
array[19938] <= 16'b0000_0000_0000_0000;
array[19939] <= 16'b0000_0000_0000_0000;
array[19940] <= 16'b0000_0000_0000_0000;
array[19941] <= 16'b0000_0000_0000_0000;
array[19942] <= 16'b0000_0000_0000_0000;
array[19943] <= 16'b0000_0000_0000_0000;
array[19944] <= 16'b0000_0000_0000_0000;
array[19945] <= 16'b0000_0000_0000_0000;
array[19946] <= 16'b0000_0000_0000_0000;
array[19947] <= 16'b0000_0000_0000_0000;
array[19948] <= 16'b0000_0000_0000_0000;
array[19949] <= 16'b0000_0000_0000_0000;
array[19950] <= 16'b0000_0000_0000_0000;
array[19951] <= 16'b0000_0000_0000_0000;
array[19952] <= 16'b0000_0000_0000_0000;
array[19953] <= 16'b0000_0000_0000_0000;
array[19954] <= 16'b0000_0000_0000_0000;
array[19955] <= 16'b0000_0000_0000_0000;
array[19956] <= 16'b0000_0000_0000_0000;
array[19957] <= 16'b0000_0000_0000_0000;
array[19958] <= 16'b0000_0000_0000_0000;
array[19959] <= 16'b0000_0000_0000_0000;
array[19960] <= 16'b0000_0000_0000_0000;
array[19961] <= 16'b0000_0000_0000_0000;
array[19962] <= 16'b0000_0000_0000_0000;
array[19963] <= 16'b0000_0000_0000_0000;
array[19964] <= 16'b0000_0000_0000_0000;
array[19965] <= 16'b0000_0000_0000_0000;
array[19966] <= 16'b0000_0000_0000_0000;
array[19967] <= 16'b0000_0000_0000_0000;
array[19968] <= 16'b0000_0000_0000_0000;
array[19969] <= 16'b0000_0000_0000_0000;
array[19970] <= 16'b0000_0000_0000_0000;
array[19971] <= 16'b0000_0000_0000_0000;
array[19972] <= 16'b0000_0000_0000_0000;
array[19973] <= 16'b0000_0000_0000_0000;
array[19974] <= 16'b0000_0000_0000_0000;
array[19975] <= 16'b0000_0000_0000_0000;
array[19976] <= 16'b0000_0000_0000_0000;
array[19977] <= 16'b0000_0000_0000_0000;
array[19978] <= 16'b0000_0000_0000_0000;
array[19979] <= 16'b0000_0000_0000_0000;
array[19980] <= 16'b0000_0000_0000_0000;
array[19981] <= 16'b0000_0000_0000_0000;
array[19982] <= 16'b0000_0000_0000_0000;
array[19983] <= 16'b0000_0000_0000_0000;
array[19984] <= 16'b0000_0000_0000_0000;
array[19985] <= 16'b0000_0000_0000_0000;
array[19986] <= 16'b0000_0000_0000_0000;
array[19987] <= 16'b0000_0000_0000_0000;
array[19988] <= 16'b0000_0000_0000_0000;
array[19989] <= 16'b0000_0000_0000_0000;
array[19990] <= 16'b0000_0000_0000_0000;
array[19991] <= 16'b0000_0000_0000_0000;
array[19992] <= 16'b0000_0000_0000_0000;
array[19993] <= 16'b0000_0000_0000_0000;
array[19994] <= 16'b0000_0000_0000_0000;
array[19995] <= 16'b0000_0000_0000_0000;
array[19996] <= 16'b0000_0000_0000_0000;
array[19997] <= 16'b0000_0000_0000_0000;
array[19998] <= 16'b0000_0000_0000_0000;
array[19999] <= 16'b0000_0000_0000_0000;
array[20000] <= 16'b0000_0000_0000_0000;
array[20001] <= 16'b0000_0000_0000_0000;
array[20002] <= 16'b0000_0000_0000_0000;
array[20003] <= 16'b0000_0000_0000_0000;
array[20004] <= 16'b0000_0000_0000_0000;
array[20005] <= 16'b0000_0000_0000_0000;
array[20006] <= 16'b0000_0000_0000_0000;
array[20007] <= 16'b0000_0000_0000_0000;
array[20008] <= 16'b0000_0000_0000_0000;
array[20009] <= 16'b0000_0000_0000_0000;
array[20010] <= 16'b0000_0000_0000_0000;
array[20011] <= 16'b0000_0000_0000_0000;
array[20012] <= 16'b0000_0000_0000_0000;
array[20013] <= 16'b0000_0000_0000_0000;
array[20014] <= 16'b0000_0000_0000_0000;
array[20015] <= 16'b0000_0000_0000_0000;
array[20016] <= 16'b0000_0000_0000_0000;
array[20017] <= 16'b0000_0000_0000_0000;
array[20018] <= 16'b0000_0000_0000_0000;
array[20019] <= 16'b0000_0000_0000_0000;
array[20020] <= 16'b0000_0000_0000_0000;
array[20021] <= 16'b0000_0000_0000_0000;
array[20022] <= 16'b0000_0000_0000_0000;
array[20023] <= 16'b0000_0000_0000_0000;
array[20024] <= 16'b0000_0000_0000_0000;
array[20025] <= 16'b0000_0000_0000_0000;
array[20026] <= 16'b0000_0000_0000_0000;
array[20027] <= 16'b0000_0000_0000_0000;
array[20028] <= 16'b0000_0000_0000_0000;
array[20029] <= 16'b0000_0000_0000_0000;
array[20030] <= 16'b0000_0000_0000_0000;
array[20031] <= 16'b0000_0000_0000_0000;
array[20032] <= 16'b0000_0000_0000_0000;
array[20033] <= 16'b0000_0000_0000_0000;
array[20034] <= 16'b0000_0000_0000_0000;
array[20035] <= 16'b0000_0000_0000_0000;
array[20036] <= 16'b0000_0000_0000_0000;
array[20037] <= 16'b0000_0000_0000_0000;
array[20038] <= 16'b0000_0000_0000_0000;
array[20039] <= 16'b0000_0000_0000_0000;
array[20040] <= 16'b0000_0000_0000_0000;
array[20041] <= 16'b0000_0000_0000_0000;
array[20042] <= 16'b0000_0000_0000_0000;
array[20043] <= 16'b0000_0000_0000_0000;
array[20044] <= 16'b0000_0000_0000_0000;
array[20045] <= 16'b0000_0000_0000_0000;
array[20046] <= 16'b0000_0000_0000_0000;
array[20047] <= 16'b0000_0000_0000_0000;
array[20048] <= 16'b0000_0000_0000_0000;
array[20049] <= 16'b0000_0000_0000_0000;
array[20050] <= 16'b0000_0000_0000_0000;
array[20051] <= 16'b0000_0000_0000_0000;
array[20052] <= 16'b0000_0000_0000_0000;
array[20053] <= 16'b0000_0000_0000_0000;
array[20054] <= 16'b0000_0000_0000_0000;
array[20055] <= 16'b0000_0000_0000_0000;
array[20056] <= 16'b0000_0000_0000_0000;
array[20057] <= 16'b0000_0000_0000_0000;
array[20058] <= 16'b0000_0000_0000_0000;
array[20059] <= 16'b0000_0000_0000_0000;
array[20060] <= 16'b0000_0000_0000_0000;
array[20061] <= 16'b0000_0000_0000_0000;
array[20062] <= 16'b0000_0000_0000_0000;
array[20063] <= 16'b0000_0000_0000_0000;
array[20064] <= 16'b0000_0000_0000_0000;
array[20065] <= 16'b0000_0000_0000_0000;
array[20066] <= 16'b0000_0000_0000_0000;
array[20067] <= 16'b0000_0000_0000_0000;
array[20068] <= 16'b0000_0000_0000_0000;
array[20069] <= 16'b0000_0000_0000_0000;
array[20070] <= 16'b0000_0000_0000_0000;
array[20071] <= 16'b0000_0000_0000_0000;
array[20072] <= 16'b0000_0000_0000_0000;
array[20073] <= 16'b0000_0000_0000_0000;
array[20074] <= 16'b0000_0000_0000_0000;
array[20075] <= 16'b0000_0000_0000_0000;
array[20076] <= 16'b0000_0000_0000_0000;
array[20077] <= 16'b0000_0000_0000_0000;
array[20078] <= 16'b0000_0000_0000_0000;
array[20079] <= 16'b0000_0000_0000_0000;
array[20080] <= 16'b0000_0000_0000_0000;
array[20081] <= 16'b0000_0000_0000_0000;
array[20082] <= 16'b0000_0000_0000_0000;
array[20083] <= 16'b0000_0000_0000_0000;
array[20084] <= 16'b0000_0000_0000_0000;
array[20085] <= 16'b0000_0000_0000_0000;
array[20086] <= 16'b0000_0000_0000_0000;
array[20087] <= 16'b0000_0000_0000_0000;
array[20088] <= 16'b0000_0000_0000_0000;
array[20089] <= 16'b0000_0000_0000_0000;
array[20090] <= 16'b0000_0000_0000_0000;
array[20091] <= 16'b0000_0000_0000_0000;
array[20092] <= 16'b0000_0000_0000_0000;
array[20093] <= 16'b0000_0000_0000_0000;
array[20094] <= 16'b0000_0000_0000_0000;
array[20095] <= 16'b0000_0000_0000_0000;
array[20096] <= 16'b0000_0000_0000_0000;
array[20097] <= 16'b0000_0000_0000_0000;
array[20098] <= 16'b0000_0000_0000_0000;
array[20099] <= 16'b0000_0000_0000_0000;
array[20100] <= 16'b0000_0000_0000_0000;
array[20101] <= 16'b0000_0000_0000_0000;
array[20102] <= 16'b0000_0000_0000_0000;
array[20103] <= 16'b0000_0000_0000_0000;
array[20104] <= 16'b0000_0000_0000_0000;
array[20105] <= 16'b0000_0000_0000_0000;
array[20106] <= 16'b0000_0000_0000_0000;
array[20107] <= 16'b0000_0000_0000_0000;
array[20108] <= 16'b0000_0000_0000_0000;
array[20109] <= 16'b0000_0000_0000_0000;
array[20110] <= 16'b0000_0000_0000_0000;
array[20111] <= 16'b0000_0000_0000_0000;
array[20112] <= 16'b0000_0000_0000_0000;
array[20113] <= 16'b0000_0000_0000_0000;
array[20114] <= 16'b0000_0000_0000_0000;
array[20115] <= 16'b0000_0000_0000_0000;
array[20116] <= 16'b0000_0000_0000_0000;
array[20117] <= 16'b0000_0000_0000_0000;
array[20118] <= 16'b0000_0000_0000_0000;
array[20119] <= 16'b0000_0000_0000_0000;
array[20120] <= 16'b0000_0000_0000_0000;
array[20121] <= 16'b0000_0000_0000_0000;
array[20122] <= 16'b0000_0000_0000_0000;
array[20123] <= 16'b0000_0000_0000_0000;
array[20124] <= 16'b0000_0000_0000_0000;
array[20125] <= 16'b0000_0000_0000_0000;
array[20126] <= 16'b0000_0000_0000_0000;
array[20127] <= 16'b0000_0000_0000_0000;
array[20128] <= 16'b0000_0000_0000_0000;
array[20129] <= 16'b0000_0000_0000_0000;
array[20130] <= 16'b0000_0000_0000_0000;
array[20131] <= 16'b0000_0000_0000_0000;
array[20132] <= 16'b0000_0000_0000_0000;
array[20133] <= 16'b0000_0000_0000_0000;
array[20134] <= 16'b0000_0000_0000_0000;
array[20135] <= 16'b0000_0000_0000_0000;
array[20136] <= 16'b0000_0000_0000_0000;
array[20137] <= 16'b0000_0000_0000_0000;
array[20138] <= 16'b0000_0000_0000_0000;
array[20139] <= 16'b0000_0000_0000_0000;
array[20140] <= 16'b0000_0000_0000_0000;
array[20141] <= 16'b0000_0000_0000_0000;
array[20142] <= 16'b0000_0000_0000_0000;
array[20143] <= 16'b0000_0000_0000_0000;
array[20144] <= 16'b0000_0000_0000_0000;
array[20145] <= 16'b0000_0000_0000_0000;
array[20146] <= 16'b0000_0000_0000_0000;
array[20147] <= 16'b0000_0000_0000_0000;
array[20148] <= 16'b0000_0000_0000_0000;
array[20149] <= 16'b0000_0000_0000_0000;
array[20150] <= 16'b0000_0000_0000_0000;
array[20151] <= 16'b0000_0000_0000_0000;
array[20152] <= 16'b0000_0000_0000_0000;
array[20153] <= 16'b0000_0000_0000_0000;
array[20154] <= 16'b0000_0000_0000_0000;
array[20155] <= 16'b0000_0000_0000_0000;
array[20156] <= 16'b0000_0000_0000_0000;
array[20157] <= 16'b0000_0000_0000_0000;
array[20158] <= 16'b0000_0000_0000_0000;
array[20159] <= 16'b0000_0000_0000_0000;
array[20160] <= 16'b0000_0000_0000_0000;
array[20161] <= 16'b0000_0000_0000_0000;
array[20162] <= 16'b0000_0000_0000_0000;
array[20163] <= 16'b0000_0000_0000_0000;
array[20164] <= 16'b0000_0000_0000_0000;
array[20165] <= 16'b0000_0000_0000_0000;
array[20166] <= 16'b0000_0000_0000_0000;
array[20167] <= 16'b0000_0000_0000_0000;
array[20168] <= 16'b0000_0000_0000_0000;
array[20169] <= 16'b0000_0000_0000_0000;
array[20170] <= 16'b0000_0000_0000_0000;
array[20171] <= 16'b0000_0000_0000_0000;
array[20172] <= 16'b0000_0000_0000_0000;
array[20173] <= 16'b0000_0000_0000_0000;
array[20174] <= 16'b0000_0000_0000_0000;
array[20175] <= 16'b0000_0000_0000_0000;
array[20176] <= 16'b0000_0000_0000_0000;
array[20177] <= 16'b0000_0000_0000_0000;
array[20178] <= 16'b0000_0000_0000_0000;
array[20179] <= 16'b0000_0000_0000_0000;
array[20180] <= 16'b0000_0000_0000_0000;
array[20181] <= 16'b0000_0000_0000_0000;
array[20182] <= 16'b0000_0000_0000_0000;
array[20183] <= 16'b0000_0000_0000_0000;
array[20184] <= 16'b0000_0000_0000_0000;
array[20185] <= 16'b0000_0000_0000_0000;
array[20186] <= 16'b0000_0000_0000_0000;
array[20187] <= 16'b0000_0000_0000_0000;
array[20188] <= 16'b0000_0000_0000_0000;
array[20189] <= 16'b0000_0000_0000_0000;
array[20190] <= 16'b0000_0000_0000_0000;
array[20191] <= 16'b0000_0000_0000_0000;
array[20192] <= 16'b0000_0000_0000_0000;
array[20193] <= 16'b0000_0000_0000_0000;
array[20194] <= 16'b0000_0000_0000_0000;
array[20195] <= 16'b0000_0000_0000_0000;
array[20196] <= 16'b0000_0000_0000_0000;
array[20197] <= 16'b0000_0000_0000_0000;
array[20198] <= 16'b0000_0000_0000_0000;
array[20199] <= 16'b0000_0000_0000_0000;
array[20200] <= 16'b0000_0000_0000_0000;
array[20201] <= 16'b0000_0000_0000_0000;
array[20202] <= 16'b0000_0000_0000_0000;
array[20203] <= 16'b0000_0000_0000_0000;
array[20204] <= 16'b0000_0000_0000_0000;
array[20205] <= 16'b0000_0000_0000_0000;
array[20206] <= 16'b0000_0000_0000_0000;
array[20207] <= 16'b0000_0000_0000_0000;
array[20208] <= 16'b0000_0000_0000_0000;
array[20209] <= 16'b0000_0000_0000_0000;
array[20210] <= 16'b0000_0000_0000_0000;
array[20211] <= 16'b0000_0000_0000_0000;
array[20212] <= 16'b0000_0000_0000_0000;
array[20213] <= 16'b0000_0000_0000_0000;
array[20214] <= 16'b0000_0000_0000_0000;
array[20215] <= 16'b0000_0000_0000_0000;
array[20216] <= 16'b0000_0000_0000_0000;
array[20217] <= 16'b0000_0000_0000_0000;
array[20218] <= 16'b0000_0000_0000_0000;
array[20219] <= 16'b0000_0000_0000_0000;
array[20220] <= 16'b0000_0000_0000_0000;
array[20221] <= 16'b0000_0000_0000_0000;
array[20222] <= 16'b0000_0000_0000_0000;
array[20223] <= 16'b0000_0000_0000_0000;
array[20224] <= 16'b0000_0000_0000_0000;
array[20225] <= 16'b0000_0000_0000_0000;
array[20226] <= 16'b0000_0000_0000_0000;
array[20227] <= 16'b0000_0000_0000_0000;
array[20228] <= 16'b0000_0000_0000_0000;
array[20229] <= 16'b0000_0000_0000_0000;
array[20230] <= 16'b0000_0000_0000_0000;
array[20231] <= 16'b0000_0000_0000_0000;
array[20232] <= 16'b0000_0000_0000_0000;
array[20233] <= 16'b0000_0000_0000_0000;
array[20234] <= 16'b0000_0000_0000_0000;
array[20235] <= 16'b0000_0000_0000_0000;
array[20236] <= 16'b0000_0000_0000_0000;
array[20237] <= 16'b0000_0000_0000_0000;
array[20238] <= 16'b0000_0000_0000_0000;
array[20239] <= 16'b0000_0000_0000_0000;
array[20240] <= 16'b0000_0000_0000_0000;
array[20241] <= 16'b0000_0000_0000_0000;
array[20242] <= 16'b0000_0000_0000_0000;
array[20243] <= 16'b0000_0000_0000_0000;
array[20244] <= 16'b0000_0000_0000_0000;
array[20245] <= 16'b0000_0000_0000_0000;
array[20246] <= 16'b0000_0000_0000_0000;
array[20247] <= 16'b0000_0000_0000_0000;
array[20248] <= 16'b0000_0000_0000_0000;
array[20249] <= 16'b0000_0000_0000_0000;
array[20250] <= 16'b0000_0000_0000_0000;
array[20251] <= 16'b0000_0000_0000_0000;
array[20252] <= 16'b0000_0000_0000_0000;
array[20253] <= 16'b0000_0000_0000_0000;
array[20254] <= 16'b0000_0000_0000_0000;
array[20255] <= 16'b0000_0000_0000_0000;
array[20256] <= 16'b0000_0000_0000_0000;
array[20257] <= 16'b0000_0000_0000_0000;
array[20258] <= 16'b0000_0000_0000_0000;
array[20259] <= 16'b0000_0000_0000_0000;
array[20260] <= 16'b0000_0000_0000_0000;
array[20261] <= 16'b0000_0000_0000_0000;
array[20262] <= 16'b0000_0000_0000_0000;
array[20263] <= 16'b0000_0000_0000_0000;
array[20264] <= 16'b0000_0000_0000_0000;
array[20265] <= 16'b0000_0000_0000_0000;
array[20266] <= 16'b0000_0000_0000_0000;
array[20267] <= 16'b0000_0000_0000_0000;
array[20268] <= 16'b0000_0000_0000_0000;
array[20269] <= 16'b0000_0000_0000_0000;
array[20270] <= 16'b0000_0000_0000_0000;
array[20271] <= 16'b0000_0000_0000_0000;
array[20272] <= 16'b0000_0000_0000_0000;
array[20273] <= 16'b0000_0000_0000_0000;
array[20274] <= 16'b0000_0000_0000_0000;
array[20275] <= 16'b0000_0000_0000_0000;
array[20276] <= 16'b0000_0000_0000_0000;
array[20277] <= 16'b0000_0000_0000_0000;
array[20278] <= 16'b0000_0000_0000_0000;
array[20279] <= 16'b0000_0000_0000_0000;
array[20280] <= 16'b0000_0000_0000_0000;
array[20281] <= 16'b0000_0000_0000_0000;
array[20282] <= 16'b0000_0000_0000_0000;
array[20283] <= 16'b0000_0000_0000_0000;
array[20284] <= 16'b0000_0000_0000_0000;
array[20285] <= 16'b0000_0000_0000_0000;
array[20286] <= 16'b0000_0000_0000_0000;
array[20287] <= 16'b0000_0000_0000_0000;
array[20288] <= 16'b0000_0000_0000_0000;
array[20289] <= 16'b0000_0000_0000_0000;
array[20290] <= 16'b0000_0000_0000_0000;
array[20291] <= 16'b0000_0000_0000_0000;
array[20292] <= 16'b0000_0000_0000_0000;
array[20293] <= 16'b0000_0000_0000_0000;
array[20294] <= 16'b0000_0000_0000_0000;
array[20295] <= 16'b0000_0000_0000_0000;
array[20296] <= 16'b0000_0000_0000_0000;
array[20297] <= 16'b0000_0000_0000_0000;
array[20298] <= 16'b0000_0000_0000_0000;
array[20299] <= 16'b0000_0000_0000_0000;
array[20300] <= 16'b0000_0000_0000_0000;
array[20301] <= 16'b0000_0000_0000_0000;
array[20302] <= 16'b0000_0000_0000_0000;
array[20303] <= 16'b0000_0000_0000_0000;
array[20304] <= 16'b0000_0000_0000_0000;
array[20305] <= 16'b0000_0000_0000_0000;
array[20306] <= 16'b0000_0000_0000_0000;
array[20307] <= 16'b0000_0000_0000_0000;
array[20308] <= 16'b0000_0000_0000_0000;
array[20309] <= 16'b0000_0000_0000_0000;
array[20310] <= 16'b0000_0000_0000_0000;
array[20311] <= 16'b0000_0000_0000_0000;
array[20312] <= 16'b0000_0000_0000_0000;
array[20313] <= 16'b0000_0000_0000_0000;
array[20314] <= 16'b0000_0000_0000_0000;
array[20315] <= 16'b0000_0000_0000_0000;
array[20316] <= 16'b0000_0000_0000_0000;
array[20317] <= 16'b0000_0000_0000_0000;
array[20318] <= 16'b0000_0000_0000_0000;
array[20319] <= 16'b0000_0000_0000_0000;
array[20320] <= 16'b0000_0000_0000_0000;
array[20321] <= 16'b0000_0000_0000_0000;
array[20322] <= 16'b0000_0000_0000_0000;
array[20323] <= 16'b0000_0000_0000_0000;
array[20324] <= 16'b0000_0000_0000_0000;
array[20325] <= 16'b0000_0000_0000_0000;
array[20326] <= 16'b0000_0000_0000_0000;
array[20327] <= 16'b0000_0000_0000_0000;
array[20328] <= 16'b0000_0000_0000_0000;
array[20329] <= 16'b0000_0000_0000_0000;
array[20330] <= 16'b0000_0000_0000_0000;
array[20331] <= 16'b0000_0000_0000_0000;
array[20332] <= 16'b0000_0000_0000_0000;
array[20333] <= 16'b0000_0000_0000_0000;
array[20334] <= 16'b0000_0000_0000_0000;
array[20335] <= 16'b0000_0000_0000_0000;
array[20336] <= 16'b0000_0000_0000_0000;
array[20337] <= 16'b0000_0000_0000_0000;
array[20338] <= 16'b0000_0000_0000_0000;
array[20339] <= 16'b0000_0000_0000_0000;
array[20340] <= 16'b0000_0000_0000_0000;
array[20341] <= 16'b0000_0000_0000_0000;
array[20342] <= 16'b0000_0000_0000_0000;
array[20343] <= 16'b0000_0000_0000_0000;
array[20344] <= 16'b0000_0000_0000_0000;
array[20345] <= 16'b0000_0000_0000_0000;
array[20346] <= 16'b0000_0000_0000_0000;
array[20347] <= 16'b0000_0000_0000_0000;
array[20348] <= 16'b0000_0000_0000_0000;
array[20349] <= 16'b0000_0000_0000_0000;
array[20350] <= 16'b0000_0000_0000_0000;
array[20351] <= 16'b0000_0000_0000_0000;
array[20352] <= 16'b0000_0000_0000_0000;
array[20353] <= 16'b0000_0000_0000_0000;
array[20354] <= 16'b0000_0000_0000_0000;
array[20355] <= 16'b0000_0000_0000_0000;
array[20356] <= 16'b0000_0000_0000_0000;
array[20357] <= 16'b0000_0000_0000_0000;
array[20358] <= 16'b0000_0000_0000_0000;
array[20359] <= 16'b0000_0000_0000_0000;
array[20360] <= 16'b0000_0000_0000_0000;
array[20361] <= 16'b0000_0000_0000_0000;
array[20362] <= 16'b0000_0000_0000_0000;
array[20363] <= 16'b0000_0000_0000_0000;
array[20364] <= 16'b0000_0000_0000_0000;
array[20365] <= 16'b0000_0000_0000_0000;
array[20366] <= 16'b0000_0000_0000_0000;
array[20367] <= 16'b0000_0000_0000_0000;
array[20368] <= 16'b0000_0000_0000_0000;
array[20369] <= 16'b0000_0000_0000_0000;
array[20370] <= 16'b0000_0000_0000_0000;
array[20371] <= 16'b0000_0000_0000_0000;
array[20372] <= 16'b0000_0000_0000_0000;
array[20373] <= 16'b0000_0000_0000_0000;
array[20374] <= 16'b0000_0000_0000_0000;
array[20375] <= 16'b0000_0000_0000_0000;
array[20376] <= 16'b0000_0000_0000_0000;
array[20377] <= 16'b0000_0000_0000_0000;
array[20378] <= 16'b0000_0000_0000_0000;
array[20379] <= 16'b0000_0000_0000_0000;
array[20380] <= 16'b0000_0000_0000_0000;
array[20381] <= 16'b0000_0000_0000_0000;
array[20382] <= 16'b0000_0000_0000_0000;
array[20383] <= 16'b0000_0000_0000_0000;
array[20384] <= 16'b0000_0000_0000_0000;
array[20385] <= 16'b0000_0000_0000_0000;
array[20386] <= 16'b0000_0000_0000_0000;
array[20387] <= 16'b0000_0000_0000_0000;
array[20388] <= 16'b0000_0000_0000_0000;
array[20389] <= 16'b0000_0000_0000_0000;
array[20390] <= 16'b0000_0000_0000_0000;
array[20391] <= 16'b0000_0000_0000_0000;
array[20392] <= 16'b0000_0000_0000_0000;
array[20393] <= 16'b0000_0000_0000_0000;
array[20394] <= 16'b0000_0000_0000_0000;
array[20395] <= 16'b0000_0000_0000_0000;
array[20396] <= 16'b0000_0000_0000_0000;
array[20397] <= 16'b0000_0000_0000_0000;
array[20398] <= 16'b0000_0000_0000_0000;
array[20399] <= 16'b0000_0000_0000_0000;
array[20400] <= 16'b0000_0000_0000_0000;
array[20401] <= 16'b0000_0000_0000_0000;
array[20402] <= 16'b0000_0000_0000_0000;
array[20403] <= 16'b0000_0000_0000_0000;
array[20404] <= 16'b0000_0000_0000_0000;
array[20405] <= 16'b0000_0000_0000_0000;
array[20406] <= 16'b0000_0000_0000_0000;
array[20407] <= 16'b0000_0000_0000_0000;
array[20408] <= 16'b0000_0000_0000_0000;
array[20409] <= 16'b0000_0000_0000_0000;
array[20410] <= 16'b0000_0000_0000_0000;
array[20411] <= 16'b0000_0000_0000_0000;
array[20412] <= 16'b0000_0000_0000_0000;
array[20413] <= 16'b0000_0000_0000_0000;
array[20414] <= 16'b0000_0000_0000_0000;
array[20415] <= 16'b0000_0000_0000_0000;
array[20416] <= 16'b0000_0000_0000_0000;
array[20417] <= 16'b0000_0000_0000_0000;
array[20418] <= 16'b0000_0000_0000_0000;
array[20419] <= 16'b0000_0000_0000_0000;
array[20420] <= 16'b0000_0000_0000_0000;
array[20421] <= 16'b0000_0000_0000_0000;
array[20422] <= 16'b0000_0000_0000_0000;
array[20423] <= 16'b0000_0000_0000_0000;
array[20424] <= 16'b0000_0000_0000_0000;
array[20425] <= 16'b0000_0000_0000_0000;
array[20426] <= 16'b0000_0000_0000_0000;
array[20427] <= 16'b0000_0000_0000_0000;
array[20428] <= 16'b0000_0000_0000_0000;
array[20429] <= 16'b0000_0000_0000_0000;
array[20430] <= 16'b0000_0000_0000_0000;
array[20431] <= 16'b0000_0000_0000_0000;
array[20432] <= 16'b0000_0000_0000_0000;
array[20433] <= 16'b0000_0000_0000_0000;
array[20434] <= 16'b0000_0000_0000_0000;
array[20435] <= 16'b0000_0000_0000_0000;
array[20436] <= 16'b0000_0000_0000_0000;
array[20437] <= 16'b0000_0000_0000_0000;
array[20438] <= 16'b0000_0000_0000_0000;
array[20439] <= 16'b0000_0000_0000_0000;
array[20440] <= 16'b0000_0000_0000_0000;
array[20441] <= 16'b0000_0000_0000_0000;
array[20442] <= 16'b0000_0000_0000_0000;
array[20443] <= 16'b0000_0000_0000_0000;
array[20444] <= 16'b0000_0000_0000_0000;
array[20445] <= 16'b0000_0000_0000_0000;
array[20446] <= 16'b0000_0000_0000_0000;
array[20447] <= 16'b0000_0000_0000_0000;
array[20448] <= 16'b0000_0000_0000_0000;
array[20449] <= 16'b0000_0000_0000_0000;
array[20450] <= 16'b0000_0000_0000_0000;
array[20451] <= 16'b0000_0000_0000_0000;
array[20452] <= 16'b0000_0000_0000_0000;
array[20453] <= 16'b0000_0000_0000_0000;
array[20454] <= 16'b0000_0000_0000_0000;
array[20455] <= 16'b0000_0000_0000_0000;
array[20456] <= 16'b0000_0000_0000_0000;
array[20457] <= 16'b0000_0000_0000_0000;
array[20458] <= 16'b0000_0000_0000_0000;
array[20459] <= 16'b0000_0000_0000_0000;
array[20460] <= 16'b0000_0000_0000_0000;
array[20461] <= 16'b0000_0000_0000_0000;
array[20462] <= 16'b0000_0000_0000_0000;
array[20463] <= 16'b0000_0000_0000_0000;
array[20464] <= 16'b0000_0000_0000_0000;
array[20465] <= 16'b0000_0000_0000_0000;
array[20466] <= 16'b0000_0000_0000_0000;
array[20467] <= 16'b0000_0000_0000_0000;
array[20468] <= 16'b0000_0000_0000_0000;
array[20469] <= 16'b0000_0000_0000_0000;
array[20470] <= 16'b0000_0000_0000_0000;
array[20471] <= 16'b0000_0000_0000_0000;
array[20472] <= 16'b0000_0000_0000_0000;
array[20473] <= 16'b0000_0000_0000_0000;
array[20474] <= 16'b0000_0000_0000_0000;
array[20475] <= 16'b0000_0000_0000_0000;
array[20476] <= 16'b0000_0000_0000_0000;
array[20477] <= 16'b0000_0000_0000_0000;
array[20478] <= 16'b0000_0000_0000_0000;
array[20479] <= 16'b0000_0000_0000_0000;
array[20480] <= 16'b0000_0000_0000_0000;
array[20481] <= 16'b0000_0000_0000_0000;
array[20482] <= 16'b0000_0000_0000_0000;
array[20483] <= 16'b0000_0000_0000_0000;
array[20484] <= 16'b0000_0000_0000_0000;
array[20485] <= 16'b0000_0000_0000_0000;
array[20486] <= 16'b0000_0000_0000_0000;
array[20487] <= 16'b0000_0000_0000_0000;
array[20488] <= 16'b0000_0000_0000_0000;
array[20489] <= 16'b0000_0000_0000_0000;
array[20490] <= 16'b0000_0000_0000_0000;
array[20491] <= 16'b0000_0000_0000_0000;
array[20492] <= 16'b0000_0000_0000_0000;
array[20493] <= 16'b0000_0000_0000_0000;
array[20494] <= 16'b0000_0000_0000_0000;
array[20495] <= 16'b0000_0000_0000_0000;
array[20496] <= 16'b0000_0000_0000_0000;
array[20497] <= 16'b0000_0000_0000_0000;
array[20498] <= 16'b0000_0000_0000_0000;
array[20499] <= 16'b0000_0000_0000_0000;
array[20500] <= 16'b0000_0000_0000_0000;
array[20501] <= 16'b0000_0000_0000_0000;
array[20502] <= 16'b0000_0000_0000_0000;
array[20503] <= 16'b0000_0000_0000_0000;
array[20504] <= 16'b0000_0000_0000_0000;
array[20505] <= 16'b0000_0000_0000_0000;
array[20506] <= 16'b0000_0000_0000_0000;
array[20507] <= 16'b0000_0000_0000_0000;
array[20508] <= 16'b0000_0000_0000_0000;
array[20509] <= 16'b0000_0000_0000_0000;
array[20510] <= 16'b0000_0000_0000_0000;
array[20511] <= 16'b0000_0000_0000_0000;
array[20512] <= 16'b0000_0000_0000_0000;
array[20513] <= 16'b0000_0000_0000_0000;
array[20514] <= 16'b0000_0000_0000_0000;
array[20515] <= 16'b0000_0000_0000_0000;
array[20516] <= 16'b0000_0000_0000_0000;
array[20517] <= 16'b0000_0000_0000_0000;
array[20518] <= 16'b0000_0000_0000_0000;
array[20519] <= 16'b0000_0000_0000_0000;
array[20520] <= 16'b0000_0000_0000_0000;
array[20521] <= 16'b0000_0000_0000_0000;
array[20522] <= 16'b0000_0000_0000_0000;
array[20523] <= 16'b0000_0000_0000_0000;
array[20524] <= 16'b0000_0000_0000_0000;
array[20525] <= 16'b0000_0000_0000_0000;
array[20526] <= 16'b0000_0000_0000_0000;
array[20527] <= 16'b0000_0000_0000_0000;
array[20528] <= 16'b0000_0000_0000_0000;
array[20529] <= 16'b0000_0000_0000_0000;
array[20530] <= 16'b0000_0000_0000_0000;
array[20531] <= 16'b0000_0000_0000_0000;
array[20532] <= 16'b0000_0000_0000_0000;
array[20533] <= 16'b0000_0000_0000_0000;
array[20534] <= 16'b0000_0000_0000_0000;
array[20535] <= 16'b0000_0000_0000_0000;
array[20536] <= 16'b0000_0000_0000_0000;
array[20537] <= 16'b0000_0000_0000_0000;
array[20538] <= 16'b0000_0000_0000_0000;
array[20539] <= 16'b0000_0000_0000_0000;
array[20540] <= 16'b0000_0000_0000_0000;
array[20541] <= 16'b0000_0000_0000_0000;
array[20542] <= 16'b0000_0000_0000_0000;
array[20543] <= 16'b0000_0000_0000_0000;
array[20544] <= 16'b0000_0000_0000_0000;
array[20545] <= 16'b0000_0000_0000_0000;
array[20546] <= 16'b0000_0000_0000_0000;
array[20547] <= 16'b0000_0000_0000_0000;
array[20548] <= 16'b0000_0000_0000_0000;
array[20549] <= 16'b0000_0000_0000_0000;
array[20550] <= 16'b0000_0000_0000_0000;
array[20551] <= 16'b0000_0000_0000_0000;
array[20552] <= 16'b0000_0000_0000_0000;
array[20553] <= 16'b0000_0000_0000_0000;
array[20554] <= 16'b0000_0000_0000_0000;
array[20555] <= 16'b0000_0000_0000_0000;
array[20556] <= 16'b0000_0000_0000_0000;
array[20557] <= 16'b0000_0000_0000_0000;
array[20558] <= 16'b0000_0000_0000_0000;
array[20559] <= 16'b0000_0000_0000_0000;
array[20560] <= 16'b0000_0000_0000_0000;
array[20561] <= 16'b0000_0000_0000_0000;
array[20562] <= 16'b0000_0000_0000_0000;
array[20563] <= 16'b0000_0000_0000_0000;
array[20564] <= 16'b0000_0000_0000_0000;
array[20565] <= 16'b0000_0000_0000_0000;
array[20566] <= 16'b0000_0000_0000_0000;
array[20567] <= 16'b0000_0000_0000_0000;
array[20568] <= 16'b0000_0000_0000_0000;
array[20569] <= 16'b0000_0000_0000_0000;
array[20570] <= 16'b0000_0000_0000_0000;
array[20571] <= 16'b0000_0000_0000_0000;
array[20572] <= 16'b0000_0000_0000_0000;
array[20573] <= 16'b0000_0000_0000_0000;
array[20574] <= 16'b0000_0000_0000_0000;
array[20575] <= 16'b0000_0000_0000_0000;
array[20576] <= 16'b0000_0000_0000_0000;
array[20577] <= 16'b0000_0000_0000_0000;
array[20578] <= 16'b0000_0000_0000_0000;
array[20579] <= 16'b0000_0000_0000_0000;
array[20580] <= 16'b0000_0000_0000_0000;
array[20581] <= 16'b0000_0000_0000_0000;
array[20582] <= 16'b0000_0000_0000_0000;
array[20583] <= 16'b0000_0000_0000_0000;
array[20584] <= 16'b0000_0000_0000_0000;
array[20585] <= 16'b0000_0000_0000_0000;
array[20586] <= 16'b0000_0000_0000_0000;
array[20587] <= 16'b0000_0000_0000_0000;
array[20588] <= 16'b0000_0000_0000_0000;
array[20589] <= 16'b0000_0000_0000_0000;
array[20590] <= 16'b0000_0000_0000_0000;
array[20591] <= 16'b0000_0000_0000_0000;
array[20592] <= 16'b0000_0000_0000_0000;
array[20593] <= 16'b0000_0000_0000_0000;
array[20594] <= 16'b0000_0000_0000_0000;
array[20595] <= 16'b0000_0000_0000_0000;
array[20596] <= 16'b0000_0000_0000_0000;
array[20597] <= 16'b0000_0000_0000_0000;
array[20598] <= 16'b0000_0000_0000_0000;
array[20599] <= 16'b0000_0000_0000_0000;
array[20600] <= 16'b0000_0000_0000_0000;
array[20601] <= 16'b0000_0000_0000_0000;
array[20602] <= 16'b0000_0000_0000_0000;
array[20603] <= 16'b0000_0000_0000_0000;
array[20604] <= 16'b0000_0000_0000_0000;
array[20605] <= 16'b0000_0000_0000_0000;
array[20606] <= 16'b0000_0000_0000_0000;
array[20607] <= 16'b0000_0000_0000_0000;
array[20608] <= 16'b0000_0000_0000_0000;
array[20609] <= 16'b0000_0000_0000_0000;
array[20610] <= 16'b0000_0000_0000_0000;
array[20611] <= 16'b0000_0000_0000_0000;
array[20612] <= 16'b0000_0000_0000_0000;
array[20613] <= 16'b0000_0000_0000_0000;
array[20614] <= 16'b0000_0000_0000_0000;
array[20615] <= 16'b0000_0000_0000_0000;
array[20616] <= 16'b0000_0000_0000_0000;
array[20617] <= 16'b0000_0000_0000_0000;
array[20618] <= 16'b0000_0000_0000_0000;
array[20619] <= 16'b0000_0000_0000_0000;
array[20620] <= 16'b0000_0000_0000_0000;
array[20621] <= 16'b0000_0000_0000_0000;
array[20622] <= 16'b0000_0000_0000_0000;
array[20623] <= 16'b0000_0000_0000_0000;
array[20624] <= 16'b0000_0000_0000_0000;
array[20625] <= 16'b0000_0000_0000_0000;
array[20626] <= 16'b0000_0000_0000_0000;
array[20627] <= 16'b0000_0000_0000_0000;
array[20628] <= 16'b0000_0000_0000_0000;
array[20629] <= 16'b0000_0000_0000_0000;
array[20630] <= 16'b0000_0000_0000_0000;
array[20631] <= 16'b0000_0000_0000_0000;
array[20632] <= 16'b0000_0000_0000_0000;
array[20633] <= 16'b0000_0000_0000_0000;
array[20634] <= 16'b0000_0000_0000_0000;
array[20635] <= 16'b0000_0000_0000_0000;
array[20636] <= 16'b0000_0000_0000_0000;
array[20637] <= 16'b0000_0000_0000_0000;
array[20638] <= 16'b0000_0000_0000_0000;
array[20639] <= 16'b0000_0000_0000_0000;
array[20640] <= 16'b0000_0000_0000_0000;
array[20641] <= 16'b0000_0000_0000_0000;
array[20642] <= 16'b0000_0000_0000_0000;
array[20643] <= 16'b0000_0000_0000_0000;
array[20644] <= 16'b0000_0000_0000_0000;
array[20645] <= 16'b0000_0000_0000_0000;
array[20646] <= 16'b0000_0000_0000_0000;
array[20647] <= 16'b0000_0000_0000_0000;
array[20648] <= 16'b0000_0000_0000_0000;
array[20649] <= 16'b0000_0000_0000_0000;
array[20650] <= 16'b0000_0000_0000_0000;
array[20651] <= 16'b0000_0000_0000_0000;
array[20652] <= 16'b0000_0000_0000_0000;
array[20653] <= 16'b0000_0000_0000_0000;
array[20654] <= 16'b0000_0000_0000_0000;
array[20655] <= 16'b0000_0000_0000_0000;
array[20656] <= 16'b0000_0000_0000_0000;
array[20657] <= 16'b0000_0000_0000_0000;
array[20658] <= 16'b0000_0000_0000_0000;
array[20659] <= 16'b0000_0000_0000_0000;
array[20660] <= 16'b0000_0000_0000_0000;
array[20661] <= 16'b0000_0000_0000_0000;
array[20662] <= 16'b0000_0000_0000_0000;
array[20663] <= 16'b0000_0000_0000_0000;
array[20664] <= 16'b0000_0000_0000_0000;
array[20665] <= 16'b0000_0000_0000_0000;
array[20666] <= 16'b0000_0000_0000_0000;
array[20667] <= 16'b0000_0000_0000_0000;
array[20668] <= 16'b0000_0000_0000_0000;
array[20669] <= 16'b0000_0000_0000_0000;
array[20670] <= 16'b0000_0000_0000_0000;
array[20671] <= 16'b0000_0000_0000_0000;
array[20672] <= 16'b0000_0000_0000_0000;
array[20673] <= 16'b0000_0000_0000_0000;
array[20674] <= 16'b0000_0000_0000_0000;
array[20675] <= 16'b0000_0000_0000_0000;
array[20676] <= 16'b0000_0000_0000_0000;
array[20677] <= 16'b0000_0000_0000_0000;
array[20678] <= 16'b0000_0000_0000_0000;
array[20679] <= 16'b0000_0000_0000_0000;
array[20680] <= 16'b0000_0000_0000_0000;
array[20681] <= 16'b0000_0000_0000_0000;
array[20682] <= 16'b0000_0000_0000_0000;
array[20683] <= 16'b0000_0000_0000_0000;
array[20684] <= 16'b0000_0000_0000_0000;
array[20685] <= 16'b0000_0000_0000_0000;
array[20686] <= 16'b0000_0000_0000_0000;
array[20687] <= 16'b0000_0000_0000_0000;
array[20688] <= 16'b0000_0000_0000_0000;
array[20689] <= 16'b0000_0000_0000_0000;
array[20690] <= 16'b0000_0000_0000_0000;
array[20691] <= 16'b0000_0000_0000_0000;
array[20692] <= 16'b0000_0000_0000_0000;
array[20693] <= 16'b0000_0000_0000_0000;
array[20694] <= 16'b0000_0000_0000_0000;
array[20695] <= 16'b0000_0000_0000_0000;
array[20696] <= 16'b0000_0000_0000_0000;
array[20697] <= 16'b0000_0000_0000_0000;
array[20698] <= 16'b0000_0000_0000_0000;
array[20699] <= 16'b0000_0000_0000_0000;
array[20700] <= 16'b0000_0000_0000_0000;
array[20701] <= 16'b0000_0000_0000_0000;
array[20702] <= 16'b0000_0000_0000_0000;
array[20703] <= 16'b0000_0000_0000_0000;
array[20704] <= 16'b0000_0000_0000_0000;
array[20705] <= 16'b0000_0000_0000_0000;
array[20706] <= 16'b0000_0000_0000_0000;
array[20707] <= 16'b0000_0000_0000_0000;
array[20708] <= 16'b0000_0000_0000_0000;
array[20709] <= 16'b0000_0000_0000_0000;
array[20710] <= 16'b0000_0000_0000_0000;
array[20711] <= 16'b0000_0000_0000_0000;
array[20712] <= 16'b0000_0000_0000_0000;
array[20713] <= 16'b0000_0000_0000_0000;
array[20714] <= 16'b0000_0000_0000_0000;
array[20715] <= 16'b0000_0000_0000_0000;
array[20716] <= 16'b0000_0000_0000_0000;
array[20717] <= 16'b0000_0000_0000_0000;
array[20718] <= 16'b0000_0000_0000_0000;
array[20719] <= 16'b0000_0000_0000_0000;
array[20720] <= 16'b0000_0000_0000_0000;
array[20721] <= 16'b0000_0000_0000_0000;
array[20722] <= 16'b0000_0000_0000_0000;
array[20723] <= 16'b0000_0000_0000_0000;
array[20724] <= 16'b0000_0000_0000_0000;
array[20725] <= 16'b0000_0000_0000_0000;
array[20726] <= 16'b0000_0000_0000_0000;
array[20727] <= 16'b0000_0000_0000_0000;
array[20728] <= 16'b0000_0000_0000_0000;
array[20729] <= 16'b0000_0000_0000_0000;
array[20730] <= 16'b0000_0000_0000_0000;
array[20731] <= 16'b0000_0000_0000_0000;
array[20732] <= 16'b0000_0000_0000_0000;
array[20733] <= 16'b0000_0000_0000_0000;
array[20734] <= 16'b0000_0000_0000_0000;
array[20735] <= 16'b0000_0000_0000_0000;
array[20736] <= 16'b0000_0000_0000_0000;
array[20737] <= 16'b0000_0000_0000_0000;
array[20738] <= 16'b0000_0000_0000_0000;
array[20739] <= 16'b0000_0000_0000_0000;
array[20740] <= 16'b0000_0000_0000_0000;
array[20741] <= 16'b0000_0000_0000_0000;
array[20742] <= 16'b0000_0000_0000_0000;
array[20743] <= 16'b0000_0000_0000_0000;
array[20744] <= 16'b0000_0000_0000_0000;
array[20745] <= 16'b0000_0000_0000_0000;
array[20746] <= 16'b0000_0000_0000_0000;
array[20747] <= 16'b0000_0000_0000_0000;
array[20748] <= 16'b0000_0000_0000_0000;
array[20749] <= 16'b0000_0000_0000_0000;
array[20750] <= 16'b0000_0000_0000_0000;
array[20751] <= 16'b0000_0000_0000_0000;
array[20752] <= 16'b0000_0000_0000_0000;
array[20753] <= 16'b0000_0000_0000_0000;
array[20754] <= 16'b0000_0000_0000_0000;
array[20755] <= 16'b0000_0000_0000_0000;
array[20756] <= 16'b0000_0000_0000_0000;
array[20757] <= 16'b0000_0000_0000_0000;
array[20758] <= 16'b0000_0000_0000_0000;
array[20759] <= 16'b0000_0000_0000_0000;
array[20760] <= 16'b0000_0000_0000_0000;
array[20761] <= 16'b0000_0000_0000_0000;
array[20762] <= 16'b0000_0000_0000_0000;
array[20763] <= 16'b0000_0000_0000_0000;
array[20764] <= 16'b0000_0000_0000_0000;
array[20765] <= 16'b0000_0000_0000_0000;
array[20766] <= 16'b0000_0000_0000_0000;
array[20767] <= 16'b0000_0000_0000_0000;
array[20768] <= 16'b0000_0000_0000_0000;
array[20769] <= 16'b0000_0000_0000_0000;
array[20770] <= 16'b0000_0000_0000_0000;
array[20771] <= 16'b0000_0000_0000_0000;
array[20772] <= 16'b0000_0000_0000_0000;
array[20773] <= 16'b0000_0000_0000_0000;
array[20774] <= 16'b0000_0000_0000_0000;
array[20775] <= 16'b0000_0000_0000_0000;
array[20776] <= 16'b0000_0000_0000_0000;
array[20777] <= 16'b0000_0000_0000_0000;
array[20778] <= 16'b0000_0000_0000_0000;
array[20779] <= 16'b0000_0000_0000_0000;
array[20780] <= 16'b0000_0000_0000_0000;
array[20781] <= 16'b0000_0000_0000_0000;
array[20782] <= 16'b0000_0000_0000_0000;
array[20783] <= 16'b0000_0000_0000_0000;
array[20784] <= 16'b0000_0000_0000_0000;
array[20785] <= 16'b0000_0000_0000_0000;
array[20786] <= 16'b0000_0000_0000_0000;
array[20787] <= 16'b0000_0000_0000_0000;
array[20788] <= 16'b0000_0000_0000_0000;
array[20789] <= 16'b0000_0000_0000_0000;
array[20790] <= 16'b0000_0000_0000_0000;
array[20791] <= 16'b0000_0000_0000_0000;
array[20792] <= 16'b0000_0000_0000_0000;
array[20793] <= 16'b0000_0000_0000_0000;
array[20794] <= 16'b0000_0000_0000_0000;
array[20795] <= 16'b0000_0000_0000_0000;
array[20796] <= 16'b0000_0000_0000_0000;
array[20797] <= 16'b0000_0000_0000_0000;
array[20798] <= 16'b0000_0000_0000_0000;
array[20799] <= 16'b0000_0000_0000_0000;
array[20800] <= 16'b0000_0000_0000_0000;
array[20801] <= 16'b0000_0000_0000_0000;
array[20802] <= 16'b0000_0000_0000_0000;
array[20803] <= 16'b0000_0000_0000_0000;
array[20804] <= 16'b0000_0000_0000_0000;
array[20805] <= 16'b0000_0000_0000_0000;
array[20806] <= 16'b0000_0000_0000_0000;
array[20807] <= 16'b0000_0000_0000_0000;
array[20808] <= 16'b0000_0000_0000_0000;
array[20809] <= 16'b0000_0000_0000_0000;
array[20810] <= 16'b0000_0000_0000_0000;
array[20811] <= 16'b0000_0000_0000_0000;
array[20812] <= 16'b0000_0000_0000_0000;
array[20813] <= 16'b0000_0000_0000_0000;
array[20814] <= 16'b0000_0000_0000_0000;
array[20815] <= 16'b0000_0000_0000_0000;
array[20816] <= 16'b0000_0000_0000_0000;
array[20817] <= 16'b0000_0000_0000_0000;
array[20818] <= 16'b0000_0000_0000_0000;
array[20819] <= 16'b0000_0000_0000_0000;
array[20820] <= 16'b0000_0000_0000_0000;
array[20821] <= 16'b0000_0000_0000_0000;
array[20822] <= 16'b0000_0000_0000_0000;
array[20823] <= 16'b0000_0000_0000_0000;
array[20824] <= 16'b0000_0000_0000_0000;
array[20825] <= 16'b0000_0000_0000_0000;
array[20826] <= 16'b0000_0000_0000_0000;
array[20827] <= 16'b0000_0000_0000_0000;
array[20828] <= 16'b0000_0000_0000_0000;
array[20829] <= 16'b0000_0000_0000_0000;
array[20830] <= 16'b0000_0000_0000_0000;
array[20831] <= 16'b0000_0000_0000_0000;
array[20832] <= 16'b0000_0000_0000_0000;
array[20833] <= 16'b0000_0000_0000_0000;
array[20834] <= 16'b0000_0000_0000_0000;
array[20835] <= 16'b0000_0000_0000_0000;
array[20836] <= 16'b0000_0000_0000_0000;
array[20837] <= 16'b0000_0000_0000_0000;
array[20838] <= 16'b0000_0000_0000_0000;
array[20839] <= 16'b0000_0000_0000_0000;
array[20840] <= 16'b0000_0000_0000_0000;
array[20841] <= 16'b0000_0000_0000_0000;
array[20842] <= 16'b0000_0000_0000_0000;
array[20843] <= 16'b0000_0000_0000_0000;
array[20844] <= 16'b0000_0000_0000_0000;
array[20845] <= 16'b0000_0000_0000_0000;
array[20846] <= 16'b0000_0000_0000_0000;
array[20847] <= 16'b0000_0000_0000_0000;
array[20848] <= 16'b0000_0000_0000_0000;
array[20849] <= 16'b0000_0000_0000_0000;
array[20850] <= 16'b0000_0000_0000_0000;
array[20851] <= 16'b0000_0000_0000_0000;
array[20852] <= 16'b0000_0000_0000_0000;
array[20853] <= 16'b0000_0000_0000_0000;
array[20854] <= 16'b0000_0000_0000_0000;
array[20855] <= 16'b0000_0000_0000_0000;
array[20856] <= 16'b0000_0000_0000_0000;
array[20857] <= 16'b0000_0000_0000_0000;
array[20858] <= 16'b0000_0000_0000_0000;
array[20859] <= 16'b0000_0000_0000_0000;
array[20860] <= 16'b0000_0000_0000_0000;
array[20861] <= 16'b0000_0000_0000_0000;
array[20862] <= 16'b0000_0000_0000_0000;
array[20863] <= 16'b0000_0000_0000_0000;
array[20864] <= 16'b0000_0000_0000_0000;
array[20865] <= 16'b0000_0000_0000_0000;
array[20866] <= 16'b0000_0000_0000_0000;
array[20867] <= 16'b0000_0000_0000_0000;
array[20868] <= 16'b0000_0000_0000_0000;
array[20869] <= 16'b0000_0000_0000_0000;
array[20870] <= 16'b0000_0000_0000_0000;
array[20871] <= 16'b0000_0000_0000_0000;
array[20872] <= 16'b0000_0000_0000_0000;
array[20873] <= 16'b0000_0000_0000_0000;
array[20874] <= 16'b0000_0000_0000_0000;
array[20875] <= 16'b0000_0000_0000_0000;
array[20876] <= 16'b0000_0000_0000_0000;
array[20877] <= 16'b0000_0000_0000_0000;
array[20878] <= 16'b0000_0000_0000_0000;
array[20879] <= 16'b0000_0000_0000_0000;
array[20880] <= 16'b0000_0000_0000_0000;
array[20881] <= 16'b0000_0000_0000_0000;
array[20882] <= 16'b0000_0000_0000_0000;
array[20883] <= 16'b0000_0000_0000_0000;
array[20884] <= 16'b0000_0000_0000_0000;
array[20885] <= 16'b0000_0000_0000_0000;
array[20886] <= 16'b0000_0000_0000_0000;
array[20887] <= 16'b0000_0000_0000_0000;
array[20888] <= 16'b0000_0000_0000_0000;
array[20889] <= 16'b0000_0000_0000_0000;
array[20890] <= 16'b0000_0000_0000_0000;
array[20891] <= 16'b0000_0000_0000_0000;
array[20892] <= 16'b0000_0000_0000_0000;
array[20893] <= 16'b0000_0000_0000_0000;
array[20894] <= 16'b0000_0000_0000_0000;
array[20895] <= 16'b0000_0000_0000_0000;
array[20896] <= 16'b0000_0000_0000_0000;
array[20897] <= 16'b0000_0000_0000_0000;
array[20898] <= 16'b0000_0000_0000_0000;
array[20899] <= 16'b0000_0000_0000_0000;
array[20900] <= 16'b0000_0000_0000_0000;
array[20901] <= 16'b0000_0000_0000_0000;
array[20902] <= 16'b0000_0000_0000_0000;
array[20903] <= 16'b0000_0000_0000_0000;
array[20904] <= 16'b0000_0000_0000_0000;
array[20905] <= 16'b0000_0000_0000_0000;
array[20906] <= 16'b0000_0000_0000_0000;
array[20907] <= 16'b0000_0000_0000_0000;
array[20908] <= 16'b0000_0000_0000_0000;
array[20909] <= 16'b0000_0000_0000_0000;
array[20910] <= 16'b0000_0000_0000_0000;
array[20911] <= 16'b0000_0000_0000_0000;
array[20912] <= 16'b0000_0000_0000_0000;
array[20913] <= 16'b0000_0000_0000_0000;
array[20914] <= 16'b0000_0000_0000_0000;
array[20915] <= 16'b0000_0000_0000_0000;
array[20916] <= 16'b0000_0000_0000_0000;
array[20917] <= 16'b0000_0000_0000_0000;
array[20918] <= 16'b0000_0000_0000_0000;
array[20919] <= 16'b0000_0000_0000_0000;
array[20920] <= 16'b0000_0000_0000_0000;
array[20921] <= 16'b0000_0000_0000_0000;
array[20922] <= 16'b0000_0000_0000_0000;
array[20923] <= 16'b0000_0000_0000_0000;
array[20924] <= 16'b0000_0000_0000_0000;
array[20925] <= 16'b0000_0000_0000_0000;
array[20926] <= 16'b0000_0000_0000_0000;
array[20927] <= 16'b0000_0000_0000_0000;
array[20928] <= 16'b0000_0000_0000_0000;
array[20929] <= 16'b0000_0000_0000_0000;
array[20930] <= 16'b0000_0000_0000_0000;
array[20931] <= 16'b0000_0000_0000_0000;
array[20932] <= 16'b0000_0000_0000_0000;
array[20933] <= 16'b0000_0000_0000_0000;
array[20934] <= 16'b0000_0000_0000_0000;
array[20935] <= 16'b0000_0000_0000_0000;
array[20936] <= 16'b0000_0000_0000_0000;
array[20937] <= 16'b0000_0000_0000_0000;
array[20938] <= 16'b0000_0000_0000_0000;
array[20939] <= 16'b0000_0000_0000_0000;
array[20940] <= 16'b0000_0000_0000_0000;
array[20941] <= 16'b0000_0000_0000_0000;
array[20942] <= 16'b0000_0000_0000_0000;
array[20943] <= 16'b0000_0000_0000_0000;
array[20944] <= 16'b0000_0000_0000_0000;
array[20945] <= 16'b0000_0000_0000_0000;
array[20946] <= 16'b0000_0000_0000_0000;
array[20947] <= 16'b0000_0000_0000_0000;
array[20948] <= 16'b0000_0000_0000_0000;
array[20949] <= 16'b0000_0000_0000_0000;
array[20950] <= 16'b0000_0000_0000_0000;
array[20951] <= 16'b0000_0000_0000_0000;
array[20952] <= 16'b0000_0000_0000_0000;
array[20953] <= 16'b0000_0000_0000_0000;
array[20954] <= 16'b0000_0000_0000_0000;
array[20955] <= 16'b0000_0000_0000_0000;
array[20956] <= 16'b0000_0000_0000_0000;
array[20957] <= 16'b0000_0000_0000_0000;
array[20958] <= 16'b0000_0000_0000_0000;
array[20959] <= 16'b0000_0000_0000_0000;
array[20960] <= 16'b0000_0000_0000_0000;
array[20961] <= 16'b0000_0000_0000_0000;
array[20962] <= 16'b0000_0000_0000_0000;
array[20963] <= 16'b0000_0000_0000_0000;
array[20964] <= 16'b0000_0000_0000_0000;
array[20965] <= 16'b0000_0000_0000_0000;
array[20966] <= 16'b0000_0000_0000_0000;
array[20967] <= 16'b0000_0000_0000_0000;
array[20968] <= 16'b0000_0000_0000_0000;
array[20969] <= 16'b0000_0000_0000_0000;
array[20970] <= 16'b0000_0000_0000_0000;
array[20971] <= 16'b0000_0000_0000_0000;
array[20972] <= 16'b0000_0000_0000_0000;
array[20973] <= 16'b0000_0000_0000_0000;
array[20974] <= 16'b0000_0000_0000_0000;
array[20975] <= 16'b0000_0000_0000_0000;
array[20976] <= 16'b0000_0000_0000_0000;
array[20977] <= 16'b0000_0000_0000_0000;
array[20978] <= 16'b0000_0000_0000_0000;
array[20979] <= 16'b0000_0000_0000_0000;
array[20980] <= 16'b0000_0000_0000_0000;
array[20981] <= 16'b0000_0000_0000_0000;
array[20982] <= 16'b0000_0000_0000_0000;
array[20983] <= 16'b0000_0000_0000_0000;
array[20984] <= 16'b0000_0000_0000_0000;
array[20985] <= 16'b0000_0000_0000_0000;
array[20986] <= 16'b0000_0000_0000_0000;
array[20987] <= 16'b0000_0000_0000_0000;
array[20988] <= 16'b0000_0000_0000_0000;
array[20989] <= 16'b0000_0000_0000_0000;
array[20990] <= 16'b0000_0000_0000_0000;
array[20991] <= 16'b0000_0000_0000_0000;
array[20992] <= 16'b0000_0000_0000_0000;
array[20993] <= 16'b0000_0000_0000_0000;
array[20994] <= 16'b0000_0000_0000_0000;
array[20995] <= 16'b0000_0000_0000_0000;
array[20996] <= 16'b0000_0000_0000_0000;
array[20997] <= 16'b0000_0000_0000_0000;
array[20998] <= 16'b0000_0000_0000_0000;
array[20999] <= 16'b0000_0000_0000_0000;
array[21000] <= 16'b0000_0000_0000_0000;
array[21001] <= 16'b0000_0000_0000_0000;
array[21002] <= 16'b0000_0000_0000_0000;
array[21003] <= 16'b0000_0000_0000_0000;
array[21004] <= 16'b0000_0000_0000_0000;
array[21005] <= 16'b0000_0000_0000_0000;
array[21006] <= 16'b0000_0000_0000_0000;
array[21007] <= 16'b0000_0000_0000_0000;
array[21008] <= 16'b0000_0000_0000_0000;
array[21009] <= 16'b0000_0000_0000_0000;
array[21010] <= 16'b0000_0000_0000_0000;
array[21011] <= 16'b0000_0000_0000_0000;
array[21012] <= 16'b0000_0000_0000_0000;
array[21013] <= 16'b0000_0000_0000_0000;
array[21014] <= 16'b0000_0000_0000_0000;
array[21015] <= 16'b0000_0000_0000_0000;
array[21016] <= 16'b0000_0000_0000_0000;
array[21017] <= 16'b0000_0000_0000_0000;
array[21018] <= 16'b0000_0000_0000_0000;
array[21019] <= 16'b0000_0000_0000_0000;
array[21020] <= 16'b0000_0000_0000_0000;
array[21021] <= 16'b0000_0000_0000_0000;
array[21022] <= 16'b0000_0000_0000_0000;
array[21023] <= 16'b0000_0000_0000_0000;
array[21024] <= 16'b0000_0000_0000_0000;
array[21025] <= 16'b0000_0000_0000_0000;
array[21026] <= 16'b0000_0000_0000_0000;
array[21027] <= 16'b0000_0000_0000_0000;
array[21028] <= 16'b0000_0000_0000_0000;
array[21029] <= 16'b0000_0000_0000_0000;
array[21030] <= 16'b0000_0000_0000_0000;
array[21031] <= 16'b0000_0000_0000_0000;
array[21032] <= 16'b0000_0000_0000_0000;
array[21033] <= 16'b0000_0000_0000_0000;
array[21034] <= 16'b0000_0000_0000_0000;
array[21035] <= 16'b0000_0000_0000_0000;
array[21036] <= 16'b0000_0000_0000_0000;
array[21037] <= 16'b0000_0000_0000_0000;
array[21038] <= 16'b0000_0000_0000_0000;
array[21039] <= 16'b0000_0000_0000_0000;
array[21040] <= 16'b0000_0000_0000_0000;
array[21041] <= 16'b0000_0000_0000_0000;
array[21042] <= 16'b0000_0000_0000_0000;
array[21043] <= 16'b0000_0000_0000_0000;
array[21044] <= 16'b0000_0000_0000_0000;
array[21045] <= 16'b0000_0000_0000_0000;
array[21046] <= 16'b0000_0000_0000_0000;
array[21047] <= 16'b0000_0000_0000_0000;
array[21048] <= 16'b0000_0000_0000_0000;
array[21049] <= 16'b0000_0000_0000_0000;
array[21050] <= 16'b0000_0000_0000_0000;
array[21051] <= 16'b0000_0000_0000_0000;
array[21052] <= 16'b0000_0000_0000_0000;
array[21053] <= 16'b0000_0000_0000_0000;
array[21054] <= 16'b0000_0000_0000_0000;
array[21055] <= 16'b0000_0000_0000_0000;
array[21056] <= 16'b0000_0000_0000_0000;
array[21057] <= 16'b0000_0000_0000_0000;
array[21058] <= 16'b0000_0000_0000_0000;
array[21059] <= 16'b0000_0000_0000_0000;
array[21060] <= 16'b0000_0000_0000_0000;
array[21061] <= 16'b0000_0000_0000_0000;
array[21062] <= 16'b0000_0000_0000_0000;
array[21063] <= 16'b0000_0000_0000_0000;
array[21064] <= 16'b0000_0000_0000_0000;
array[21065] <= 16'b0000_0000_0000_0000;
array[21066] <= 16'b0000_0000_0000_0000;
array[21067] <= 16'b0000_0000_0000_0000;
array[21068] <= 16'b0000_0000_0000_0000;
array[21069] <= 16'b0000_0000_0000_0000;
array[21070] <= 16'b0000_0000_0000_0000;
array[21071] <= 16'b0000_0000_0000_0000;
array[21072] <= 16'b0000_0000_0000_0000;
array[21073] <= 16'b0000_0000_0000_0000;
array[21074] <= 16'b0000_0000_0000_0000;
array[21075] <= 16'b0000_0000_0000_0000;
array[21076] <= 16'b0000_0000_0000_0000;
array[21077] <= 16'b0000_0000_0000_0000;
array[21078] <= 16'b0000_0000_0000_0000;
array[21079] <= 16'b0000_0000_0000_0000;
array[21080] <= 16'b0000_0000_0000_0000;
array[21081] <= 16'b0000_0000_0000_0000;
array[21082] <= 16'b0000_0000_0000_0000;
array[21083] <= 16'b0000_0000_0000_0000;
array[21084] <= 16'b0000_0000_0000_0000;
array[21085] <= 16'b0000_0000_0000_0000;
array[21086] <= 16'b0000_0000_0000_0000;
array[21087] <= 16'b0000_0000_0000_0000;
array[21088] <= 16'b0000_0000_0000_0000;
array[21089] <= 16'b0000_0000_0000_0000;
array[21090] <= 16'b0000_0000_0000_0000;
array[21091] <= 16'b0000_0000_0000_0000;
array[21092] <= 16'b0000_0000_0000_0000;
array[21093] <= 16'b0000_0000_0000_0000;
array[21094] <= 16'b0000_0000_0000_0000;
array[21095] <= 16'b0000_0000_0000_0000;
array[21096] <= 16'b0000_0000_0000_0000;
array[21097] <= 16'b0000_0000_0000_0000;
array[21098] <= 16'b0000_0000_0000_0000;
array[21099] <= 16'b0000_0000_0000_0000;
array[21100] <= 16'b0000_0000_0000_0000;
array[21101] <= 16'b0000_0000_0000_0000;
array[21102] <= 16'b0000_0000_0000_0000;
array[21103] <= 16'b0000_0000_0000_0000;
array[21104] <= 16'b0000_0000_0000_0000;
array[21105] <= 16'b0000_0000_0000_0000;
array[21106] <= 16'b0000_0000_0000_0000;
array[21107] <= 16'b0000_0000_0000_0000;
array[21108] <= 16'b0000_0000_0000_0000;
array[21109] <= 16'b0000_0000_0000_0000;
array[21110] <= 16'b0000_0000_0000_0000;
array[21111] <= 16'b0000_0000_0000_0000;
array[21112] <= 16'b0000_0000_0000_0000;
array[21113] <= 16'b0000_0000_0000_0000;
array[21114] <= 16'b0000_0000_0000_0000;
array[21115] <= 16'b0000_0000_0000_0000;
array[21116] <= 16'b0000_0000_0000_0000;
array[21117] <= 16'b0000_0000_0000_0000;
array[21118] <= 16'b0000_0000_0000_0000;
array[21119] <= 16'b0000_0000_0000_0000;
array[21120] <= 16'b0000_0000_0000_0000;
array[21121] <= 16'b0000_0000_0000_0000;
array[21122] <= 16'b0000_0000_0000_0000;
array[21123] <= 16'b0000_0000_0000_0000;
array[21124] <= 16'b0000_0000_0000_0000;
array[21125] <= 16'b0000_0000_0000_0000;
array[21126] <= 16'b0000_0000_0000_0000;
array[21127] <= 16'b0000_0000_0000_0000;
array[21128] <= 16'b0000_0000_0000_0000;
array[21129] <= 16'b0000_0000_0000_0000;
array[21130] <= 16'b0000_0000_0000_0000;
array[21131] <= 16'b0000_0000_0000_0000;
array[21132] <= 16'b0000_0000_0000_0000;
array[21133] <= 16'b0000_0000_0000_0000;
array[21134] <= 16'b0000_0000_0000_0000;
array[21135] <= 16'b0000_0000_0000_0000;
array[21136] <= 16'b0000_0000_0000_0000;
array[21137] <= 16'b0000_0000_0000_0000;
array[21138] <= 16'b0000_0000_0000_0000;
array[21139] <= 16'b0000_0000_0000_0000;
array[21140] <= 16'b0000_0000_0000_0000;
array[21141] <= 16'b0000_0000_0000_0000;
array[21142] <= 16'b0000_0000_0000_0000;
array[21143] <= 16'b0000_0000_0000_0000;
array[21144] <= 16'b0000_0000_0000_0000;
array[21145] <= 16'b0000_0000_0000_0000;
array[21146] <= 16'b0000_0000_0000_0000;
array[21147] <= 16'b0000_0000_0000_0000;
array[21148] <= 16'b0000_0000_0000_0000;
array[21149] <= 16'b0000_0000_0000_0000;
array[21150] <= 16'b0000_0000_0000_0000;
array[21151] <= 16'b0000_0000_0000_0000;
array[21152] <= 16'b0000_0000_0000_0000;
array[21153] <= 16'b0000_0000_0000_0000;
array[21154] <= 16'b0000_0000_0000_0000;
array[21155] <= 16'b0000_0000_0000_0000;
array[21156] <= 16'b0000_0000_0000_0000;
array[21157] <= 16'b0000_0000_0000_0000;
array[21158] <= 16'b0000_0000_0000_0000;
array[21159] <= 16'b0000_0000_0000_0000;
array[21160] <= 16'b0000_0000_0000_0000;
array[21161] <= 16'b0000_0000_0000_0000;
array[21162] <= 16'b0000_0000_0000_0000;
array[21163] <= 16'b0000_0000_0000_0000;
array[21164] <= 16'b0000_0000_0000_0000;
array[21165] <= 16'b0000_0000_0000_0000;
array[21166] <= 16'b0000_0000_0000_0000;
array[21167] <= 16'b0000_0000_0000_0000;
array[21168] <= 16'b0000_0000_0000_0000;
array[21169] <= 16'b0000_0000_0000_0000;
array[21170] <= 16'b0000_0000_0000_0000;
array[21171] <= 16'b0000_0000_0000_0000;
array[21172] <= 16'b0000_0000_0000_0000;
array[21173] <= 16'b0000_0000_0000_0000;
array[21174] <= 16'b0000_0000_0000_0000;
array[21175] <= 16'b0000_0000_0000_0000;
array[21176] <= 16'b0000_0000_0000_0000;
array[21177] <= 16'b0000_0000_0000_0000;
array[21178] <= 16'b0000_0000_0000_0000;
array[21179] <= 16'b0000_0000_0000_0000;
array[21180] <= 16'b0000_0000_0000_0000;
array[21181] <= 16'b0000_0000_0000_0000;
array[21182] <= 16'b0000_0000_0000_0000;
array[21183] <= 16'b0000_0000_0000_0000;
array[21184] <= 16'b0000_0000_0000_0000;
array[21185] <= 16'b0000_0000_0000_0000;
array[21186] <= 16'b0000_0000_0000_0000;
array[21187] <= 16'b0000_0000_0000_0000;
array[21188] <= 16'b0000_0000_0000_0000;
array[21189] <= 16'b0000_0000_0000_0000;
array[21190] <= 16'b0000_0000_0000_0000;
array[21191] <= 16'b0000_0000_0000_0000;
array[21192] <= 16'b0000_0000_0000_0000;
array[21193] <= 16'b0000_0000_0000_0000;
array[21194] <= 16'b0000_0000_0000_0000;
array[21195] <= 16'b0000_0000_0000_0000;
array[21196] <= 16'b0000_0000_0000_0000;
array[21197] <= 16'b0000_0000_0000_0000;
array[21198] <= 16'b0000_0000_0000_0000;
array[21199] <= 16'b0000_0000_0000_0000;
array[21200] <= 16'b0000_0000_0000_0000;
array[21201] <= 16'b0000_0000_0000_0000;
array[21202] <= 16'b0000_0000_0000_0000;
array[21203] <= 16'b0000_0000_0000_0000;
array[21204] <= 16'b0000_0000_0000_0000;
array[21205] <= 16'b0000_0000_0000_0000;
array[21206] <= 16'b0000_0000_0000_0000;
array[21207] <= 16'b0000_0000_0000_0000;
array[21208] <= 16'b0000_0000_0000_0000;
array[21209] <= 16'b0000_0000_0000_0000;
array[21210] <= 16'b0000_0000_0000_0000;
array[21211] <= 16'b0000_0000_0000_0000;
array[21212] <= 16'b0000_0000_0000_0000;
array[21213] <= 16'b0000_0000_0000_0000;
array[21214] <= 16'b0000_0000_0000_0000;
array[21215] <= 16'b0000_0000_0000_0000;
array[21216] <= 16'b0000_0000_0000_0000;
array[21217] <= 16'b0000_0000_0000_0000;
array[21218] <= 16'b0000_0000_0000_0000;
array[21219] <= 16'b0000_0000_0000_0000;
array[21220] <= 16'b0000_0000_0000_0000;
array[21221] <= 16'b0000_0000_0000_0000;
array[21222] <= 16'b0000_0000_0000_0000;
array[21223] <= 16'b0000_0000_0000_0000;
array[21224] <= 16'b0000_0000_0000_0000;
array[21225] <= 16'b0000_0000_0000_0000;
array[21226] <= 16'b0000_0000_0000_0000;
array[21227] <= 16'b0000_0000_0000_0000;
array[21228] <= 16'b0000_0000_0000_0000;
array[21229] <= 16'b0000_0000_0000_0000;
array[21230] <= 16'b0000_0000_0000_0000;
array[21231] <= 16'b0000_0000_0000_0000;
array[21232] <= 16'b0000_0000_0000_0000;
array[21233] <= 16'b0000_0000_0000_0000;
array[21234] <= 16'b0000_0000_0000_0000;
array[21235] <= 16'b0000_0000_0000_0000;
array[21236] <= 16'b0000_0000_0000_0000;
array[21237] <= 16'b0000_0000_0000_0000;
array[21238] <= 16'b0000_0000_0000_0000;
array[21239] <= 16'b0000_0000_0000_0000;
array[21240] <= 16'b0000_0000_0000_0000;
array[21241] <= 16'b0000_0000_0000_0000;
array[21242] <= 16'b0000_0000_0000_0000;
array[21243] <= 16'b0000_0000_0000_0000;
array[21244] <= 16'b0000_0000_0000_0000;
array[21245] <= 16'b0000_0000_0000_0000;
array[21246] <= 16'b0000_0000_0000_0000;
array[21247] <= 16'b0000_0000_0000_0000;
array[21248] <= 16'b0000_0000_0000_0000;
array[21249] <= 16'b0000_0000_0000_0000;
array[21250] <= 16'b0000_0000_0000_0000;
array[21251] <= 16'b0000_0000_0000_0000;
array[21252] <= 16'b0000_0000_0000_0000;
array[21253] <= 16'b0000_0000_0000_0000;
array[21254] <= 16'b0000_0000_0000_0000;
array[21255] <= 16'b0000_0000_0000_0000;
array[21256] <= 16'b0000_0000_0000_0000;
array[21257] <= 16'b0000_0000_0000_0000;
array[21258] <= 16'b0000_0000_0000_0000;
array[21259] <= 16'b0000_0000_0000_0000;
array[21260] <= 16'b0000_0000_0000_0000;
array[21261] <= 16'b0000_0000_0000_0000;
array[21262] <= 16'b0000_0000_0000_0000;
array[21263] <= 16'b0000_0000_0000_0000;
array[21264] <= 16'b0000_0000_0000_0000;
array[21265] <= 16'b0000_0000_0000_0000;
array[21266] <= 16'b0000_0000_0000_0000;
array[21267] <= 16'b0000_0000_0000_0000;
array[21268] <= 16'b0000_0000_0000_0000;
array[21269] <= 16'b0000_0000_0000_0000;
array[21270] <= 16'b0000_0000_0000_0000;
array[21271] <= 16'b0000_0000_0000_0000;
array[21272] <= 16'b0000_0000_0000_0000;
array[21273] <= 16'b0000_0000_0000_0000;
array[21274] <= 16'b0000_0000_0000_0000;
array[21275] <= 16'b0000_0000_0000_0000;
array[21276] <= 16'b0000_0000_0000_0000;
array[21277] <= 16'b0000_0000_0000_0000;
array[21278] <= 16'b0000_0000_0000_0000;
array[21279] <= 16'b0000_0000_0000_0000;
array[21280] <= 16'b0000_0000_0000_0000;
array[21281] <= 16'b0000_0000_0000_0000;
array[21282] <= 16'b0000_0000_0000_0000;
array[21283] <= 16'b0000_0000_0000_0000;
array[21284] <= 16'b0000_0000_0000_0000;
array[21285] <= 16'b0000_0000_0000_0000;
array[21286] <= 16'b0000_0000_0000_0000;
array[21287] <= 16'b0000_0000_0000_0000;
array[21288] <= 16'b0000_0000_0000_0000;
array[21289] <= 16'b0000_0000_0000_0000;
array[21290] <= 16'b0000_0000_0000_0000;
array[21291] <= 16'b0000_0000_0000_0000;
array[21292] <= 16'b0000_0000_0000_0000;
array[21293] <= 16'b0000_0000_0000_0000;
array[21294] <= 16'b0000_0000_0000_0000;
array[21295] <= 16'b0000_0000_0000_0000;
array[21296] <= 16'b0000_0000_0000_0000;
array[21297] <= 16'b0000_0000_0000_0000;
array[21298] <= 16'b0000_0000_0000_0000;
array[21299] <= 16'b0000_0000_0000_0000;
array[21300] <= 16'b0000_0000_0000_0000;
array[21301] <= 16'b0000_0000_0000_0000;
array[21302] <= 16'b0000_0000_0000_0000;
array[21303] <= 16'b0000_0000_0000_0000;
array[21304] <= 16'b0000_0000_0000_0000;
array[21305] <= 16'b0000_0000_0000_0000;
array[21306] <= 16'b0000_0000_0000_0000;
array[21307] <= 16'b0000_0000_0000_0000;
array[21308] <= 16'b0000_0000_0000_0000;
array[21309] <= 16'b0000_0000_0000_0000;
array[21310] <= 16'b0000_0000_0000_0000;
array[21311] <= 16'b0000_0000_0000_0000;
array[21312] <= 16'b0000_0000_0000_0000;
array[21313] <= 16'b0000_0000_0000_0000;
array[21314] <= 16'b0000_0000_0000_0000;
array[21315] <= 16'b0000_0000_0000_0000;
array[21316] <= 16'b0000_0000_0000_0000;
array[21317] <= 16'b0000_0000_0000_0000;
array[21318] <= 16'b0000_0000_0000_0000;
array[21319] <= 16'b0000_0000_0000_0000;
array[21320] <= 16'b0000_0000_0000_0000;
array[21321] <= 16'b0000_0000_0000_0000;
array[21322] <= 16'b0000_0000_0000_0000;
array[21323] <= 16'b0000_0000_0000_0000;
array[21324] <= 16'b0000_0000_0000_0000;
array[21325] <= 16'b0000_0000_0000_0000;
array[21326] <= 16'b0000_0000_0000_0000;
array[21327] <= 16'b0000_0000_0000_0000;
array[21328] <= 16'b0000_0000_0000_0000;
array[21329] <= 16'b0000_0000_0000_0000;
array[21330] <= 16'b0000_0000_0000_0000;
array[21331] <= 16'b0000_0000_0000_0000;
array[21332] <= 16'b0000_0000_0000_0000;
array[21333] <= 16'b0000_0000_0000_0000;
array[21334] <= 16'b0000_0000_0000_0000;
array[21335] <= 16'b0000_0000_0000_0000;
array[21336] <= 16'b0000_0000_0000_0000;
array[21337] <= 16'b0000_0000_0000_0000;
array[21338] <= 16'b0000_0000_0000_0000;
array[21339] <= 16'b0000_0000_0000_0000;
array[21340] <= 16'b0000_0000_0000_0000;
array[21341] <= 16'b0000_0000_0000_0000;
array[21342] <= 16'b0000_0000_0000_0000;
array[21343] <= 16'b0000_0000_0000_0000;
array[21344] <= 16'b0000_0000_0000_0000;
array[21345] <= 16'b0000_0000_0000_0000;
array[21346] <= 16'b0000_0000_0000_0000;
array[21347] <= 16'b0000_0000_0000_0000;
array[21348] <= 16'b0000_0000_0000_0000;
array[21349] <= 16'b0000_0000_0000_0000;
array[21350] <= 16'b0000_0000_0000_0000;
array[21351] <= 16'b0000_0000_0000_0000;
array[21352] <= 16'b0000_0000_0000_0000;
array[21353] <= 16'b0000_0000_0000_0000;
array[21354] <= 16'b0000_0000_0000_0000;
array[21355] <= 16'b0000_0000_0000_0000;
array[21356] <= 16'b0000_0000_0000_0000;
array[21357] <= 16'b0000_0000_0000_0000;
array[21358] <= 16'b0000_0000_0000_0000;
array[21359] <= 16'b0000_0000_0000_0000;
array[21360] <= 16'b0000_0000_0000_0000;
array[21361] <= 16'b0000_0000_0000_0000;
array[21362] <= 16'b0000_0000_0000_0000;
array[21363] <= 16'b0000_0000_0000_0000;
array[21364] <= 16'b0000_0000_0000_0000;
array[21365] <= 16'b0000_0000_0000_0000;
array[21366] <= 16'b0000_0000_0000_0000;
array[21367] <= 16'b0000_0000_0000_0000;
array[21368] <= 16'b0000_0000_0000_0000;
array[21369] <= 16'b0000_0000_0000_0000;
array[21370] <= 16'b0000_0000_0000_0000;
array[21371] <= 16'b0000_0000_0000_0000;
array[21372] <= 16'b0000_0000_0000_0000;
array[21373] <= 16'b0000_0000_0000_0000;
array[21374] <= 16'b0000_0000_0000_0000;
array[21375] <= 16'b0000_0000_0000_0000;
array[21376] <= 16'b0000_0000_0000_0000;
array[21377] <= 16'b0000_0000_0000_0000;
array[21378] <= 16'b0000_0000_0000_0000;
array[21379] <= 16'b0000_0000_0000_0000;
array[21380] <= 16'b0000_0000_0000_0000;
array[21381] <= 16'b0000_0000_0000_0000;
array[21382] <= 16'b0000_0000_0000_0000;
array[21383] <= 16'b0000_0000_0000_0000;
array[21384] <= 16'b0000_0000_0000_0000;
array[21385] <= 16'b0000_0000_0000_0000;
array[21386] <= 16'b0000_0000_0000_0000;
array[21387] <= 16'b0000_0000_0000_0000;
array[21388] <= 16'b0000_0000_0000_0000;
array[21389] <= 16'b0000_0000_0000_0000;
array[21390] <= 16'b0000_0000_0000_0000;
array[21391] <= 16'b0000_0000_0000_0000;
array[21392] <= 16'b0000_0000_0000_0000;
array[21393] <= 16'b0000_0000_0000_0000;
array[21394] <= 16'b0000_0000_0000_0000;
array[21395] <= 16'b0000_0000_0000_0000;
array[21396] <= 16'b0000_0000_0000_0000;
array[21397] <= 16'b0000_0000_0000_0000;
array[21398] <= 16'b0000_0000_0000_0000;
array[21399] <= 16'b0000_0000_0000_0000;
array[21400] <= 16'b0000_0000_0000_0000;
array[21401] <= 16'b0000_0000_0000_0000;
array[21402] <= 16'b0000_0000_0000_0000;
array[21403] <= 16'b0000_0000_0000_0000;
array[21404] <= 16'b0000_0000_0000_0000;
array[21405] <= 16'b0000_0000_0000_0000;
array[21406] <= 16'b0000_0000_0000_0000;
array[21407] <= 16'b0000_0000_0000_0000;
array[21408] <= 16'b0000_0000_0000_0000;
array[21409] <= 16'b0000_0000_0000_0000;
array[21410] <= 16'b0000_0000_0000_0000;
array[21411] <= 16'b0000_0000_0000_0000;
array[21412] <= 16'b0000_0000_0000_0000;
array[21413] <= 16'b0000_0000_0000_0000;
array[21414] <= 16'b0000_0000_0000_0000;
array[21415] <= 16'b0000_0000_0000_0000;
array[21416] <= 16'b0000_0000_0000_0000;
array[21417] <= 16'b0000_0000_0000_0000;
array[21418] <= 16'b0000_0000_0000_0000;
array[21419] <= 16'b0000_0000_0000_0000;
array[21420] <= 16'b0000_0000_0000_0000;
array[21421] <= 16'b0000_0000_0000_0000;
array[21422] <= 16'b0000_0000_0000_0000;
array[21423] <= 16'b0000_0000_0000_0000;
array[21424] <= 16'b0000_0000_0000_0000;
array[21425] <= 16'b0000_0000_0000_0000;
array[21426] <= 16'b0000_0000_0000_0000;
array[21427] <= 16'b0000_0000_0000_0000;
array[21428] <= 16'b0000_0000_0000_0000;
array[21429] <= 16'b0000_0000_0000_0000;
array[21430] <= 16'b0000_0000_0000_0000;
array[21431] <= 16'b0000_0000_0000_0000;
array[21432] <= 16'b0000_0000_0000_0000;
array[21433] <= 16'b0000_0000_0000_0000;
array[21434] <= 16'b0000_0000_0000_0000;
array[21435] <= 16'b0000_0000_0000_0000;
array[21436] <= 16'b0000_0000_0000_0000;
array[21437] <= 16'b0000_0000_0000_0000;
array[21438] <= 16'b0000_0000_0000_0000;
array[21439] <= 16'b0000_0000_0000_0000;
array[21440] <= 16'b0000_0000_0000_0000;
array[21441] <= 16'b0000_0000_0000_0000;
array[21442] <= 16'b0000_0000_0000_0000;
array[21443] <= 16'b0000_0000_0000_0000;
array[21444] <= 16'b0000_0000_0000_0000;
array[21445] <= 16'b0000_0000_0000_0000;
array[21446] <= 16'b0000_0000_0000_0000;
array[21447] <= 16'b0000_0000_0000_0000;
array[21448] <= 16'b0000_0000_0000_0000;
array[21449] <= 16'b0000_0000_0000_0000;
array[21450] <= 16'b0000_0000_0000_0000;
array[21451] <= 16'b0000_0000_0000_0000;
array[21452] <= 16'b0000_0000_0000_0000;
array[21453] <= 16'b0000_0000_0000_0000;
array[21454] <= 16'b0000_0000_0000_0000;
array[21455] <= 16'b0000_0000_0000_0000;
array[21456] <= 16'b0000_0000_0000_0000;
array[21457] <= 16'b0000_0000_0000_0000;
array[21458] <= 16'b0000_0000_0000_0000;
array[21459] <= 16'b0000_0000_0000_0000;
array[21460] <= 16'b0000_0000_0000_0000;
array[21461] <= 16'b0000_0000_0000_0000;
array[21462] <= 16'b0000_0000_0000_0000;
array[21463] <= 16'b0000_0000_0000_0000;
array[21464] <= 16'b0000_0000_0000_0000;
array[21465] <= 16'b0000_0000_0000_0000;
array[21466] <= 16'b0000_0000_0000_0000;
array[21467] <= 16'b0000_0000_0000_0000;
array[21468] <= 16'b0000_0000_0000_0000;
array[21469] <= 16'b0000_0000_0000_0000;
array[21470] <= 16'b0000_0000_0000_0000;
array[21471] <= 16'b0000_0000_0000_0000;
array[21472] <= 16'b0000_0000_0000_0000;
array[21473] <= 16'b0000_0000_0000_0000;
array[21474] <= 16'b0000_0000_0000_0000;
array[21475] <= 16'b0000_0000_0000_0000;
array[21476] <= 16'b0000_0000_0000_0000;
array[21477] <= 16'b0000_0000_0000_0000;
array[21478] <= 16'b0000_0000_0000_0000;
array[21479] <= 16'b0000_0000_0000_0000;
array[21480] <= 16'b0000_0000_0000_0000;
array[21481] <= 16'b0000_0000_0000_0000;
array[21482] <= 16'b0000_0000_0000_0000;
array[21483] <= 16'b0000_0000_0000_0000;
array[21484] <= 16'b0000_0000_0000_0000;
array[21485] <= 16'b0000_0000_0000_0000;
array[21486] <= 16'b0000_0000_0000_0000;
array[21487] <= 16'b0000_0000_0000_0000;
array[21488] <= 16'b0000_0000_0000_0000;
array[21489] <= 16'b0000_0000_0000_0000;
array[21490] <= 16'b0000_0000_0000_0000;
array[21491] <= 16'b0000_0000_0000_0000;
array[21492] <= 16'b0000_0000_0000_0000;
array[21493] <= 16'b0000_0000_0000_0000;
array[21494] <= 16'b0000_0000_0000_0000;
array[21495] <= 16'b0000_0000_0000_0000;
array[21496] <= 16'b0000_0000_0000_0000;
array[21497] <= 16'b0000_0000_0000_0000;
array[21498] <= 16'b0000_0000_0000_0000;
array[21499] <= 16'b0000_0000_0000_0000;
array[21500] <= 16'b0000_0000_0000_0000;
array[21501] <= 16'b0000_0000_0000_0000;
array[21502] <= 16'b0000_0000_0000_0000;
array[21503] <= 16'b0000_0000_0000_0000;
array[21504] <= 16'b0000_0000_0000_0000;
array[21505] <= 16'b0000_0000_0000_0000;
array[21506] <= 16'b0000_0000_0000_0000;
array[21507] <= 16'b0000_0000_0000_0000;
array[21508] <= 16'b0000_0000_0000_0000;
array[21509] <= 16'b0000_0000_0000_0000;
array[21510] <= 16'b0000_0000_0000_0000;
array[21511] <= 16'b0000_0000_0000_0000;
array[21512] <= 16'b0000_0000_0000_0000;
array[21513] <= 16'b0000_0000_0000_0000;
array[21514] <= 16'b0000_0000_0000_0000;
array[21515] <= 16'b0000_0000_0000_0000;
array[21516] <= 16'b0000_0000_0000_0000;
array[21517] <= 16'b0000_0000_0000_0000;
array[21518] <= 16'b0000_0000_0000_0000;
array[21519] <= 16'b0000_0000_0000_0000;
array[21520] <= 16'b0000_0000_0000_0000;
array[21521] <= 16'b0000_0000_0000_0000;
array[21522] <= 16'b0000_0000_0000_0000;
array[21523] <= 16'b0000_0000_0000_0000;
array[21524] <= 16'b0000_0000_0000_0000;
array[21525] <= 16'b0000_0000_0000_0000;
array[21526] <= 16'b0000_0000_0000_0000;
array[21527] <= 16'b0000_0000_0000_0000;
array[21528] <= 16'b0000_0000_0000_0000;
array[21529] <= 16'b0000_0000_0000_0000;
array[21530] <= 16'b0000_0000_0000_0000;
array[21531] <= 16'b0000_0000_0000_0000;
array[21532] <= 16'b0000_0000_0000_0000;
array[21533] <= 16'b0000_0000_0000_0000;
array[21534] <= 16'b0000_0000_0000_0000;
array[21535] <= 16'b0000_0000_0000_0000;
array[21536] <= 16'b0000_0000_0000_0000;
array[21537] <= 16'b0000_0000_0000_0000;
array[21538] <= 16'b0000_0000_0000_0000;
array[21539] <= 16'b0000_0000_0000_0000;
array[21540] <= 16'b0000_0000_0000_0000;
array[21541] <= 16'b0000_0000_0000_0000;
array[21542] <= 16'b0000_0000_0000_0000;
array[21543] <= 16'b0000_0000_0000_0000;
array[21544] <= 16'b0000_0000_0000_0000;
array[21545] <= 16'b0000_0000_0000_0000;
array[21546] <= 16'b0000_0000_0000_0000;
array[21547] <= 16'b0000_0000_0000_0000;
array[21548] <= 16'b0000_0000_0000_0000;
array[21549] <= 16'b0000_0000_0000_0000;
array[21550] <= 16'b0000_0000_0000_0000;
array[21551] <= 16'b0000_0000_0000_0000;
array[21552] <= 16'b0000_0000_0000_0000;
array[21553] <= 16'b0000_0000_0000_0000;
array[21554] <= 16'b0000_0000_0000_0000;
array[21555] <= 16'b0000_0000_0000_0000;
array[21556] <= 16'b0000_0000_0000_0000;
array[21557] <= 16'b0000_0000_0000_0000;
array[21558] <= 16'b0000_0000_0000_0000;
array[21559] <= 16'b0000_0000_0000_0000;
array[21560] <= 16'b0000_0000_0000_0000;
array[21561] <= 16'b0000_0000_0000_0000;
array[21562] <= 16'b0000_0000_0000_0000;
array[21563] <= 16'b0000_0000_0000_0000;
array[21564] <= 16'b0000_0000_0000_0000;
array[21565] <= 16'b0000_0000_0000_0000;
array[21566] <= 16'b0000_0000_0000_0000;
array[21567] <= 16'b0000_0000_0000_0000;
array[21568] <= 16'b0000_0000_0000_0000;
array[21569] <= 16'b0000_0000_0000_0000;
array[21570] <= 16'b0000_0000_0000_0000;
array[21571] <= 16'b0000_0000_0000_0000;
array[21572] <= 16'b0000_0000_0000_0000;
array[21573] <= 16'b0000_0000_0000_0000;
array[21574] <= 16'b0000_0000_0000_0000;
array[21575] <= 16'b0000_0000_0000_0000;
array[21576] <= 16'b0000_0000_0000_0000;
array[21577] <= 16'b0000_0000_0000_0000;
array[21578] <= 16'b0000_0000_0000_0000;
array[21579] <= 16'b0000_0000_0000_0000;
array[21580] <= 16'b0000_0000_0000_0000;
array[21581] <= 16'b0000_0000_0000_0000;
array[21582] <= 16'b0000_0000_0000_0000;
array[21583] <= 16'b0000_0000_0000_0000;
array[21584] <= 16'b0000_0000_0000_0000;
array[21585] <= 16'b0000_0000_0000_0000;
array[21586] <= 16'b0000_0000_0000_0000;
array[21587] <= 16'b0000_0000_0000_0000;
array[21588] <= 16'b0000_0000_0000_0000;
array[21589] <= 16'b0000_0000_0000_0000;
array[21590] <= 16'b0000_0000_0000_0000;
array[21591] <= 16'b0000_0000_0000_0000;
array[21592] <= 16'b0000_0000_0000_0000;
array[21593] <= 16'b0000_0000_0000_0000;
array[21594] <= 16'b0000_0000_0000_0000;
array[21595] <= 16'b0000_0000_0000_0000;
array[21596] <= 16'b0000_0000_0000_0000;
array[21597] <= 16'b0000_0000_0000_0000;
array[21598] <= 16'b0000_0000_0000_0000;
array[21599] <= 16'b0000_0000_0000_0000;
array[21600] <= 16'b0000_0000_0000_0000;
array[21601] <= 16'b0000_0000_0000_0000;
array[21602] <= 16'b0000_0000_0000_0000;
array[21603] <= 16'b0000_0000_0000_0000;
array[21604] <= 16'b0000_0000_0000_0000;
array[21605] <= 16'b0000_0000_0000_0000;
array[21606] <= 16'b0000_0000_0000_0000;
array[21607] <= 16'b0000_0000_0000_0000;
array[21608] <= 16'b0000_0000_0000_0000;
array[21609] <= 16'b0000_0000_0000_0000;
array[21610] <= 16'b0000_0000_0000_0000;
array[21611] <= 16'b0000_0000_0000_0000;
array[21612] <= 16'b0000_0000_0000_0000;
array[21613] <= 16'b0000_0000_0000_0000;
array[21614] <= 16'b0000_0000_0000_0000;
array[21615] <= 16'b0000_0000_0000_0000;
array[21616] <= 16'b0000_0000_0000_0000;
array[21617] <= 16'b0000_0000_0000_0000;
array[21618] <= 16'b0000_0000_0000_0000;
array[21619] <= 16'b0000_0000_0000_0000;
array[21620] <= 16'b0000_0000_0000_0000;
array[21621] <= 16'b0000_0000_0000_0000;
array[21622] <= 16'b0000_0000_0000_0000;
array[21623] <= 16'b0000_0000_0000_0000;
array[21624] <= 16'b0000_0000_0000_0000;
array[21625] <= 16'b0000_0000_0000_0000;
array[21626] <= 16'b0000_0000_0000_0000;
array[21627] <= 16'b0000_0000_0000_0000;
array[21628] <= 16'b0000_0000_0000_0000;
array[21629] <= 16'b0000_0000_0000_0000;
array[21630] <= 16'b0000_0000_0000_0000;
array[21631] <= 16'b0000_0000_0000_0000;
array[21632] <= 16'b0000_0000_0000_0000;
array[21633] <= 16'b0000_0000_0000_0000;
array[21634] <= 16'b0000_0000_0000_0000;
array[21635] <= 16'b0000_0000_0000_0000;
array[21636] <= 16'b0000_0000_0000_0000;
array[21637] <= 16'b0000_0000_0000_0000;
array[21638] <= 16'b0000_0000_0000_0000;
array[21639] <= 16'b0000_0000_0000_0000;
array[21640] <= 16'b0000_0000_0000_0000;
array[21641] <= 16'b0000_0000_0000_0000;
array[21642] <= 16'b0000_0000_0000_0000;
array[21643] <= 16'b0000_0000_0000_0000;
array[21644] <= 16'b0000_0000_0000_0000;
array[21645] <= 16'b0000_0000_0000_0000;
array[21646] <= 16'b0000_0000_0000_0000;
array[21647] <= 16'b0000_0000_0000_0000;
array[21648] <= 16'b0000_0000_0000_0000;
array[21649] <= 16'b0000_0000_0000_0000;
array[21650] <= 16'b0000_0000_0000_0000;
array[21651] <= 16'b0000_0000_0000_0000;
array[21652] <= 16'b0000_0000_0000_0000;
array[21653] <= 16'b0000_0000_0000_0000;
array[21654] <= 16'b0000_0000_0000_0000;
array[21655] <= 16'b0000_0000_0000_0000;
array[21656] <= 16'b0000_0000_0000_0000;
array[21657] <= 16'b0000_0000_0000_0000;
array[21658] <= 16'b0000_0000_0000_0000;
array[21659] <= 16'b0000_0000_0000_0000;
array[21660] <= 16'b0000_0000_0000_0000;
array[21661] <= 16'b0000_0000_0000_0000;
array[21662] <= 16'b0000_0000_0000_0000;
array[21663] <= 16'b0000_0000_0000_0000;
array[21664] <= 16'b0000_0000_0000_0000;
array[21665] <= 16'b0000_0000_0000_0000;
array[21666] <= 16'b0000_0000_0000_0000;
array[21667] <= 16'b0000_0000_0000_0000;
array[21668] <= 16'b0000_0000_0000_0000;
array[21669] <= 16'b0000_0000_0000_0000;
array[21670] <= 16'b0000_0000_0000_0000;
array[21671] <= 16'b0000_0000_0000_0000;
array[21672] <= 16'b0000_0000_0000_0000;
array[21673] <= 16'b0000_0000_0000_0000;
array[21674] <= 16'b0000_0000_0000_0000;
array[21675] <= 16'b0000_0000_0000_0000;
array[21676] <= 16'b0000_0000_0000_0000;
array[21677] <= 16'b0000_0000_0000_0000;
array[21678] <= 16'b0000_0000_0000_0000;
array[21679] <= 16'b0000_0000_0000_0000;
array[21680] <= 16'b0000_0000_0000_0000;
array[21681] <= 16'b0000_0000_0000_0000;
array[21682] <= 16'b0000_0000_0000_0000;
array[21683] <= 16'b0000_0000_0000_0000;
array[21684] <= 16'b0000_0000_0000_0000;
array[21685] <= 16'b0000_0000_0000_0000;
array[21686] <= 16'b0000_0000_0000_0000;
array[21687] <= 16'b0000_0000_0000_0000;
array[21688] <= 16'b0000_0000_0000_0000;
array[21689] <= 16'b0000_0000_0000_0000;
array[21690] <= 16'b0000_0000_0000_0000;
array[21691] <= 16'b0000_0000_0000_0000;
array[21692] <= 16'b0000_0000_0000_0000;
array[21693] <= 16'b0000_0000_0000_0000;
array[21694] <= 16'b0000_0000_0000_0000;
array[21695] <= 16'b0000_0000_0000_0000;
array[21696] <= 16'b0000_0000_0000_0000;
array[21697] <= 16'b0000_0000_0000_0000;
array[21698] <= 16'b0000_0000_0000_0000;
array[21699] <= 16'b0000_0000_0000_0000;
array[21700] <= 16'b0000_0000_0000_0000;
array[21701] <= 16'b0000_0000_0000_0000;
array[21702] <= 16'b0000_0000_0000_0000;
array[21703] <= 16'b0000_0000_0000_0000;
array[21704] <= 16'b0000_0000_0000_0000;
array[21705] <= 16'b0000_0000_0000_0000;
array[21706] <= 16'b0000_0000_0000_0000;
array[21707] <= 16'b0000_0000_0000_0000;
array[21708] <= 16'b0000_0000_0000_0000;
array[21709] <= 16'b0000_0000_0000_0000;
array[21710] <= 16'b0000_0000_0000_0000;
array[21711] <= 16'b0000_0000_0000_0000;
array[21712] <= 16'b0000_0000_0000_0000;
array[21713] <= 16'b0000_0000_0000_0000;
array[21714] <= 16'b0000_0000_0000_0000;
array[21715] <= 16'b0000_0000_0000_0000;
array[21716] <= 16'b0000_0000_0000_0000;
array[21717] <= 16'b0000_0000_0000_0000;
array[21718] <= 16'b0000_0000_0000_0000;
array[21719] <= 16'b0000_0000_0000_0000;
array[21720] <= 16'b0000_0000_0000_0000;
array[21721] <= 16'b0000_0000_0000_0000;
array[21722] <= 16'b0000_0000_0000_0000;
array[21723] <= 16'b0000_0000_0000_0000;
array[21724] <= 16'b0000_0000_0000_0000;
array[21725] <= 16'b0000_0000_0000_0000;
array[21726] <= 16'b0000_0000_0000_0000;
array[21727] <= 16'b0000_0000_0000_0000;
array[21728] <= 16'b0000_0000_0000_0000;
array[21729] <= 16'b0000_0000_0000_0000;
array[21730] <= 16'b0000_0000_0000_0000;
array[21731] <= 16'b0000_0000_0000_0000;
array[21732] <= 16'b0000_0000_0000_0000;
array[21733] <= 16'b0000_0000_0000_0000;
array[21734] <= 16'b0000_0000_0000_0000;
array[21735] <= 16'b0000_0000_0000_0000;
array[21736] <= 16'b0000_0000_0000_0000;
array[21737] <= 16'b0000_0000_0000_0000;
array[21738] <= 16'b0000_0000_0000_0000;
array[21739] <= 16'b0000_0000_0000_0000;
array[21740] <= 16'b0000_0000_0000_0000;
array[21741] <= 16'b0000_0000_0000_0000;
array[21742] <= 16'b0000_0000_0000_0000;
array[21743] <= 16'b0000_0000_0000_0000;
array[21744] <= 16'b0000_0000_0000_0000;
array[21745] <= 16'b0000_0000_0000_0000;
array[21746] <= 16'b0000_0000_0000_0000;
array[21747] <= 16'b0000_0000_0000_0000;
array[21748] <= 16'b0000_0000_0000_0000;
array[21749] <= 16'b0000_0000_0000_0000;
array[21750] <= 16'b0000_0000_0000_0000;
array[21751] <= 16'b0000_0000_0000_0000;
array[21752] <= 16'b0000_0000_0000_0000;
array[21753] <= 16'b0000_0000_0000_0000;
array[21754] <= 16'b0000_0000_0000_0000;
array[21755] <= 16'b0000_0000_0000_0000;
array[21756] <= 16'b0000_0000_0000_0000;
array[21757] <= 16'b0000_0000_0000_0000;
array[21758] <= 16'b0000_0000_0000_0000;
array[21759] <= 16'b0000_0000_0000_0000;
array[21760] <= 16'b0000_0000_0000_0000;
array[21761] <= 16'b0000_0000_0000_0000;
array[21762] <= 16'b0000_0000_0000_0000;
array[21763] <= 16'b0000_0000_0000_0000;
array[21764] <= 16'b0000_0000_0000_0000;
array[21765] <= 16'b0000_0000_0000_0000;
array[21766] <= 16'b0000_0000_0000_0000;
array[21767] <= 16'b0000_0000_0000_0000;
array[21768] <= 16'b0000_0000_0000_0000;
array[21769] <= 16'b0000_0000_0000_0000;
array[21770] <= 16'b0000_0000_0000_0000;
array[21771] <= 16'b0000_0000_0000_0000;
array[21772] <= 16'b0000_0000_0000_0000;
array[21773] <= 16'b0000_0000_0000_0000;
array[21774] <= 16'b0000_0000_0000_0000;
array[21775] <= 16'b0000_0000_0000_0000;
array[21776] <= 16'b0000_0000_0000_0000;
array[21777] <= 16'b0000_0000_0000_0000;
array[21778] <= 16'b0000_0000_0000_0000;
array[21779] <= 16'b0000_0000_0000_0000;
array[21780] <= 16'b0000_0000_0000_0000;
array[21781] <= 16'b0000_0000_0000_0000;
array[21782] <= 16'b0000_0000_0000_0000;
array[21783] <= 16'b0000_0000_0000_0000;
array[21784] <= 16'b0000_0000_0000_0000;
array[21785] <= 16'b0000_0000_0000_0000;
array[21786] <= 16'b0000_0000_0000_0000;
array[21787] <= 16'b0000_0000_0000_0000;
array[21788] <= 16'b0000_0000_0000_0000;
array[21789] <= 16'b0000_0000_0000_0000;
array[21790] <= 16'b0000_0000_0000_0000;
array[21791] <= 16'b0000_0000_0000_0000;
array[21792] <= 16'b0000_0000_0000_0000;
array[21793] <= 16'b0000_0000_0000_0000;
array[21794] <= 16'b0000_0000_0000_0000;
array[21795] <= 16'b0000_0000_0000_0000;
array[21796] <= 16'b0000_0000_0000_0000;
array[21797] <= 16'b0000_0000_0000_0000;
array[21798] <= 16'b0000_0000_0000_0000;
array[21799] <= 16'b0000_0000_0000_0000;
array[21800] <= 16'b0000_0000_0000_0000;
array[21801] <= 16'b0000_0000_0000_0000;
array[21802] <= 16'b0000_0000_0000_0000;
array[21803] <= 16'b0000_0000_0000_0000;
array[21804] <= 16'b0000_0000_0000_0000;
array[21805] <= 16'b0000_0000_0000_0000;
array[21806] <= 16'b0000_0000_0000_0000;
array[21807] <= 16'b0000_0000_0000_0000;
array[21808] <= 16'b0000_0000_0000_0000;
array[21809] <= 16'b0000_0000_0000_0000;
array[21810] <= 16'b0000_0000_0000_0000;
array[21811] <= 16'b0000_0000_0000_0000;
array[21812] <= 16'b0000_0000_0000_0000;
array[21813] <= 16'b0000_0000_0000_0000;
array[21814] <= 16'b0000_0000_0000_0000;
array[21815] <= 16'b0000_0000_0000_0000;
array[21816] <= 16'b0000_0000_0000_0000;
array[21817] <= 16'b0000_0000_0000_0000;
array[21818] <= 16'b0000_0000_0000_0000;
array[21819] <= 16'b0000_0000_0000_0000;
array[21820] <= 16'b0000_0000_0000_0000;
array[21821] <= 16'b0000_0000_0000_0000;
array[21822] <= 16'b0000_0000_0000_0000;
array[21823] <= 16'b0000_0000_0000_0000;
array[21824] <= 16'b0000_0000_0000_0000;
array[21825] <= 16'b0000_0000_0000_0000;
array[21826] <= 16'b0000_0000_0000_0000;
array[21827] <= 16'b0000_0000_0000_0000;
array[21828] <= 16'b0000_0000_0000_0000;
array[21829] <= 16'b0000_0000_0000_0000;
array[21830] <= 16'b0000_0000_0000_0000;
array[21831] <= 16'b0000_0000_0000_0000;
array[21832] <= 16'b0000_0000_0000_0000;
array[21833] <= 16'b0000_0000_0000_0000;
array[21834] <= 16'b0000_0000_0000_0000;
array[21835] <= 16'b0000_0000_0000_0000;
array[21836] <= 16'b0000_0000_0000_0000;
array[21837] <= 16'b0000_0000_0000_0000;
array[21838] <= 16'b0000_0000_0000_0000;
array[21839] <= 16'b0000_0000_0000_0000;
array[21840] <= 16'b0000_0000_0000_0000;
array[21841] <= 16'b0000_0000_0000_0000;
array[21842] <= 16'b0000_0000_0000_0000;
array[21843] <= 16'b0000_0000_0000_0000;
array[21844] <= 16'b0000_0000_0000_0000;
array[21845] <= 16'b0000_0000_0000_0000;
array[21846] <= 16'b0000_0000_0000_0000;
array[21847] <= 16'b0000_0000_0000_0000;
array[21848] <= 16'b0000_0000_0000_0000;
array[21849] <= 16'b0000_0000_0000_0000;
array[21850] <= 16'b0000_0000_0000_0000;
array[21851] <= 16'b0000_0000_0000_0000;
array[21852] <= 16'b0000_0000_0000_0000;
array[21853] <= 16'b0000_0000_0000_0000;
array[21854] <= 16'b0000_0000_0000_0000;
array[21855] <= 16'b0000_0000_0000_0000;
array[21856] <= 16'b0000_0000_0000_0000;
array[21857] <= 16'b0000_0000_0000_0000;
array[21858] <= 16'b0000_0000_0000_0000;
array[21859] <= 16'b0000_0000_0000_0000;
array[21860] <= 16'b0000_0000_0000_0000;
array[21861] <= 16'b0000_0000_0000_0000;
array[21862] <= 16'b0000_0000_0000_0000;
array[21863] <= 16'b0000_0000_0000_0000;
array[21864] <= 16'b0000_0000_0000_0000;
array[21865] <= 16'b0000_0000_0000_0000;
array[21866] <= 16'b0000_0000_0000_0000;
array[21867] <= 16'b0000_0000_0000_0000;
array[21868] <= 16'b0000_0000_0000_0000;
array[21869] <= 16'b0000_0000_0000_0000;
array[21870] <= 16'b0000_0000_0000_0000;
array[21871] <= 16'b0000_0000_0000_0000;
array[21872] <= 16'b0000_0000_0000_0000;
array[21873] <= 16'b0000_0000_0000_0000;
array[21874] <= 16'b0000_0000_0000_0000;
array[21875] <= 16'b0000_0000_0000_0000;
array[21876] <= 16'b0000_0000_0000_0000;
array[21877] <= 16'b0000_0000_0000_0000;
array[21878] <= 16'b0000_0000_0000_0000;
array[21879] <= 16'b0000_0000_0000_0000;
array[21880] <= 16'b0000_0000_0000_0000;
array[21881] <= 16'b0000_0000_0000_0000;
array[21882] <= 16'b0000_0000_0000_0000;
array[21883] <= 16'b0000_0000_0000_0000;
array[21884] <= 16'b0000_0000_0000_0000;
array[21885] <= 16'b0000_0000_0000_0000;
array[21886] <= 16'b0000_0000_0000_0000;
array[21887] <= 16'b0000_0000_0000_0000;
array[21888] <= 16'b0000_0000_0000_0000;
array[21889] <= 16'b0000_0000_0000_0000;
array[21890] <= 16'b0000_0000_0000_0000;
array[21891] <= 16'b0000_0000_0000_0000;
array[21892] <= 16'b0000_0000_0000_0000;
array[21893] <= 16'b0000_0000_0000_0000;
array[21894] <= 16'b0000_0000_0000_0000;
array[21895] <= 16'b0000_0000_0000_0000;
array[21896] <= 16'b0000_0000_0000_0000;
array[21897] <= 16'b0000_0000_0000_0000;
array[21898] <= 16'b0000_0000_0000_0000;
array[21899] <= 16'b0000_0000_0000_0000;
array[21900] <= 16'b0000_0000_0000_0000;
array[21901] <= 16'b0000_0000_0000_0000;
array[21902] <= 16'b0000_0000_0000_0000;
array[21903] <= 16'b0000_0000_0000_0000;
array[21904] <= 16'b0000_0000_0000_0000;
array[21905] <= 16'b0000_0000_0000_0000;
array[21906] <= 16'b0000_0000_0000_0000;
array[21907] <= 16'b0000_0000_0000_0000;
array[21908] <= 16'b0000_0000_0000_0000;
array[21909] <= 16'b0000_0000_0000_0000;
array[21910] <= 16'b0000_0000_0000_0000;
array[21911] <= 16'b0000_0000_0000_0000;
array[21912] <= 16'b0000_0000_0000_0000;
array[21913] <= 16'b0000_0000_0000_0000;
array[21914] <= 16'b0000_0000_0000_0000;
array[21915] <= 16'b0000_0000_0000_0000;
array[21916] <= 16'b0000_0000_0000_0000;
array[21917] <= 16'b0000_0000_0000_0000;
array[21918] <= 16'b0000_0000_0000_0000;
array[21919] <= 16'b0000_0000_0000_0000;
array[21920] <= 16'b0000_0000_0000_0000;
array[21921] <= 16'b0000_0000_0000_0000;
array[21922] <= 16'b0000_0000_0000_0000;
array[21923] <= 16'b0000_0000_0000_0000;
array[21924] <= 16'b0000_0000_0000_0000;
array[21925] <= 16'b0000_0000_0000_0000;
array[21926] <= 16'b0000_0000_0000_0000;
array[21927] <= 16'b0000_0000_0000_0000;
array[21928] <= 16'b0000_0000_0000_0000;
array[21929] <= 16'b0000_0000_0000_0000;
array[21930] <= 16'b0000_0000_0000_0000;
array[21931] <= 16'b0000_0000_0000_0000;
array[21932] <= 16'b0000_0000_0000_0000;
array[21933] <= 16'b0000_0000_0000_0000;
array[21934] <= 16'b0000_0000_0000_0000;
array[21935] <= 16'b0000_0000_0000_0000;
array[21936] <= 16'b0000_0000_0000_0000;
array[21937] <= 16'b0000_0000_0000_0000;
array[21938] <= 16'b0000_0000_0000_0000;
array[21939] <= 16'b0000_0000_0000_0000;
array[21940] <= 16'b0000_0000_0000_0000;
array[21941] <= 16'b0000_0000_0000_0000;
array[21942] <= 16'b0000_0000_0000_0000;
array[21943] <= 16'b0000_0000_0000_0000;
array[21944] <= 16'b0000_0000_0000_0000;
array[21945] <= 16'b0000_0000_0000_0000;
array[21946] <= 16'b0000_0000_0000_0000;
array[21947] <= 16'b0000_0000_0000_0000;
array[21948] <= 16'b0000_0000_0000_0000;
array[21949] <= 16'b0000_0000_0000_0000;
array[21950] <= 16'b0000_0000_0000_0000;
array[21951] <= 16'b0000_0000_0000_0000;
array[21952] <= 16'b0000_0000_0000_0000;
array[21953] <= 16'b0000_0000_0000_0000;
array[21954] <= 16'b0000_0000_0000_0000;
array[21955] <= 16'b0000_0000_0000_0000;
array[21956] <= 16'b0000_0000_0000_0000;
array[21957] <= 16'b0000_0000_0000_0000;
array[21958] <= 16'b0000_0000_0000_0000;
array[21959] <= 16'b0000_0000_0000_0000;
array[21960] <= 16'b0000_0000_0000_0000;
array[21961] <= 16'b0000_0000_0000_0000;
array[21962] <= 16'b0000_0000_0000_0000;
array[21963] <= 16'b0000_0000_0000_0000;
array[21964] <= 16'b0000_0000_0000_0000;
array[21965] <= 16'b0000_0000_0000_0000;
array[21966] <= 16'b0000_0000_0000_0000;
array[21967] <= 16'b0000_0000_0000_0000;
array[21968] <= 16'b0000_0000_0000_0000;
array[21969] <= 16'b0000_0000_0000_0000;
array[21970] <= 16'b0000_0000_0000_0000;
array[21971] <= 16'b0000_0000_0000_0000;
array[21972] <= 16'b0000_0000_0000_0000;
array[21973] <= 16'b0000_0000_0000_0000;
array[21974] <= 16'b0000_0000_0000_0000;
array[21975] <= 16'b0000_0000_0000_0000;
array[21976] <= 16'b0000_0000_0000_0000;
array[21977] <= 16'b0000_0000_0000_0000;
array[21978] <= 16'b0000_0000_0000_0000;
array[21979] <= 16'b0000_0000_0000_0000;
array[21980] <= 16'b0000_0000_0000_0000;
array[21981] <= 16'b0000_0000_0000_0000;
array[21982] <= 16'b0000_0000_0000_0000;
array[21983] <= 16'b0000_0000_0000_0000;
array[21984] <= 16'b0000_0000_0000_0000;
array[21985] <= 16'b0000_0000_0000_0000;
array[21986] <= 16'b0000_0000_0000_0000;
array[21987] <= 16'b0000_0000_0000_0000;
array[21988] <= 16'b0000_0000_0000_0000;
array[21989] <= 16'b0000_0000_0000_0000;
array[21990] <= 16'b0000_0000_0000_0000;
array[21991] <= 16'b0000_0000_0000_0000;
array[21992] <= 16'b0000_0000_0000_0000;
array[21993] <= 16'b0000_0000_0000_0000;
array[21994] <= 16'b0000_0000_0000_0000;
array[21995] <= 16'b0000_0000_0000_0000;
array[21996] <= 16'b0000_0000_0000_0000;
array[21997] <= 16'b0000_0000_0000_0000;
array[21998] <= 16'b0000_0000_0000_0000;
array[21999] <= 16'b0000_0000_0000_0000;
array[22000] <= 16'b0000_0000_0000_0000;
array[22001] <= 16'b0000_0000_0000_0000;
array[22002] <= 16'b0000_0000_0000_0000;
array[22003] <= 16'b0000_0000_0000_0000;
array[22004] <= 16'b0000_0000_0000_0000;
array[22005] <= 16'b0000_0000_0000_0000;
array[22006] <= 16'b0000_0000_0000_0000;
array[22007] <= 16'b0000_0000_0000_0000;
array[22008] <= 16'b0000_0000_0000_0000;
array[22009] <= 16'b0000_0000_0000_0000;
array[22010] <= 16'b0000_0000_0000_0000;
array[22011] <= 16'b0000_0000_0000_0000;
array[22012] <= 16'b0000_0000_0000_0000;
array[22013] <= 16'b0000_0000_0000_0000;
array[22014] <= 16'b0000_0000_0000_0000;
array[22015] <= 16'b0000_0000_0000_0000;
array[22016] <= 16'b0000_0000_0000_0000;
array[22017] <= 16'b0000_0000_0000_0000;
array[22018] <= 16'b0000_0000_0000_0000;
array[22019] <= 16'b0000_0000_0000_0000;
array[22020] <= 16'b0000_0000_0000_0000;
array[22021] <= 16'b0000_0000_0000_0000;
array[22022] <= 16'b0000_0000_0000_0000;
array[22023] <= 16'b0000_0000_0000_0000;
array[22024] <= 16'b0000_0000_0000_0000;
array[22025] <= 16'b0000_0000_0000_0000;
array[22026] <= 16'b0000_0000_0000_0000;
array[22027] <= 16'b0000_0000_0000_0000;
array[22028] <= 16'b0000_0000_0000_0000;
array[22029] <= 16'b0000_0000_0000_0000;
array[22030] <= 16'b0000_0000_0000_0000;
array[22031] <= 16'b0000_0000_0000_0000;
array[22032] <= 16'b0000_0000_0000_0000;
array[22033] <= 16'b0000_0000_0000_0000;
array[22034] <= 16'b0000_0000_0000_0000;
array[22035] <= 16'b0000_0000_0000_0000;
array[22036] <= 16'b0000_0000_0000_0000;
array[22037] <= 16'b0000_0000_0000_0000;
array[22038] <= 16'b0000_0000_0000_0000;
array[22039] <= 16'b0000_0000_0000_0000;
array[22040] <= 16'b0000_0000_0000_0000;
array[22041] <= 16'b0000_0000_0000_0000;
array[22042] <= 16'b0000_0000_0000_0000;
array[22043] <= 16'b0000_0000_0000_0000;
array[22044] <= 16'b0000_0000_0000_0000;
array[22045] <= 16'b0000_0000_0000_0000;
array[22046] <= 16'b0000_0000_0000_0000;
array[22047] <= 16'b0000_0000_0000_0000;
array[22048] <= 16'b0000_0000_0000_0000;
array[22049] <= 16'b0000_0000_0000_0000;
array[22050] <= 16'b0000_0000_0000_0000;
array[22051] <= 16'b0000_0000_0000_0000;
array[22052] <= 16'b0000_0000_0000_0000;
array[22053] <= 16'b0000_0000_0000_0000;
array[22054] <= 16'b0000_0000_0000_0000;
array[22055] <= 16'b0000_0000_0000_0000;
array[22056] <= 16'b0000_0000_0000_0000;
array[22057] <= 16'b0000_0000_0000_0000;
array[22058] <= 16'b0000_0000_0000_0000;
array[22059] <= 16'b0000_0000_0000_0000;
array[22060] <= 16'b0000_0000_0000_0000;
array[22061] <= 16'b0000_0000_0000_0000;
array[22062] <= 16'b0000_0000_0000_0000;
array[22063] <= 16'b0000_0000_0000_0000;
array[22064] <= 16'b0000_0000_0000_0000;
array[22065] <= 16'b0000_0000_0000_0000;
array[22066] <= 16'b0000_0000_0000_0000;
array[22067] <= 16'b0000_0000_0000_0000;
array[22068] <= 16'b0000_0000_0000_0000;
array[22069] <= 16'b0000_0000_0000_0000;
array[22070] <= 16'b0000_0000_0000_0000;
array[22071] <= 16'b0000_0000_0000_0000;
array[22072] <= 16'b0000_0000_0000_0000;
array[22073] <= 16'b0000_0000_0000_0000;
array[22074] <= 16'b0000_0000_0000_0000;
array[22075] <= 16'b0000_0000_0000_0000;
array[22076] <= 16'b0000_0000_0000_0000;
array[22077] <= 16'b0000_0000_0000_0000;
array[22078] <= 16'b0000_0000_0000_0000;
array[22079] <= 16'b0000_0000_0000_0000;
array[22080] <= 16'b0000_0000_0000_0000;
array[22081] <= 16'b0000_0000_0000_0000;
array[22082] <= 16'b0000_0000_0000_0000;
array[22083] <= 16'b0000_0000_0000_0000;
array[22084] <= 16'b0000_0000_0000_0000;
array[22085] <= 16'b0000_0000_0000_0000;
array[22086] <= 16'b0000_0000_0000_0000;
array[22087] <= 16'b0000_0000_0000_0000;
array[22088] <= 16'b0000_0000_0000_0000;
array[22089] <= 16'b0000_0000_0000_0000;
array[22090] <= 16'b0000_0000_0000_0000;
array[22091] <= 16'b0000_0000_0000_0000;
array[22092] <= 16'b0000_0000_0000_0000;
array[22093] <= 16'b0000_0000_0000_0000;
array[22094] <= 16'b0000_0000_0000_0000;
array[22095] <= 16'b0000_0000_0000_0000;
array[22096] <= 16'b0000_0000_0000_0000;
array[22097] <= 16'b0000_0000_0000_0000;
array[22098] <= 16'b0000_0000_0000_0000;
array[22099] <= 16'b0000_0000_0000_0000;
array[22100] <= 16'b0000_0000_0000_0000;
array[22101] <= 16'b0000_0000_0000_0000;
array[22102] <= 16'b0000_0000_0000_0000;
array[22103] <= 16'b0000_0000_0000_0000;
array[22104] <= 16'b0000_0000_0000_0000;
array[22105] <= 16'b0000_0000_0000_0000;
array[22106] <= 16'b0000_0000_0000_0000;
array[22107] <= 16'b0000_0000_0000_0000;
array[22108] <= 16'b0000_0000_0000_0000;
array[22109] <= 16'b0000_0000_0000_0000;
array[22110] <= 16'b0000_0000_0000_0000;
array[22111] <= 16'b0000_0000_0000_0000;
array[22112] <= 16'b0000_0000_0000_0000;
array[22113] <= 16'b0000_0000_0000_0000;
array[22114] <= 16'b0000_0000_0000_0000;
array[22115] <= 16'b0000_0000_0000_0000;
array[22116] <= 16'b0000_0000_0000_0000;
array[22117] <= 16'b0000_0000_0000_0000;
array[22118] <= 16'b0000_0000_0000_0000;
array[22119] <= 16'b0000_0000_0000_0000;
array[22120] <= 16'b0000_0000_0000_0000;
array[22121] <= 16'b0000_0000_0000_0000;
array[22122] <= 16'b0000_0000_0000_0000;
array[22123] <= 16'b0000_0000_0000_0000;
array[22124] <= 16'b0000_0000_0000_0000;
array[22125] <= 16'b0000_0000_0000_0000;
array[22126] <= 16'b0000_0000_0000_0000;
array[22127] <= 16'b0000_0000_0000_0000;
array[22128] <= 16'b0000_0000_0000_0000;
array[22129] <= 16'b0000_0000_0000_0000;
array[22130] <= 16'b0000_0000_0000_0000;
array[22131] <= 16'b0000_0000_0000_0000;
array[22132] <= 16'b0000_0000_0000_0000;
array[22133] <= 16'b0000_0000_0000_0000;
array[22134] <= 16'b0000_0000_0000_0000;
array[22135] <= 16'b0000_0000_0000_0000;
array[22136] <= 16'b0000_0000_0000_0000;
array[22137] <= 16'b0000_0000_0000_0000;
array[22138] <= 16'b0000_0000_0000_0000;
array[22139] <= 16'b0000_0000_0000_0000;
array[22140] <= 16'b0000_0000_0000_0000;
array[22141] <= 16'b0000_0000_0000_0000;
array[22142] <= 16'b0000_0000_0000_0000;
array[22143] <= 16'b0000_0000_0000_0000;
array[22144] <= 16'b0000_0000_0000_0000;
array[22145] <= 16'b0000_0000_0000_0000;
array[22146] <= 16'b0000_0000_0000_0000;
array[22147] <= 16'b0000_0000_0000_0000;
array[22148] <= 16'b0000_0000_0000_0000;
array[22149] <= 16'b0000_0000_0000_0000;
array[22150] <= 16'b0000_0000_0000_0000;
array[22151] <= 16'b0000_0000_0000_0000;
array[22152] <= 16'b0000_0000_0000_0000;
array[22153] <= 16'b0000_0000_0000_0000;
array[22154] <= 16'b0000_0000_0000_0000;
array[22155] <= 16'b0000_0000_0000_0000;
array[22156] <= 16'b0000_0000_0000_0000;
array[22157] <= 16'b0000_0000_0000_0000;
array[22158] <= 16'b0000_0000_0000_0000;
array[22159] <= 16'b0000_0000_0000_0000;
array[22160] <= 16'b0000_0000_0000_0000;
array[22161] <= 16'b0000_0000_0000_0000;
array[22162] <= 16'b0000_0000_0000_0000;
array[22163] <= 16'b0000_0000_0000_0000;
array[22164] <= 16'b0000_0000_0000_0000;
array[22165] <= 16'b0000_0000_0000_0000;
array[22166] <= 16'b0000_0000_0000_0000;
array[22167] <= 16'b0000_0000_0000_0000;
array[22168] <= 16'b0000_0000_0000_0000;
array[22169] <= 16'b0000_0000_0000_0000;
array[22170] <= 16'b0000_0000_0000_0000;
array[22171] <= 16'b0000_0000_0000_0000;
array[22172] <= 16'b0000_0000_0000_0000;
array[22173] <= 16'b0000_0000_0000_0000;
array[22174] <= 16'b0000_0000_0000_0000;
array[22175] <= 16'b0000_0000_0000_0000;
array[22176] <= 16'b0000_0000_0000_0000;
array[22177] <= 16'b0000_0000_0000_0000;
array[22178] <= 16'b0000_0000_0000_0000;
array[22179] <= 16'b0000_0000_0000_0000;
array[22180] <= 16'b0000_0000_0000_0000;
array[22181] <= 16'b0000_0000_0000_0000;
array[22182] <= 16'b0000_0000_0000_0000;
array[22183] <= 16'b0000_0000_0000_0000;
array[22184] <= 16'b0000_0000_0000_0000;
array[22185] <= 16'b0000_0000_0000_0000;
array[22186] <= 16'b0000_0000_0000_0000;
array[22187] <= 16'b0000_0000_0000_0000;
array[22188] <= 16'b0000_0000_0000_0000;
array[22189] <= 16'b0000_0000_0000_0000;
array[22190] <= 16'b0000_0000_0000_0000;
array[22191] <= 16'b0000_0000_0000_0000;
array[22192] <= 16'b0000_0000_0000_0000;
array[22193] <= 16'b0000_0000_0000_0000;
array[22194] <= 16'b0000_0000_0000_0000;
array[22195] <= 16'b0000_0000_0000_0000;
array[22196] <= 16'b0000_0000_0000_0000;
array[22197] <= 16'b0000_0000_0000_0000;
array[22198] <= 16'b0000_0000_0000_0000;
array[22199] <= 16'b0000_0000_0000_0000;
array[22200] <= 16'b0000_0000_0000_0000;
array[22201] <= 16'b0000_0000_0000_0000;
array[22202] <= 16'b0000_0000_0000_0000;
array[22203] <= 16'b0000_0000_0000_0000;
array[22204] <= 16'b0000_0000_0000_0000;
array[22205] <= 16'b0000_0000_0000_0000;
array[22206] <= 16'b0000_0000_0000_0000;
array[22207] <= 16'b0000_0000_0000_0000;
array[22208] <= 16'b0000_0000_0000_0000;
array[22209] <= 16'b0000_0000_0000_0000;
array[22210] <= 16'b0000_0000_0000_0000;
array[22211] <= 16'b0000_0000_0000_0000;
array[22212] <= 16'b0000_0000_0000_0000;
array[22213] <= 16'b0000_0000_0000_0000;
array[22214] <= 16'b0000_0000_0000_0000;
array[22215] <= 16'b0000_0000_0000_0000;
array[22216] <= 16'b0000_0000_0000_0000;
array[22217] <= 16'b0000_0000_0000_0000;
array[22218] <= 16'b0000_0000_0000_0000;
array[22219] <= 16'b0000_0000_0000_0000;
array[22220] <= 16'b0000_0000_0000_0000;
array[22221] <= 16'b0000_0000_0000_0000;
array[22222] <= 16'b0000_0000_0000_0000;
array[22223] <= 16'b0000_0000_0000_0000;
array[22224] <= 16'b0000_0000_0000_0000;
array[22225] <= 16'b0000_0000_0000_0000;
array[22226] <= 16'b0000_0000_0000_0000;
array[22227] <= 16'b0000_0000_0000_0000;
array[22228] <= 16'b0000_0000_0000_0000;
array[22229] <= 16'b0000_0000_0000_0000;
array[22230] <= 16'b0000_0000_0000_0000;
array[22231] <= 16'b0000_0000_0000_0000;
array[22232] <= 16'b0000_0000_0000_0000;
array[22233] <= 16'b0000_0000_0000_0000;
array[22234] <= 16'b0000_0000_0000_0000;
array[22235] <= 16'b0000_0000_0000_0000;
array[22236] <= 16'b0000_0000_0000_0000;
array[22237] <= 16'b0000_0000_0000_0000;
array[22238] <= 16'b0000_0000_0000_0000;
array[22239] <= 16'b0000_0000_0000_0000;
array[22240] <= 16'b0000_0000_0000_0000;
array[22241] <= 16'b0000_0000_0000_0000;
array[22242] <= 16'b0000_0000_0000_0000;
array[22243] <= 16'b0000_0000_0000_0000;
array[22244] <= 16'b0000_0000_0000_0000;
array[22245] <= 16'b0000_0000_0000_0000;
array[22246] <= 16'b0000_0000_0000_0000;
array[22247] <= 16'b0000_0000_0000_0000;
array[22248] <= 16'b0000_0000_0000_0000;
array[22249] <= 16'b0000_0000_0000_0000;
array[22250] <= 16'b0000_0000_0000_0000;
array[22251] <= 16'b0000_0000_0000_0000;
array[22252] <= 16'b0000_0000_0000_0000;
array[22253] <= 16'b0000_0000_0000_0000;
array[22254] <= 16'b0000_0000_0000_0000;
array[22255] <= 16'b0000_0000_0000_0000;
array[22256] <= 16'b0000_0000_0000_0000;
array[22257] <= 16'b0000_0000_0000_0000;
array[22258] <= 16'b0000_0000_0000_0000;
array[22259] <= 16'b0000_0000_0000_0000;
array[22260] <= 16'b0000_0000_0000_0000;
array[22261] <= 16'b0000_0000_0000_0000;
array[22262] <= 16'b0000_0000_0000_0000;
array[22263] <= 16'b0000_0000_0000_0000;
array[22264] <= 16'b0000_0000_0000_0000;
array[22265] <= 16'b0000_0000_0000_0000;
array[22266] <= 16'b0000_0000_0000_0000;
array[22267] <= 16'b0000_0000_0000_0000;
array[22268] <= 16'b0000_0000_0000_0000;
array[22269] <= 16'b0000_0000_0000_0000;
array[22270] <= 16'b0000_0000_0000_0000;
array[22271] <= 16'b0000_0000_0000_0000;
array[22272] <= 16'b0000_0000_0000_0000;
array[22273] <= 16'b0000_0000_0000_0000;
array[22274] <= 16'b0000_0000_0000_0000;
array[22275] <= 16'b0000_0000_0000_0000;
array[22276] <= 16'b0000_0000_0000_0000;
array[22277] <= 16'b0000_0000_0000_0000;
array[22278] <= 16'b0000_0000_0000_0000;
array[22279] <= 16'b0000_0000_0000_0000;
array[22280] <= 16'b0000_0000_0000_0000;
array[22281] <= 16'b0000_0000_0000_0000;
array[22282] <= 16'b0000_0000_0000_0000;
array[22283] <= 16'b0000_0000_0000_0000;
array[22284] <= 16'b0000_0000_0000_0000;
array[22285] <= 16'b0000_0000_0000_0000;
array[22286] <= 16'b0000_0000_0000_0000;
array[22287] <= 16'b0000_0000_0000_0000;
array[22288] <= 16'b0000_0000_0000_0000;
array[22289] <= 16'b0000_0000_0000_0000;
array[22290] <= 16'b0000_0000_0000_0000;
array[22291] <= 16'b0000_0000_0000_0000;
array[22292] <= 16'b0000_0000_0000_0000;
array[22293] <= 16'b0000_0000_0000_0000;
array[22294] <= 16'b0000_0000_0000_0000;
array[22295] <= 16'b0000_0000_0000_0000;
array[22296] <= 16'b0000_0000_0000_0000;
array[22297] <= 16'b0000_0000_0000_0000;
array[22298] <= 16'b0000_0000_0000_0000;
array[22299] <= 16'b0000_0000_0000_0000;
array[22300] <= 16'b0000_0000_0000_0000;
array[22301] <= 16'b0000_0000_0000_0000;
array[22302] <= 16'b0000_0000_0000_0000;
array[22303] <= 16'b0000_0000_0000_0000;
array[22304] <= 16'b0000_0000_0000_0000;
array[22305] <= 16'b0000_0000_0000_0000;
array[22306] <= 16'b0000_0000_0000_0000;
array[22307] <= 16'b0000_0000_0000_0000;
array[22308] <= 16'b0000_0000_0000_0000;
array[22309] <= 16'b0000_0000_0000_0000;
array[22310] <= 16'b0000_0000_0000_0000;
array[22311] <= 16'b0000_0000_0000_0000;
array[22312] <= 16'b0000_0000_0000_0000;
array[22313] <= 16'b0000_0000_0000_0000;
array[22314] <= 16'b0000_0000_0000_0000;
array[22315] <= 16'b0000_0000_0000_0000;
array[22316] <= 16'b0000_0000_0000_0000;
array[22317] <= 16'b0000_0000_0000_0000;
array[22318] <= 16'b0000_0000_0000_0000;
array[22319] <= 16'b0000_0000_0000_0000;
array[22320] <= 16'b0000_0000_0000_0000;
array[22321] <= 16'b0000_0000_0000_0000;
array[22322] <= 16'b0000_0000_0000_0000;
array[22323] <= 16'b0000_0000_0000_0000;
array[22324] <= 16'b0000_0000_0000_0000;
array[22325] <= 16'b0000_0000_0000_0000;
array[22326] <= 16'b0000_0000_0000_0000;
array[22327] <= 16'b0000_0000_0000_0000;
array[22328] <= 16'b0000_0000_0000_0000;
array[22329] <= 16'b0000_0000_0000_0000;
array[22330] <= 16'b0000_0000_0000_0000;
array[22331] <= 16'b0000_0000_0000_0000;
array[22332] <= 16'b0000_0000_0000_0000;
array[22333] <= 16'b0000_0000_0000_0000;
array[22334] <= 16'b0000_0000_0000_0000;
array[22335] <= 16'b0000_0000_0000_0000;
array[22336] <= 16'b0000_0000_0000_0000;
array[22337] <= 16'b0000_0000_0000_0000;
array[22338] <= 16'b0000_0000_0000_0000;
array[22339] <= 16'b0000_0000_0000_0000;
array[22340] <= 16'b0000_0000_0000_0000;
array[22341] <= 16'b0000_0000_0000_0000;
array[22342] <= 16'b0000_0000_0000_0000;
array[22343] <= 16'b0000_0000_0000_0000;
array[22344] <= 16'b0000_0000_0000_0000;
array[22345] <= 16'b0000_0000_0000_0000;
array[22346] <= 16'b0000_0000_0000_0000;
array[22347] <= 16'b0000_0000_0000_0000;
array[22348] <= 16'b0000_0000_0000_0000;
array[22349] <= 16'b0000_0000_0000_0000;
array[22350] <= 16'b0000_0000_0000_0000;
array[22351] <= 16'b0000_0000_0000_0000;
array[22352] <= 16'b0000_0000_0000_0000;
array[22353] <= 16'b0000_0000_0000_0000;
array[22354] <= 16'b0000_0000_0000_0000;
array[22355] <= 16'b0000_0000_0000_0000;
array[22356] <= 16'b0000_0000_0000_0000;
array[22357] <= 16'b0000_0000_0000_0000;
array[22358] <= 16'b0000_0000_0000_0000;
array[22359] <= 16'b0000_0000_0000_0000;
array[22360] <= 16'b0000_0000_0000_0000;
array[22361] <= 16'b0000_0000_0000_0000;
array[22362] <= 16'b0000_0000_0000_0000;
array[22363] <= 16'b0000_0000_0000_0000;
array[22364] <= 16'b0000_0000_0000_0000;
array[22365] <= 16'b0000_0000_0000_0000;
array[22366] <= 16'b0000_0000_0000_0000;
array[22367] <= 16'b0000_0000_0000_0000;
array[22368] <= 16'b0000_0000_0000_0000;
array[22369] <= 16'b0000_0000_0000_0000;
array[22370] <= 16'b0000_0000_0000_0000;
array[22371] <= 16'b0000_0000_0000_0000;
array[22372] <= 16'b0000_0000_0000_0000;
array[22373] <= 16'b0000_0000_0000_0000;
array[22374] <= 16'b0000_0000_0000_0000;
array[22375] <= 16'b0000_0000_0000_0000;
array[22376] <= 16'b0000_0000_0000_0000;
array[22377] <= 16'b0000_0000_0000_0000;
array[22378] <= 16'b0000_0000_0000_0000;
array[22379] <= 16'b0000_0000_0000_0000;
array[22380] <= 16'b0000_0000_0000_0000;
array[22381] <= 16'b0000_0000_0000_0000;
array[22382] <= 16'b0000_0000_0000_0000;
array[22383] <= 16'b0000_0000_0000_0000;
array[22384] <= 16'b0000_0000_0000_0000;
array[22385] <= 16'b0000_0000_0000_0000;
array[22386] <= 16'b0000_0000_0000_0000;
array[22387] <= 16'b0000_0000_0000_0000;
array[22388] <= 16'b0000_0000_0000_0000;
array[22389] <= 16'b0000_0000_0000_0000;
array[22390] <= 16'b0000_0000_0000_0000;
array[22391] <= 16'b0000_0000_0000_0000;
array[22392] <= 16'b0000_0000_0000_0000;
array[22393] <= 16'b0000_0000_0000_0000;
array[22394] <= 16'b0000_0000_0000_0000;
array[22395] <= 16'b0000_0000_0000_0000;
array[22396] <= 16'b0000_0000_0000_0000;
array[22397] <= 16'b0000_0000_0000_0000;
array[22398] <= 16'b0000_0000_0000_0000;
array[22399] <= 16'b0000_0000_0000_0000;
array[22400] <= 16'b0000_0000_0000_0000;
array[22401] <= 16'b0000_0000_0000_0000;
array[22402] <= 16'b0000_0000_0000_0000;
array[22403] <= 16'b0000_0000_0000_0000;
array[22404] <= 16'b0000_0000_0000_0000;
array[22405] <= 16'b0000_0000_0000_0000;
array[22406] <= 16'b0000_0000_0000_0000;
array[22407] <= 16'b0000_0000_0000_0000;
array[22408] <= 16'b0000_0000_0000_0000;
array[22409] <= 16'b0000_0000_0000_0000;
array[22410] <= 16'b0000_0000_0000_0000;
array[22411] <= 16'b0000_0000_0000_0000;
array[22412] <= 16'b0000_0000_0000_0000;
array[22413] <= 16'b0000_0000_0000_0000;
array[22414] <= 16'b0000_0000_0000_0000;
array[22415] <= 16'b0000_0000_0000_0000;
array[22416] <= 16'b0000_0000_0000_0000;
array[22417] <= 16'b0000_0000_0000_0000;
array[22418] <= 16'b0000_0000_0000_0000;
array[22419] <= 16'b0000_0000_0000_0000;
array[22420] <= 16'b0000_0000_0000_0000;
array[22421] <= 16'b0000_0000_0000_0000;
array[22422] <= 16'b0000_0000_0000_0000;
array[22423] <= 16'b0000_0000_0000_0000;
array[22424] <= 16'b0000_0000_0000_0000;
array[22425] <= 16'b0000_0000_0000_0000;
array[22426] <= 16'b0000_0000_0000_0000;
array[22427] <= 16'b0000_0000_0000_0000;
array[22428] <= 16'b0000_0000_0000_0000;
array[22429] <= 16'b0000_0000_0000_0000;
array[22430] <= 16'b0000_0000_0000_0000;
array[22431] <= 16'b0000_0000_0000_0000;
array[22432] <= 16'b0000_0000_0000_0000;
array[22433] <= 16'b0000_0000_0000_0000;
array[22434] <= 16'b0000_0000_0000_0000;
array[22435] <= 16'b0000_0000_0000_0000;
array[22436] <= 16'b0000_0000_0000_0000;
array[22437] <= 16'b0000_0000_0000_0000;
array[22438] <= 16'b0000_0000_0000_0000;
array[22439] <= 16'b0000_0000_0000_0000;
array[22440] <= 16'b0000_0000_0000_0000;
array[22441] <= 16'b0000_0000_0000_0000;
array[22442] <= 16'b0000_0000_0000_0000;
array[22443] <= 16'b0000_0000_0000_0000;
array[22444] <= 16'b0000_0000_0000_0000;
array[22445] <= 16'b0000_0000_0000_0000;
array[22446] <= 16'b0000_0000_0000_0000;
array[22447] <= 16'b0000_0000_0000_0000;
array[22448] <= 16'b0000_0000_0000_0000;
array[22449] <= 16'b0000_0000_0000_0000;
array[22450] <= 16'b0000_0000_0000_0000;
array[22451] <= 16'b0000_0000_0000_0000;
array[22452] <= 16'b0000_0000_0000_0000;
array[22453] <= 16'b0000_0000_0000_0000;
array[22454] <= 16'b0000_0000_0000_0000;
array[22455] <= 16'b0000_0000_0000_0000;
array[22456] <= 16'b0000_0000_0000_0000;
array[22457] <= 16'b0000_0000_0000_0000;
array[22458] <= 16'b0000_0000_0000_0000;
array[22459] <= 16'b0000_0000_0000_0000;
array[22460] <= 16'b0000_0000_0000_0000;
array[22461] <= 16'b0000_0000_0000_0000;
array[22462] <= 16'b0000_0000_0000_0000;
array[22463] <= 16'b0000_0000_0000_0000;
array[22464] <= 16'b0000_0000_0000_0000;
array[22465] <= 16'b0000_0000_0000_0000;
array[22466] <= 16'b0000_0000_0000_0000;
array[22467] <= 16'b0000_0000_0000_0000;
array[22468] <= 16'b0000_0000_0000_0000;
array[22469] <= 16'b0000_0000_0000_0000;
array[22470] <= 16'b0000_0000_0000_0000;
array[22471] <= 16'b0000_0000_0000_0000;
array[22472] <= 16'b0000_0000_0000_0000;
array[22473] <= 16'b0000_0000_0000_0000;
array[22474] <= 16'b0000_0000_0000_0000;
array[22475] <= 16'b0000_0000_0000_0000;
array[22476] <= 16'b0000_0000_0000_0000;
array[22477] <= 16'b0000_0000_0000_0000;
array[22478] <= 16'b0000_0000_0000_0000;
array[22479] <= 16'b0000_0000_0000_0000;
array[22480] <= 16'b0000_0000_0000_0000;
array[22481] <= 16'b0000_0000_0000_0000;
array[22482] <= 16'b0000_0000_0000_0000;
array[22483] <= 16'b0000_0000_0000_0000;
array[22484] <= 16'b0000_0000_0000_0000;
array[22485] <= 16'b0000_0000_0000_0000;
array[22486] <= 16'b0000_0000_0000_0000;
array[22487] <= 16'b0000_0000_0000_0000;
array[22488] <= 16'b0000_0000_0000_0000;
array[22489] <= 16'b0000_0000_0000_0000;
array[22490] <= 16'b0000_0000_0000_0000;
array[22491] <= 16'b0000_0000_0000_0000;
array[22492] <= 16'b0000_0000_0000_0000;
array[22493] <= 16'b0000_0000_0000_0000;
array[22494] <= 16'b0000_0000_0000_0000;
array[22495] <= 16'b0000_0000_0000_0000;
array[22496] <= 16'b0000_0000_0000_0000;
array[22497] <= 16'b0000_0000_0000_0000;
array[22498] <= 16'b0000_0000_0000_0000;
array[22499] <= 16'b0000_0000_0000_0000;
array[22500] <= 16'b0000_0000_0000_0000;
array[22501] <= 16'b0000_0000_0000_0000;
array[22502] <= 16'b0000_0000_0000_0000;
array[22503] <= 16'b0000_0000_0000_0000;
array[22504] <= 16'b0000_0000_0000_0000;
array[22505] <= 16'b0000_0000_0000_0000;
array[22506] <= 16'b0000_0000_0000_0000;
array[22507] <= 16'b0000_0000_0000_0000;
array[22508] <= 16'b0000_0000_0000_0000;
array[22509] <= 16'b0000_0000_0000_0000;
array[22510] <= 16'b0000_0000_0000_0000;
array[22511] <= 16'b0000_0000_0000_0000;
array[22512] <= 16'b0000_0000_0000_0000;
array[22513] <= 16'b0000_0000_0000_0000;
array[22514] <= 16'b0000_0000_0000_0000;
array[22515] <= 16'b0000_0000_0000_0000;
array[22516] <= 16'b0000_0000_0000_0000;
array[22517] <= 16'b0000_0000_0000_0000;
array[22518] <= 16'b0000_0000_0000_0000;
array[22519] <= 16'b0000_0000_0000_0000;
array[22520] <= 16'b0000_0000_0000_0000;
array[22521] <= 16'b0000_0000_0000_0000;
array[22522] <= 16'b0000_0000_0000_0000;
array[22523] <= 16'b0000_0000_0000_0000;
array[22524] <= 16'b0000_0000_0000_0000;
array[22525] <= 16'b0000_0000_0000_0000;
array[22526] <= 16'b0000_0000_0000_0000;
array[22527] <= 16'b0000_0000_0000_0000;
array[22528] <= 16'b0000_0000_0000_0000;
array[22529] <= 16'b0000_0000_0000_0000;
array[22530] <= 16'b0000_0000_0000_0000;
array[22531] <= 16'b0000_0000_0000_0000;
array[22532] <= 16'b0000_0000_0000_0000;
array[22533] <= 16'b0000_0000_0000_0000;
array[22534] <= 16'b0000_0000_0000_0000;
array[22535] <= 16'b0000_0000_0000_0000;
array[22536] <= 16'b0000_0000_0000_0000;
array[22537] <= 16'b0000_0000_0000_0000;
array[22538] <= 16'b0000_0000_0000_0000;
array[22539] <= 16'b0000_0000_0000_0000;
array[22540] <= 16'b0000_0000_0000_0000;
array[22541] <= 16'b0000_0000_0000_0000;
array[22542] <= 16'b0000_0000_0000_0000;
array[22543] <= 16'b0000_0000_0000_0000;
array[22544] <= 16'b0000_0000_0000_0000;
array[22545] <= 16'b0000_0000_0000_0000;
array[22546] <= 16'b0000_0000_0000_0000;
array[22547] <= 16'b0000_0000_0000_0000;
array[22548] <= 16'b0000_0000_0000_0000;
array[22549] <= 16'b0000_0000_0000_0000;
array[22550] <= 16'b0000_0000_0000_0000;
array[22551] <= 16'b0000_0000_0000_0000;
array[22552] <= 16'b0000_0000_0000_0000;
array[22553] <= 16'b0000_0000_0000_0000;
array[22554] <= 16'b0000_0000_0000_0000;
array[22555] <= 16'b0000_0000_0000_0000;
array[22556] <= 16'b0000_0000_0000_0000;
array[22557] <= 16'b0000_0000_0000_0000;
array[22558] <= 16'b0000_0000_0000_0000;
array[22559] <= 16'b0000_0000_0000_0000;
array[22560] <= 16'b0000_0000_0000_0000;
array[22561] <= 16'b0000_0000_0000_0000;
array[22562] <= 16'b0000_0000_0000_0000;
array[22563] <= 16'b0000_0000_0000_0000;
array[22564] <= 16'b0000_0000_0000_0000;
array[22565] <= 16'b0000_0000_0000_0000;
array[22566] <= 16'b0000_0000_0000_0000;
array[22567] <= 16'b0000_0000_0000_0000;
array[22568] <= 16'b0000_0000_0000_0000;
array[22569] <= 16'b0000_0000_0000_0000;
array[22570] <= 16'b0000_0000_0000_0000;
array[22571] <= 16'b0000_0000_0000_0000;
array[22572] <= 16'b0000_0000_0000_0000;
array[22573] <= 16'b0000_0000_0000_0000;
array[22574] <= 16'b0000_0000_0000_0000;
array[22575] <= 16'b0000_0000_0000_0000;
array[22576] <= 16'b0000_0000_0000_0000;
array[22577] <= 16'b0000_0000_0000_0000;
array[22578] <= 16'b0000_0000_0000_0000;
array[22579] <= 16'b0000_0000_0000_0000;
array[22580] <= 16'b0000_0000_0000_0000;
array[22581] <= 16'b0000_0000_0000_0000;
array[22582] <= 16'b0000_0000_0000_0000;
array[22583] <= 16'b0000_0000_0000_0000;
array[22584] <= 16'b0000_0000_0000_0000;
array[22585] <= 16'b0000_0000_0000_0000;
array[22586] <= 16'b0000_0000_0000_0000;
array[22587] <= 16'b0000_0000_0000_0000;
array[22588] <= 16'b0000_0000_0000_0000;
array[22589] <= 16'b0000_0000_0000_0000;
array[22590] <= 16'b0000_0000_0000_0000;
array[22591] <= 16'b0000_0000_0000_0000;
array[22592] <= 16'b0000_0000_0000_0000;
array[22593] <= 16'b0000_0000_0000_0000;
array[22594] <= 16'b0000_0000_0000_0000;
array[22595] <= 16'b0000_0000_0000_0000;
array[22596] <= 16'b0000_0000_0000_0000;
array[22597] <= 16'b0000_0000_0000_0000;
array[22598] <= 16'b0000_0000_0000_0000;
array[22599] <= 16'b0000_0000_0000_0000;
array[22600] <= 16'b0000_0000_0000_0000;
array[22601] <= 16'b0000_0000_0000_0000;
array[22602] <= 16'b0000_0000_0000_0000;
array[22603] <= 16'b0000_0000_0000_0000;
array[22604] <= 16'b0000_0000_0000_0000;
array[22605] <= 16'b0000_0000_0000_0000;
array[22606] <= 16'b0000_0000_0000_0000;
array[22607] <= 16'b0000_0000_0000_0000;
array[22608] <= 16'b0000_0000_0000_0000;
array[22609] <= 16'b0000_0000_0000_0000;
array[22610] <= 16'b0000_0000_0000_0000;
array[22611] <= 16'b0000_0000_0000_0000;
array[22612] <= 16'b0000_0000_0000_0000;
array[22613] <= 16'b0000_0000_0000_0000;
array[22614] <= 16'b0000_0000_0000_0000;
array[22615] <= 16'b0000_0000_0000_0000;
array[22616] <= 16'b0000_0000_0000_0000;
array[22617] <= 16'b0000_0000_0000_0000;
array[22618] <= 16'b0000_0000_0000_0000;
array[22619] <= 16'b0000_0000_0000_0000;
array[22620] <= 16'b0000_0000_0000_0000;
array[22621] <= 16'b0000_0000_0000_0000;
array[22622] <= 16'b0000_0000_0000_0000;
array[22623] <= 16'b0000_0000_0000_0000;
array[22624] <= 16'b0000_0000_0000_0000;
array[22625] <= 16'b0000_0000_0000_0000;
array[22626] <= 16'b0000_0000_0000_0000;
array[22627] <= 16'b0000_0000_0000_0000;
array[22628] <= 16'b0000_0000_0000_0000;
array[22629] <= 16'b0000_0000_0000_0000;
array[22630] <= 16'b0000_0000_0000_0000;
array[22631] <= 16'b0000_0000_0000_0000;
array[22632] <= 16'b0000_0000_0000_0000;
array[22633] <= 16'b0000_0000_0000_0000;
array[22634] <= 16'b0000_0000_0000_0000;
array[22635] <= 16'b0000_0000_0000_0000;
array[22636] <= 16'b0000_0000_0000_0000;
array[22637] <= 16'b0000_0000_0000_0000;
array[22638] <= 16'b0000_0000_0000_0000;
array[22639] <= 16'b0000_0000_0000_0000;
array[22640] <= 16'b0000_0000_0000_0000;
array[22641] <= 16'b0000_0000_0000_0000;
array[22642] <= 16'b0000_0000_0000_0000;
array[22643] <= 16'b0000_0000_0000_0000;
array[22644] <= 16'b0000_0000_0000_0000;
array[22645] <= 16'b0000_0000_0000_0000;
array[22646] <= 16'b0000_0000_0000_0000;
array[22647] <= 16'b0000_0000_0000_0000;
array[22648] <= 16'b0000_0000_0000_0000;
array[22649] <= 16'b0000_0000_0000_0000;
array[22650] <= 16'b0000_0000_0000_0000;
array[22651] <= 16'b0000_0000_0000_0000;
array[22652] <= 16'b0000_0000_0000_0000;
array[22653] <= 16'b0000_0000_0000_0000;
array[22654] <= 16'b0000_0000_0000_0000;
array[22655] <= 16'b0000_0000_0000_0000;
array[22656] <= 16'b0000_0000_0000_0000;
array[22657] <= 16'b0000_0000_0000_0000;
array[22658] <= 16'b0000_0000_0000_0000;
array[22659] <= 16'b0000_0000_0000_0000;
array[22660] <= 16'b0000_0000_0000_0000;
array[22661] <= 16'b0000_0000_0000_0000;
array[22662] <= 16'b0000_0000_0000_0000;
array[22663] <= 16'b0000_0000_0000_0000;
array[22664] <= 16'b0000_0000_0000_0000;
array[22665] <= 16'b0000_0000_0000_0000;
array[22666] <= 16'b0000_0000_0000_0000;
array[22667] <= 16'b0000_0000_0000_0000;
array[22668] <= 16'b0000_0000_0000_0000;
array[22669] <= 16'b0000_0000_0000_0000;
array[22670] <= 16'b0000_0000_0000_0000;
array[22671] <= 16'b0000_0000_0000_0000;
array[22672] <= 16'b0000_0000_0000_0000;
array[22673] <= 16'b0000_0000_0000_0000;
array[22674] <= 16'b0000_0000_0000_0000;
array[22675] <= 16'b0000_0000_0000_0000;
array[22676] <= 16'b0000_0000_0000_0000;
array[22677] <= 16'b0000_0000_0000_0000;
array[22678] <= 16'b0000_0000_0000_0000;
array[22679] <= 16'b0000_0000_0000_0000;
array[22680] <= 16'b0000_0000_0000_0000;
array[22681] <= 16'b0000_0000_0000_0000;
array[22682] <= 16'b0000_0000_0000_0000;
array[22683] <= 16'b0000_0000_0000_0000;
array[22684] <= 16'b0000_0000_0000_0000;
array[22685] <= 16'b0000_0000_0000_0000;
array[22686] <= 16'b0000_0000_0000_0000;
array[22687] <= 16'b0000_0000_0000_0000;
array[22688] <= 16'b0000_0000_0000_0000;
array[22689] <= 16'b0000_0000_0000_0000;
array[22690] <= 16'b0000_0000_0000_0000;
array[22691] <= 16'b0000_0000_0000_0000;
array[22692] <= 16'b0000_0000_0000_0000;
array[22693] <= 16'b0000_0000_0000_0000;
array[22694] <= 16'b0000_0000_0000_0000;
array[22695] <= 16'b0000_0000_0000_0000;
array[22696] <= 16'b0000_0000_0000_0000;
array[22697] <= 16'b0000_0000_0000_0000;
array[22698] <= 16'b0000_0000_0000_0000;
array[22699] <= 16'b0000_0000_0000_0000;
array[22700] <= 16'b0000_0000_0000_0000;
array[22701] <= 16'b0000_0000_0000_0000;
array[22702] <= 16'b0000_0000_0000_0000;
array[22703] <= 16'b0000_0000_0000_0000;
array[22704] <= 16'b0000_0000_0000_0000;
array[22705] <= 16'b0000_0000_0000_0000;
array[22706] <= 16'b0000_0000_0000_0000;
array[22707] <= 16'b0000_0000_0000_0000;
array[22708] <= 16'b0000_0000_0000_0000;
array[22709] <= 16'b0000_0000_0000_0000;
array[22710] <= 16'b0000_0000_0000_0000;
array[22711] <= 16'b0000_0000_0000_0000;
array[22712] <= 16'b0000_0000_0000_0000;
array[22713] <= 16'b0000_0000_0000_0000;
array[22714] <= 16'b0000_0000_0000_0000;
array[22715] <= 16'b0000_0000_0000_0000;
array[22716] <= 16'b0000_0000_0000_0000;
array[22717] <= 16'b0000_0000_0000_0000;
array[22718] <= 16'b0000_0000_0000_0000;
array[22719] <= 16'b0000_0000_0000_0000;
array[22720] <= 16'b0000_0000_0000_0000;
array[22721] <= 16'b0000_0000_0000_0000;
array[22722] <= 16'b0000_0000_0000_0000;
array[22723] <= 16'b0000_0000_0000_0000;
array[22724] <= 16'b0000_0000_0000_0000;
array[22725] <= 16'b0000_0000_0000_0000;
array[22726] <= 16'b0000_0000_0000_0000;
array[22727] <= 16'b0000_0000_0000_0000;
array[22728] <= 16'b0000_0000_0000_0000;
array[22729] <= 16'b0000_0000_0000_0000;
array[22730] <= 16'b0000_0000_0000_0000;
array[22731] <= 16'b0000_0000_0000_0000;
array[22732] <= 16'b0000_0000_0000_0000;
array[22733] <= 16'b0000_0000_0000_0000;
array[22734] <= 16'b0000_0000_0000_0000;
array[22735] <= 16'b0000_0000_0000_0000;
array[22736] <= 16'b0000_0000_0000_0000;
array[22737] <= 16'b0000_0000_0000_0000;
array[22738] <= 16'b0000_0000_0000_0000;
array[22739] <= 16'b0000_0000_0000_0000;
array[22740] <= 16'b0000_0000_0000_0000;
array[22741] <= 16'b0000_0000_0000_0000;
array[22742] <= 16'b0000_0000_0000_0000;
array[22743] <= 16'b0000_0000_0000_0000;
array[22744] <= 16'b0000_0000_0000_0000;
array[22745] <= 16'b0000_0000_0000_0000;
array[22746] <= 16'b0000_0000_0000_0000;
array[22747] <= 16'b0000_0000_0000_0000;
array[22748] <= 16'b0000_0000_0000_0000;
array[22749] <= 16'b0000_0000_0000_0000;
array[22750] <= 16'b0000_0000_0000_0000;
array[22751] <= 16'b0000_0000_0000_0000;
array[22752] <= 16'b0000_0000_0000_0000;
array[22753] <= 16'b0000_0000_0000_0000;
array[22754] <= 16'b0000_0000_0000_0000;
array[22755] <= 16'b0000_0000_0000_0000;
array[22756] <= 16'b0000_0000_0000_0000;
array[22757] <= 16'b0000_0000_0000_0000;
array[22758] <= 16'b0000_0000_0000_0000;
array[22759] <= 16'b0000_0000_0000_0000;
array[22760] <= 16'b0000_0000_0000_0000;
array[22761] <= 16'b0000_0000_0000_0000;
array[22762] <= 16'b0000_0000_0000_0000;
array[22763] <= 16'b0000_0000_0000_0000;
array[22764] <= 16'b0000_0000_0000_0000;
array[22765] <= 16'b0000_0000_0000_0000;
array[22766] <= 16'b0000_0000_0000_0000;
array[22767] <= 16'b0000_0000_0000_0000;
array[22768] <= 16'b0000_0000_0000_0000;
array[22769] <= 16'b0000_0000_0000_0000;
array[22770] <= 16'b0000_0000_0000_0000;
array[22771] <= 16'b0000_0000_0000_0000;
array[22772] <= 16'b0000_0000_0000_0000;
array[22773] <= 16'b0000_0000_0000_0000;
array[22774] <= 16'b0000_0000_0000_0000;
array[22775] <= 16'b0000_0000_0000_0000;
array[22776] <= 16'b0000_0000_0000_0000;
array[22777] <= 16'b0000_0000_0000_0000;
array[22778] <= 16'b0000_0000_0000_0000;
array[22779] <= 16'b0000_0000_0000_0000;
array[22780] <= 16'b0000_0000_0000_0000;
array[22781] <= 16'b0000_0000_0000_0000;
array[22782] <= 16'b0000_0000_0000_0000;
array[22783] <= 16'b0000_0000_0000_0000;
array[22784] <= 16'b0000_0000_0000_0000;
array[22785] <= 16'b0000_0000_0000_0000;
array[22786] <= 16'b0000_0000_0000_0000;
array[22787] <= 16'b0000_0000_0000_0000;
array[22788] <= 16'b0000_0000_0000_0000;
array[22789] <= 16'b0000_0000_0000_0000;
array[22790] <= 16'b0000_0000_0000_0000;
array[22791] <= 16'b0000_0000_0000_0000;
array[22792] <= 16'b0000_0000_0000_0000;
array[22793] <= 16'b0000_0000_0000_0000;
array[22794] <= 16'b0000_0000_0000_0000;
array[22795] <= 16'b0000_0000_0000_0000;
array[22796] <= 16'b0000_0000_0000_0000;
array[22797] <= 16'b0000_0000_0000_0000;
array[22798] <= 16'b0000_0000_0000_0000;
array[22799] <= 16'b0000_0000_0000_0000;
array[22800] <= 16'b0000_0000_0000_0000;
array[22801] <= 16'b0000_0000_0000_0000;
array[22802] <= 16'b0000_0000_0000_0000;
array[22803] <= 16'b0000_0000_0000_0000;
array[22804] <= 16'b0000_0000_0000_0000;
array[22805] <= 16'b0000_0000_0000_0000;
array[22806] <= 16'b0000_0000_0000_0000;
array[22807] <= 16'b0000_0000_0000_0000;
array[22808] <= 16'b0000_0000_0000_0000;
array[22809] <= 16'b0000_0000_0000_0000;
array[22810] <= 16'b0000_0000_0000_0000;
array[22811] <= 16'b0000_0000_0000_0000;
array[22812] <= 16'b0000_0000_0000_0000;
array[22813] <= 16'b0000_0000_0000_0000;
array[22814] <= 16'b0000_0000_0000_0000;
array[22815] <= 16'b0000_0000_0000_0000;
array[22816] <= 16'b0000_0000_0000_0000;
array[22817] <= 16'b0000_0000_0000_0000;
array[22818] <= 16'b0000_0000_0000_0000;
array[22819] <= 16'b0000_0000_0000_0000;
array[22820] <= 16'b0000_0000_0000_0000;
array[22821] <= 16'b0000_0000_0000_0000;
array[22822] <= 16'b0000_0000_0000_0000;
array[22823] <= 16'b0000_0000_0000_0000;
array[22824] <= 16'b0000_0000_0000_0000;
array[22825] <= 16'b0000_0000_0000_0000;
array[22826] <= 16'b0000_0000_0000_0000;
array[22827] <= 16'b0000_0000_0000_0000;
array[22828] <= 16'b0000_0000_0000_0000;
array[22829] <= 16'b0000_0000_0000_0000;
array[22830] <= 16'b0000_0000_0000_0000;
array[22831] <= 16'b0000_0000_0000_0000;
array[22832] <= 16'b0000_0000_0000_0000;
array[22833] <= 16'b0000_0000_0000_0000;
array[22834] <= 16'b0000_0000_0000_0000;
array[22835] <= 16'b0000_0000_0000_0000;
array[22836] <= 16'b0000_0000_0000_0000;
array[22837] <= 16'b0000_0000_0000_0000;
array[22838] <= 16'b0000_0000_0000_0000;
array[22839] <= 16'b0000_0000_0000_0000;
array[22840] <= 16'b0000_0000_0000_0000;
array[22841] <= 16'b0000_0000_0000_0000;
array[22842] <= 16'b0000_0000_0000_0000;
array[22843] <= 16'b0000_0000_0000_0000;
array[22844] <= 16'b0000_0000_0000_0000;
array[22845] <= 16'b0000_0000_0000_0000;
array[22846] <= 16'b0000_0000_0000_0000;
array[22847] <= 16'b0000_0000_0000_0000;
array[22848] <= 16'b0000_0000_0000_0000;
array[22849] <= 16'b0000_0000_0000_0000;
array[22850] <= 16'b0000_0000_0000_0000;
array[22851] <= 16'b0000_0000_0000_0000;
array[22852] <= 16'b0000_0000_0000_0000;
array[22853] <= 16'b0000_0000_0000_0000;
array[22854] <= 16'b0000_0000_0000_0000;
array[22855] <= 16'b0000_0000_0000_0000;
array[22856] <= 16'b0000_0000_0000_0000;
array[22857] <= 16'b0000_0000_0000_0000;
array[22858] <= 16'b0000_0000_0000_0000;
array[22859] <= 16'b0000_0000_0000_0000;
array[22860] <= 16'b0000_0000_0000_0000;
array[22861] <= 16'b0000_0000_0000_0000;
array[22862] <= 16'b0000_0000_0000_0000;
array[22863] <= 16'b0000_0000_0000_0000;
array[22864] <= 16'b0000_0000_0000_0000;
array[22865] <= 16'b0000_0000_0000_0000;
array[22866] <= 16'b0000_0000_0000_0000;
array[22867] <= 16'b0000_0000_0000_0000;
array[22868] <= 16'b0000_0000_0000_0000;
array[22869] <= 16'b0000_0000_0000_0000;
array[22870] <= 16'b0000_0000_0000_0000;
array[22871] <= 16'b0000_0000_0000_0000;
array[22872] <= 16'b0000_0000_0000_0000;
array[22873] <= 16'b0000_0000_0000_0000;
array[22874] <= 16'b0000_0000_0000_0000;
array[22875] <= 16'b0000_0000_0000_0000;
array[22876] <= 16'b0000_0000_0000_0000;
array[22877] <= 16'b0000_0000_0000_0000;
array[22878] <= 16'b0000_0000_0000_0000;
array[22879] <= 16'b0000_0000_0000_0000;
array[22880] <= 16'b0000_0000_0000_0000;
array[22881] <= 16'b0000_0000_0000_0000;
array[22882] <= 16'b0000_0000_0000_0000;
array[22883] <= 16'b0000_0000_0000_0000;
array[22884] <= 16'b0000_0000_0000_0000;
array[22885] <= 16'b0000_0000_0000_0000;
array[22886] <= 16'b0000_0000_0000_0000;
array[22887] <= 16'b0000_0000_0000_0000;
array[22888] <= 16'b0000_0000_0000_0000;
array[22889] <= 16'b0000_0000_0000_0000;
array[22890] <= 16'b0000_0000_0000_0000;
array[22891] <= 16'b0000_0000_0000_0000;
array[22892] <= 16'b0000_0000_0000_0000;
array[22893] <= 16'b0000_0000_0000_0000;
array[22894] <= 16'b0000_0000_0000_0000;
array[22895] <= 16'b0000_0000_0000_0000;
array[22896] <= 16'b0000_0000_0000_0000;
array[22897] <= 16'b0000_0000_0000_0000;
array[22898] <= 16'b0000_0000_0000_0000;
array[22899] <= 16'b0000_0000_0000_0000;
array[22900] <= 16'b0000_0000_0000_0000;
array[22901] <= 16'b0000_0000_0000_0000;
array[22902] <= 16'b0000_0000_0000_0000;
array[22903] <= 16'b0000_0000_0000_0000;
array[22904] <= 16'b0000_0000_0000_0000;
array[22905] <= 16'b0000_0000_0000_0000;
array[22906] <= 16'b0000_0000_0000_0000;
array[22907] <= 16'b0000_0000_0000_0000;
array[22908] <= 16'b0000_0000_0000_0000;
array[22909] <= 16'b0000_0000_0000_0000;
array[22910] <= 16'b0000_0000_0000_0000;
array[22911] <= 16'b0000_0000_0000_0000;
array[22912] <= 16'b0000_0000_0000_0000;
array[22913] <= 16'b0000_0000_0000_0000;
array[22914] <= 16'b0000_0000_0000_0000;
array[22915] <= 16'b0000_0000_0000_0000;
array[22916] <= 16'b0000_0000_0000_0000;
array[22917] <= 16'b0000_0000_0000_0000;
array[22918] <= 16'b0000_0000_0000_0000;
array[22919] <= 16'b0000_0000_0000_0000;
array[22920] <= 16'b0000_0000_0000_0000;
array[22921] <= 16'b0000_0000_0000_0000;
array[22922] <= 16'b0000_0000_0000_0000;
array[22923] <= 16'b0000_0000_0000_0000;
array[22924] <= 16'b0000_0000_0000_0000;
array[22925] <= 16'b0000_0000_0000_0000;
array[22926] <= 16'b0000_0000_0000_0000;
array[22927] <= 16'b0000_0000_0000_0000;
array[22928] <= 16'b0000_0000_0000_0000;
array[22929] <= 16'b0000_0000_0000_0000;
array[22930] <= 16'b0000_0000_0000_0000;
array[22931] <= 16'b0000_0000_0000_0000;
array[22932] <= 16'b0000_0000_0000_0000;
array[22933] <= 16'b0000_0000_0000_0000;
array[22934] <= 16'b0000_0000_0000_0000;
array[22935] <= 16'b0000_0000_0000_0000;
array[22936] <= 16'b0000_0000_0000_0000;
array[22937] <= 16'b0000_0000_0000_0000;
array[22938] <= 16'b0000_0000_0000_0000;
array[22939] <= 16'b0000_0000_0000_0000;
array[22940] <= 16'b0000_0000_0000_0000;
array[22941] <= 16'b0000_0000_0000_0000;
array[22942] <= 16'b0000_0000_0000_0000;
array[22943] <= 16'b0000_0000_0000_0000;
array[22944] <= 16'b0000_0000_0000_0000;
array[22945] <= 16'b0000_0000_0000_0000;
array[22946] <= 16'b0000_0000_0000_0000;
array[22947] <= 16'b0000_0000_0000_0000;
array[22948] <= 16'b0000_0000_0000_0000;
array[22949] <= 16'b0000_0000_0000_0000;
array[22950] <= 16'b0000_0000_0000_0000;
array[22951] <= 16'b0000_0000_0000_0000;
array[22952] <= 16'b0000_0000_0000_0000;
array[22953] <= 16'b0000_0000_0000_0000;
array[22954] <= 16'b0000_0000_0000_0000;
array[22955] <= 16'b0000_0000_0000_0000;
array[22956] <= 16'b0000_0000_0000_0000;
array[22957] <= 16'b0000_0000_0000_0000;
array[22958] <= 16'b0000_0000_0000_0000;
array[22959] <= 16'b0000_0000_0000_0000;
array[22960] <= 16'b0000_0000_0000_0000;
array[22961] <= 16'b0000_0000_0000_0000;
array[22962] <= 16'b0000_0000_0000_0000;
array[22963] <= 16'b0000_0000_0000_0000;
array[22964] <= 16'b0000_0000_0000_0000;
array[22965] <= 16'b0000_0000_0000_0000;
array[22966] <= 16'b0000_0000_0000_0000;
array[22967] <= 16'b0000_0000_0000_0000;
array[22968] <= 16'b0000_0000_0000_0000;
array[22969] <= 16'b0000_0000_0000_0000;
array[22970] <= 16'b0000_0000_0000_0000;
array[22971] <= 16'b0000_0000_0000_0000;
array[22972] <= 16'b0000_0000_0000_0000;
array[22973] <= 16'b0000_0000_0000_0000;
array[22974] <= 16'b0000_0000_0000_0000;
array[22975] <= 16'b0000_0000_0000_0000;
array[22976] <= 16'b0000_0000_0000_0000;
array[22977] <= 16'b0000_0000_0000_0000;
array[22978] <= 16'b0000_0000_0000_0000;
array[22979] <= 16'b0000_0000_0000_0000;
array[22980] <= 16'b0000_0000_0000_0000;
array[22981] <= 16'b0000_0000_0000_0000;
array[22982] <= 16'b0000_0000_0000_0000;
array[22983] <= 16'b0000_0000_0000_0000;
array[22984] <= 16'b0000_0000_0000_0000;
array[22985] <= 16'b0000_0000_0000_0000;
array[22986] <= 16'b0000_0000_0000_0000;
array[22987] <= 16'b0000_0000_0000_0000;
array[22988] <= 16'b0000_0000_0000_0000;
array[22989] <= 16'b0000_0000_0000_0000;
array[22990] <= 16'b0000_0000_0000_0000;
array[22991] <= 16'b0000_0000_0000_0000;
array[22992] <= 16'b0000_0000_0000_0000;
array[22993] <= 16'b0000_0000_0000_0000;
array[22994] <= 16'b0000_0000_0000_0000;
array[22995] <= 16'b0000_0000_0000_0000;
array[22996] <= 16'b0000_0000_0000_0000;
array[22997] <= 16'b0000_0000_0000_0000;
array[22998] <= 16'b0000_0000_0000_0000;
array[22999] <= 16'b0000_0000_0000_0000;
array[23000] <= 16'b0000_0000_0000_0000;
array[23001] <= 16'b0000_0000_0000_0000;
array[23002] <= 16'b0000_0000_0000_0000;
array[23003] <= 16'b0000_0000_0000_0000;
array[23004] <= 16'b0000_0000_0000_0000;
array[23005] <= 16'b0000_0000_0000_0000;
array[23006] <= 16'b0000_0000_0000_0000;
array[23007] <= 16'b0000_0000_0000_0000;
array[23008] <= 16'b0000_0000_0000_0000;
array[23009] <= 16'b0000_0000_0000_0000;
array[23010] <= 16'b0000_0000_0000_0000;
array[23011] <= 16'b0000_0000_0000_0000;
array[23012] <= 16'b0000_0000_0000_0000;
array[23013] <= 16'b0000_0000_0000_0000;
array[23014] <= 16'b0000_0000_0000_0000;
array[23015] <= 16'b0000_0000_0000_0000;
array[23016] <= 16'b0000_0000_0000_0000;
array[23017] <= 16'b0000_0000_0000_0000;
array[23018] <= 16'b0000_0000_0000_0000;
array[23019] <= 16'b0000_0000_0000_0000;
array[23020] <= 16'b0000_0000_0000_0000;
array[23021] <= 16'b0000_0000_0000_0000;
array[23022] <= 16'b0000_0000_0000_0000;
array[23023] <= 16'b0000_0000_0000_0000;
array[23024] <= 16'b0000_0000_0000_0000;
array[23025] <= 16'b0000_0000_0000_0000;
array[23026] <= 16'b0000_0000_0000_0000;
array[23027] <= 16'b0000_0000_0000_0000;
array[23028] <= 16'b0000_0000_0000_0000;
array[23029] <= 16'b0000_0000_0000_0000;
array[23030] <= 16'b0000_0000_0000_0000;
array[23031] <= 16'b0000_0000_0000_0000;
array[23032] <= 16'b0000_0000_0000_0000;
array[23033] <= 16'b0000_0000_0000_0000;
array[23034] <= 16'b0000_0000_0000_0000;
array[23035] <= 16'b0000_0000_0000_0000;
array[23036] <= 16'b0000_0000_0000_0000;
array[23037] <= 16'b0000_0000_0000_0000;
array[23038] <= 16'b0000_0000_0000_0000;
array[23039] <= 16'b0000_0000_0000_0000;
array[23040] <= 16'b0000_0000_0000_0000;
array[23041] <= 16'b0000_0000_0000_0000;
array[23042] <= 16'b0000_0000_0000_0000;
array[23043] <= 16'b0000_0000_0000_0000;
array[23044] <= 16'b0000_0000_0000_0000;
array[23045] <= 16'b0000_0000_0000_0000;
array[23046] <= 16'b0000_0000_0000_0000;
array[23047] <= 16'b0000_0000_0000_0000;
array[23048] <= 16'b0000_0000_0000_0000;
array[23049] <= 16'b0000_0000_0000_0000;
array[23050] <= 16'b0000_0000_0000_0000;
array[23051] <= 16'b0000_0000_0000_0000;
array[23052] <= 16'b0000_0000_0000_0000;
array[23053] <= 16'b0000_0000_0000_0000;
array[23054] <= 16'b0000_0000_0000_0000;
array[23055] <= 16'b0000_0000_0000_0000;
array[23056] <= 16'b0000_0000_0000_0000;
array[23057] <= 16'b0000_0000_0000_0000;
array[23058] <= 16'b0000_0000_0000_0000;
array[23059] <= 16'b0000_0000_0000_0000;
array[23060] <= 16'b0000_0000_0000_0000;
array[23061] <= 16'b0000_0000_0000_0000;
array[23062] <= 16'b0000_0000_0000_0000;
array[23063] <= 16'b0000_0000_0000_0000;
array[23064] <= 16'b0000_0000_0000_0000;
array[23065] <= 16'b0000_0000_0000_0000;
array[23066] <= 16'b0000_0000_0000_0000;
array[23067] <= 16'b0000_0000_0000_0000;
array[23068] <= 16'b0000_0000_0000_0000;
array[23069] <= 16'b0000_0000_0000_0000;
array[23070] <= 16'b0000_0000_0000_0000;
array[23071] <= 16'b0000_0000_0000_0000;
array[23072] <= 16'b0000_0000_0000_0000;
array[23073] <= 16'b0000_0000_0000_0000;
array[23074] <= 16'b0000_0000_0000_0000;
array[23075] <= 16'b0000_0000_0000_0000;
array[23076] <= 16'b0000_0000_0000_0000;
array[23077] <= 16'b0000_0000_0000_0000;
array[23078] <= 16'b0000_0000_0000_0000;
array[23079] <= 16'b0000_0000_0000_0000;
array[23080] <= 16'b0000_0000_0000_0000;
array[23081] <= 16'b0000_0000_0000_0000;
array[23082] <= 16'b0000_0000_0000_0000;
array[23083] <= 16'b0000_0000_0000_0000;
array[23084] <= 16'b0000_0000_0000_0000;
array[23085] <= 16'b0000_0000_0000_0000;
array[23086] <= 16'b0000_0000_0000_0000;
array[23087] <= 16'b0000_0000_0000_0000;
array[23088] <= 16'b0000_0000_0000_0000;
array[23089] <= 16'b0000_0000_0000_0000;
array[23090] <= 16'b0000_0000_0000_0000;
array[23091] <= 16'b0000_0000_0000_0000;
array[23092] <= 16'b0000_0000_0000_0000;
array[23093] <= 16'b0000_0000_0000_0000;
array[23094] <= 16'b0000_0000_0000_0000;
array[23095] <= 16'b0000_0000_0000_0000;
array[23096] <= 16'b0000_0000_0000_0000;
array[23097] <= 16'b0000_0000_0000_0000;
array[23098] <= 16'b0000_0000_0000_0000;
array[23099] <= 16'b0000_0000_0000_0000;
array[23100] <= 16'b0000_0000_0000_0000;
array[23101] <= 16'b0000_0000_0000_0000;
array[23102] <= 16'b0000_0000_0000_0000;
array[23103] <= 16'b0000_0000_0000_0000;
array[23104] <= 16'b0000_0000_0000_0000;
array[23105] <= 16'b0000_0000_0000_0000;
array[23106] <= 16'b0000_0000_0000_0000;
array[23107] <= 16'b0000_0000_0000_0000;
array[23108] <= 16'b0000_0000_0000_0000;
array[23109] <= 16'b0000_0000_0000_0000;
array[23110] <= 16'b0000_0000_0000_0000;
array[23111] <= 16'b0000_0000_0000_0000;
array[23112] <= 16'b0000_0000_0000_0000;
array[23113] <= 16'b0000_0000_0000_0000;
array[23114] <= 16'b0000_0000_0000_0000;
array[23115] <= 16'b0000_0000_0000_0000;
array[23116] <= 16'b0000_0000_0000_0000;
array[23117] <= 16'b0000_0000_0000_0000;
array[23118] <= 16'b0000_0000_0000_0000;
array[23119] <= 16'b0000_0000_0000_0000;
array[23120] <= 16'b0000_0000_0000_0000;
array[23121] <= 16'b0000_0000_0000_0000;
array[23122] <= 16'b0000_0000_0000_0000;
array[23123] <= 16'b0000_0000_0000_0000;
array[23124] <= 16'b0000_0000_0000_0000;
array[23125] <= 16'b0000_0000_0000_0000;
array[23126] <= 16'b0000_0000_0000_0000;
array[23127] <= 16'b0000_0000_0000_0000;
array[23128] <= 16'b0000_0000_0000_0000;
array[23129] <= 16'b0000_0000_0000_0000;
array[23130] <= 16'b0000_0000_0000_0000;
array[23131] <= 16'b0000_0000_0000_0000;
array[23132] <= 16'b0000_0000_0000_0000;
array[23133] <= 16'b0000_0000_0000_0000;
array[23134] <= 16'b0000_0000_0000_0000;
array[23135] <= 16'b0000_0000_0000_0000;
array[23136] <= 16'b0000_0000_0000_0000;
array[23137] <= 16'b0000_0000_0000_0000;
array[23138] <= 16'b0000_0000_0000_0000;
array[23139] <= 16'b0000_0000_0000_0000;
array[23140] <= 16'b0000_0000_0000_0000;
array[23141] <= 16'b0000_0000_0000_0000;
array[23142] <= 16'b0000_0000_0000_0000;
array[23143] <= 16'b0000_0000_0000_0000;
array[23144] <= 16'b0000_0000_0000_0000;
array[23145] <= 16'b0000_0000_0000_0000;
array[23146] <= 16'b0000_0000_0000_0000;
array[23147] <= 16'b0000_0000_0000_0000;
array[23148] <= 16'b0000_0000_0000_0000;
array[23149] <= 16'b0000_0000_0000_0000;
array[23150] <= 16'b0000_0000_0000_0000;
array[23151] <= 16'b0000_0000_0000_0000;
array[23152] <= 16'b0000_0000_0000_0000;
array[23153] <= 16'b0000_0000_0000_0000;
array[23154] <= 16'b0000_0000_0000_0000;
array[23155] <= 16'b0000_0000_0000_0000;
array[23156] <= 16'b0000_0000_0000_0000;
array[23157] <= 16'b0000_0000_0000_0000;
array[23158] <= 16'b0000_0000_0000_0000;
array[23159] <= 16'b0000_0000_0000_0000;
array[23160] <= 16'b0000_0000_0000_0000;
array[23161] <= 16'b0000_0000_0000_0000;
array[23162] <= 16'b0000_0000_0000_0000;
array[23163] <= 16'b0000_0000_0000_0000;
array[23164] <= 16'b0000_0000_0000_0000;
array[23165] <= 16'b0000_0000_0000_0000;
array[23166] <= 16'b0000_0000_0000_0000;
array[23167] <= 16'b0000_0000_0000_0000;
array[23168] <= 16'b0000_0000_0000_0000;
array[23169] <= 16'b0000_0000_0000_0000;
array[23170] <= 16'b0000_0000_0000_0000;
array[23171] <= 16'b0000_0000_0000_0000;
array[23172] <= 16'b0000_0000_0000_0000;
array[23173] <= 16'b0000_0000_0000_0000;
array[23174] <= 16'b0000_0000_0000_0000;
array[23175] <= 16'b0000_0000_0000_0000;
array[23176] <= 16'b0000_0000_0000_0000;
array[23177] <= 16'b0000_0000_0000_0000;
array[23178] <= 16'b0000_0000_0000_0000;
array[23179] <= 16'b0000_0000_0000_0000;
array[23180] <= 16'b0000_0000_0000_0000;
array[23181] <= 16'b0000_0000_0000_0000;
array[23182] <= 16'b0000_0000_0000_0000;
array[23183] <= 16'b0000_0000_0000_0000;
array[23184] <= 16'b0000_0000_0000_0000;
array[23185] <= 16'b0000_0000_0000_0000;
array[23186] <= 16'b0000_0000_0000_0000;
array[23187] <= 16'b0000_0000_0000_0000;
array[23188] <= 16'b0000_0000_0000_0000;
array[23189] <= 16'b0000_0000_0000_0000;
array[23190] <= 16'b0000_0000_0000_0000;
array[23191] <= 16'b0000_0000_0000_0000;
array[23192] <= 16'b0000_0000_0000_0000;
array[23193] <= 16'b0000_0000_0000_0000;
array[23194] <= 16'b0000_0000_0000_0000;
array[23195] <= 16'b0000_0000_0000_0000;
array[23196] <= 16'b0000_0000_0000_0000;
array[23197] <= 16'b0000_0000_0000_0000;
array[23198] <= 16'b0000_0000_0000_0000;
array[23199] <= 16'b0000_0000_0000_0000;
array[23200] <= 16'b0000_0000_0000_0000;
array[23201] <= 16'b0000_0000_0000_0000;
array[23202] <= 16'b0000_0000_0000_0000;
array[23203] <= 16'b0000_0000_0000_0000;
array[23204] <= 16'b0000_0000_0000_0000;
array[23205] <= 16'b0000_0000_0000_0000;
array[23206] <= 16'b0000_0000_0000_0000;
array[23207] <= 16'b0000_0000_0000_0000;
array[23208] <= 16'b0000_0000_0000_0000;
array[23209] <= 16'b0000_0000_0000_0000;
array[23210] <= 16'b0000_0000_0000_0000;
array[23211] <= 16'b0000_0000_0000_0000;
array[23212] <= 16'b0000_0000_0000_0000;
array[23213] <= 16'b0000_0000_0000_0000;
array[23214] <= 16'b0000_0000_0000_0000;
array[23215] <= 16'b0000_0000_0000_0000;
array[23216] <= 16'b0000_0000_0000_0000;
array[23217] <= 16'b0000_0000_0000_0000;
array[23218] <= 16'b0000_0000_0000_0000;
array[23219] <= 16'b0000_0000_0000_0000;
array[23220] <= 16'b0000_0000_0000_0000;
array[23221] <= 16'b0000_0000_0000_0000;
array[23222] <= 16'b0000_0000_0000_0000;
array[23223] <= 16'b0000_0000_0000_0000;
array[23224] <= 16'b0000_0000_0000_0000;
array[23225] <= 16'b0000_0000_0000_0000;
array[23226] <= 16'b0000_0000_0000_0000;
array[23227] <= 16'b0000_0000_0000_0000;
array[23228] <= 16'b0000_0000_0000_0000;
array[23229] <= 16'b0000_0000_0000_0000;
array[23230] <= 16'b0000_0000_0000_0000;
array[23231] <= 16'b0000_0000_0000_0000;
array[23232] <= 16'b0000_0000_0000_0000;
array[23233] <= 16'b0000_0000_0000_0000;
array[23234] <= 16'b0000_0000_0000_0000;
array[23235] <= 16'b0000_0000_0000_0000;
array[23236] <= 16'b0000_0000_0000_0000;
array[23237] <= 16'b0000_0000_0000_0000;
array[23238] <= 16'b0000_0000_0000_0000;
array[23239] <= 16'b0000_0000_0000_0000;
array[23240] <= 16'b0000_0000_0000_0000;
array[23241] <= 16'b0000_0000_0000_0000;
array[23242] <= 16'b0000_0000_0000_0000;
array[23243] <= 16'b0000_0000_0000_0000;
array[23244] <= 16'b0000_0000_0000_0000;
array[23245] <= 16'b0000_0000_0000_0000;
array[23246] <= 16'b0000_0000_0000_0000;
array[23247] <= 16'b0000_0000_0000_0000;
array[23248] <= 16'b0000_0000_0000_0000;
array[23249] <= 16'b0000_0000_0000_0000;
array[23250] <= 16'b0000_0000_0000_0000;
array[23251] <= 16'b0000_0000_0000_0000;
array[23252] <= 16'b0000_0000_0000_0000;
array[23253] <= 16'b0000_0000_0000_0000;
array[23254] <= 16'b0000_0000_0000_0000;
array[23255] <= 16'b0000_0000_0000_0000;
array[23256] <= 16'b0000_0000_0000_0000;
array[23257] <= 16'b0000_0000_0000_0000;
array[23258] <= 16'b0000_0000_0000_0000;
array[23259] <= 16'b0000_0000_0000_0000;
array[23260] <= 16'b0000_0000_0000_0000;
array[23261] <= 16'b0000_0000_0000_0000;
array[23262] <= 16'b0000_0000_0000_0000;
array[23263] <= 16'b0000_0000_0000_0000;
array[23264] <= 16'b0000_0000_0000_0000;
array[23265] <= 16'b0000_0000_0000_0000;
array[23266] <= 16'b0000_0000_0000_0000;
array[23267] <= 16'b0000_0000_0000_0000;
array[23268] <= 16'b0000_0000_0000_0000;
array[23269] <= 16'b0000_0000_0000_0000;
array[23270] <= 16'b0000_0000_0000_0000;
array[23271] <= 16'b0000_0000_0000_0000;
array[23272] <= 16'b0000_0000_0000_0000;
array[23273] <= 16'b0000_0000_0000_0000;
array[23274] <= 16'b0000_0000_0000_0000;
array[23275] <= 16'b0000_0000_0000_0000;
array[23276] <= 16'b0000_0000_0000_0000;
array[23277] <= 16'b0000_0000_0000_0000;
array[23278] <= 16'b0000_0000_0000_0000;
array[23279] <= 16'b0000_0000_0000_0000;
array[23280] <= 16'b0000_0000_0000_0000;
array[23281] <= 16'b0000_0000_0000_0000;
array[23282] <= 16'b0000_0000_0000_0000;
array[23283] <= 16'b0000_0000_0000_0000;
array[23284] <= 16'b0000_0000_0000_0000;
array[23285] <= 16'b0000_0000_0000_0000;
array[23286] <= 16'b0000_0000_0000_0000;
array[23287] <= 16'b0000_0000_0000_0000;
array[23288] <= 16'b0000_0000_0000_0000;
array[23289] <= 16'b0000_0000_0000_0000;
array[23290] <= 16'b0000_0000_0000_0000;
array[23291] <= 16'b0000_0000_0000_0000;
array[23292] <= 16'b0000_0000_0000_0000;
array[23293] <= 16'b0000_0000_0000_0000;
array[23294] <= 16'b0000_0000_0000_0000;
array[23295] <= 16'b0000_0000_0000_0000;
array[23296] <= 16'b0000_0000_0000_0000;
array[23297] <= 16'b0000_0000_0000_0000;
array[23298] <= 16'b0000_0000_0000_0000;
array[23299] <= 16'b0000_0000_0000_0000;
array[23300] <= 16'b0000_0000_0000_0000;
array[23301] <= 16'b0000_0000_0000_0000;
array[23302] <= 16'b0000_0000_0000_0000;
array[23303] <= 16'b0000_0000_0000_0000;
array[23304] <= 16'b0000_0000_0000_0000;
array[23305] <= 16'b0000_0000_0000_0000;
array[23306] <= 16'b0000_0000_0000_0000;
array[23307] <= 16'b0000_0000_0000_0000;
array[23308] <= 16'b0000_0000_0000_0000;
array[23309] <= 16'b0000_0000_0000_0000;
array[23310] <= 16'b0000_0000_0000_0000;
array[23311] <= 16'b0000_0000_0000_0000;
array[23312] <= 16'b0000_0000_0000_0000;
array[23313] <= 16'b0000_0000_0000_0000;
array[23314] <= 16'b0000_0000_0000_0000;
array[23315] <= 16'b0000_0000_0000_0000;
array[23316] <= 16'b0000_0000_0000_0000;
array[23317] <= 16'b0000_0000_0000_0000;
array[23318] <= 16'b0000_0000_0000_0000;
array[23319] <= 16'b0000_0000_0000_0000;
array[23320] <= 16'b0000_0000_0000_0000;
array[23321] <= 16'b0000_0000_0000_0000;
array[23322] <= 16'b0000_0000_0000_0000;
array[23323] <= 16'b0000_0000_0000_0000;
array[23324] <= 16'b0000_0000_0000_0000;
array[23325] <= 16'b0000_0000_0000_0000;
array[23326] <= 16'b0000_0000_0000_0000;
array[23327] <= 16'b0000_0000_0000_0000;
array[23328] <= 16'b0000_0000_0000_0000;
array[23329] <= 16'b0000_0000_0000_0000;
array[23330] <= 16'b0000_0000_0000_0000;
array[23331] <= 16'b0000_0000_0000_0000;
array[23332] <= 16'b0000_0000_0000_0000;
array[23333] <= 16'b0000_0000_0000_0000;
array[23334] <= 16'b0000_0000_0000_0000;
array[23335] <= 16'b0000_0000_0000_0000;
array[23336] <= 16'b0000_0000_0000_0000;
array[23337] <= 16'b0000_0000_0000_0000;
array[23338] <= 16'b0000_0000_0000_0000;
array[23339] <= 16'b0000_0000_0000_0000;
array[23340] <= 16'b0000_0000_0000_0000;
array[23341] <= 16'b0000_0000_0000_0000;
array[23342] <= 16'b0000_0000_0000_0000;
array[23343] <= 16'b0000_0000_0000_0000;
array[23344] <= 16'b0000_0000_0000_0000;
array[23345] <= 16'b0000_0000_0000_0000;
array[23346] <= 16'b0000_0000_0000_0000;
array[23347] <= 16'b0000_0000_0000_0000;
array[23348] <= 16'b0000_0000_0000_0000;
array[23349] <= 16'b0000_0000_0000_0000;
array[23350] <= 16'b0000_0000_0000_0000;
array[23351] <= 16'b0000_0000_0000_0000;
array[23352] <= 16'b0000_0000_0000_0000;
array[23353] <= 16'b0000_0000_0000_0000;
array[23354] <= 16'b0000_0000_0000_0000;
array[23355] <= 16'b0000_0000_0000_0000;
array[23356] <= 16'b0000_0000_0000_0000;
array[23357] <= 16'b0000_0000_0000_0000;
array[23358] <= 16'b0000_0000_0000_0000;
array[23359] <= 16'b0000_0000_0000_0000;
array[23360] <= 16'b0000_0000_0000_0000;
array[23361] <= 16'b0000_0000_0000_0000;
array[23362] <= 16'b0000_0000_0000_0000;
array[23363] <= 16'b0000_0000_0000_0000;
array[23364] <= 16'b0000_0000_0000_0000;
array[23365] <= 16'b0000_0000_0000_0000;
array[23366] <= 16'b0000_0000_0000_0000;
array[23367] <= 16'b0000_0000_0000_0000;
array[23368] <= 16'b0000_0000_0000_0000;
array[23369] <= 16'b0000_0000_0000_0000;
array[23370] <= 16'b0000_0000_0000_0000;
array[23371] <= 16'b0000_0000_0000_0000;
array[23372] <= 16'b0000_0000_0000_0000;
array[23373] <= 16'b0000_0000_0000_0000;
array[23374] <= 16'b0000_0000_0000_0000;
array[23375] <= 16'b0000_0000_0000_0000;
array[23376] <= 16'b0000_0000_0000_0000;
array[23377] <= 16'b0000_0000_0000_0000;
array[23378] <= 16'b0000_0000_0000_0000;
array[23379] <= 16'b0000_0000_0000_0000;
array[23380] <= 16'b0000_0000_0000_0000;
array[23381] <= 16'b0000_0000_0000_0000;
array[23382] <= 16'b0000_0000_0000_0000;
array[23383] <= 16'b0000_0000_0000_0000;
array[23384] <= 16'b0000_0000_0000_0000;
array[23385] <= 16'b0000_0000_0000_0000;
array[23386] <= 16'b0000_0000_0000_0000;
array[23387] <= 16'b0000_0000_0000_0000;
array[23388] <= 16'b0000_0000_0000_0000;
array[23389] <= 16'b0000_0000_0000_0000;
array[23390] <= 16'b0000_0000_0000_0000;
array[23391] <= 16'b0000_0000_0000_0000;
array[23392] <= 16'b0000_0000_0000_0000;
array[23393] <= 16'b0000_0000_0000_0000;
array[23394] <= 16'b0000_0000_0000_0000;
array[23395] <= 16'b0000_0000_0000_0000;
array[23396] <= 16'b0000_0000_0000_0000;
array[23397] <= 16'b0000_0000_0000_0000;
array[23398] <= 16'b0000_0000_0000_0000;
array[23399] <= 16'b0000_0000_0000_0000;
array[23400] <= 16'b0000_0000_0000_0000;
array[23401] <= 16'b0000_0000_0000_0000;
array[23402] <= 16'b0000_0000_0000_0000;
array[23403] <= 16'b0000_0000_0000_0000;
array[23404] <= 16'b0000_0000_0000_0000;
array[23405] <= 16'b0000_0000_0000_0000;
array[23406] <= 16'b0000_0000_0000_0000;
array[23407] <= 16'b0000_0000_0000_0000;
array[23408] <= 16'b0000_0000_0000_0000;
array[23409] <= 16'b0000_0000_0000_0000;
array[23410] <= 16'b0000_0000_0000_0000;
array[23411] <= 16'b0000_0000_0000_0000;
array[23412] <= 16'b0000_0000_0000_0000;
array[23413] <= 16'b0000_0000_0000_0000;
array[23414] <= 16'b0000_0000_0000_0000;
array[23415] <= 16'b0000_0000_0000_0000;
array[23416] <= 16'b0000_0000_0000_0000;
array[23417] <= 16'b0000_0000_0000_0000;
array[23418] <= 16'b0000_0000_0000_0000;
array[23419] <= 16'b0000_0000_0000_0000;
array[23420] <= 16'b0000_0000_0000_0000;
array[23421] <= 16'b0000_0000_0000_0000;
array[23422] <= 16'b0000_0000_0000_0000;
array[23423] <= 16'b0000_0000_0000_0000;
array[23424] <= 16'b0000_0000_0000_0000;
array[23425] <= 16'b0000_0000_0000_0000;
array[23426] <= 16'b0000_0000_0000_0000;
array[23427] <= 16'b0000_0000_0000_0000;
array[23428] <= 16'b0000_0000_0000_0000;
array[23429] <= 16'b0000_0000_0000_0000;
array[23430] <= 16'b0000_0000_0000_0000;
array[23431] <= 16'b0000_0000_0000_0000;
array[23432] <= 16'b0000_0000_0000_0000;
array[23433] <= 16'b0000_0000_0000_0000;
array[23434] <= 16'b0000_0000_0000_0000;
array[23435] <= 16'b0000_0000_0000_0000;
array[23436] <= 16'b0000_0000_0000_0000;
array[23437] <= 16'b0000_0000_0000_0000;
array[23438] <= 16'b0000_0000_0000_0000;
array[23439] <= 16'b0000_0000_0000_0000;
array[23440] <= 16'b0000_0000_0000_0000;
array[23441] <= 16'b0000_0000_0000_0000;
array[23442] <= 16'b0000_0000_0000_0000;
array[23443] <= 16'b0000_0000_0000_0000;
array[23444] <= 16'b0000_0000_0000_0000;
array[23445] <= 16'b0000_0000_0000_0000;
array[23446] <= 16'b0000_0000_0000_0000;
array[23447] <= 16'b0000_0000_0000_0000;
array[23448] <= 16'b0000_0000_0000_0000;
array[23449] <= 16'b0000_0000_0000_0000;
array[23450] <= 16'b0000_0000_0000_0000;
array[23451] <= 16'b0000_0000_0000_0000;
array[23452] <= 16'b0000_0000_0000_0000;
array[23453] <= 16'b0000_0000_0000_0000;
array[23454] <= 16'b0000_0000_0000_0000;
array[23455] <= 16'b0000_0000_0000_0000;
array[23456] <= 16'b0000_0000_0000_0000;
array[23457] <= 16'b0000_0000_0000_0000;
array[23458] <= 16'b0000_0000_0000_0000;
array[23459] <= 16'b0000_0000_0000_0000;
array[23460] <= 16'b0000_0000_0000_0000;
array[23461] <= 16'b0000_0000_0000_0000;
array[23462] <= 16'b0000_0000_0000_0000;
array[23463] <= 16'b0000_0000_0000_0000;
array[23464] <= 16'b0000_0000_0000_0000;
array[23465] <= 16'b0000_0000_0000_0000;
array[23466] <= 16'b0000_0000_0000_0000;
array[23467] <= 16'b0000_0000_0000_0000;
array[23468] <= 16'b0000_0000_0000_0000;
array[23469] <= 16'b0000_0000_0000_0000;
array[23470] <= 16'b0000_0000_0000_0000;
array[23471] <= 16'b0000_0000_0000_0000;
array[23472] <= 16'b0000_0000_0000_0000;
array[23473] <= 16'b0000_0000_0000_0000;
array[23474] <= 16'b0000_0000_0000_0000;
array[23475] <= 16'b0000_0000_0000_0000;
array[23476] <= 16'b0000_0000_0000_0000;
array[23477] <= 16'b0000_0000_0000_0000;
array[23478] <= 16'b0000_0000_0000_0000;
array[23479] <= 16'b0000_0000_0000_0000;
array[23480] <= 16'b0000_0000_0000_0000;
array[23481] <= 16'b0000_0000_0000_0000;
array[23482] <= 16'b0000_0000_0000_0000;
array[23483] <= 16'b0000_0000_0000_0000;
array[23484] <= 16'b0000_0000_0000_0000;
array[23485] <= 16'b0000_0000_0000_0000;
array[23486] <= 16'b0000_0000_0000_0000;
array[23487] <= 16'b0000_0000_0000_0000;
array[23488] <= 16'b0000_0000_0000_0000;
array[23489] <= 16'b0000_0000_0000_0000;
array[23490] <= 16'b0000_0000_0000_0000;
array[23491] <= 16'b0000_0000_0000_0000;
array[23492] <= 16'b0000_0000_0000_0000;
array[23493] <= 16'b0000_0000_0000_0000;
array[23494] <= 16'b0000_0000_0000_0000;
array[23495] <= 16'b0000_0000_0000_0000;
array[23496] <= 16'b0000_0000_0000_0000;
array[23497] <= 16'b0000_0000_0000_0000;
array[23498] <= 16'b0000_0000_0000_0000;
array[23499] <= 16'b0000_0000_0000_0000;
array[23500] <= 16'b0000_0000_0000_0000;
array[23501] <= 16'b0000_0000_0000_0000;
array[23502] <= 16'b0000_0000_0000_0000;
array[23503] <= 16'b0000_0000_0000_0000;
array[23504] <= 16'b0000_0000_0000_0000;
array[23505] <= 16'b0000_0000_0000_0000;
array[23506] <= 16'b0000_0000_0000_0000;
array[23507] <= 16'b0000_0000_0000_0000;
array[23508] <= 16'b0000_0000_0000_0000;
array[23509] <= 16'b0000_0000_0000_0000;
array[23510] <= 16'b0000_0000_0000_0000;
array[23511] <= 16'b0000_0000_0000_0000;
array[23512] <= 16'b0000_0000_0000_0000;
array[23513] <= 16'b0000_0000_0000_0000;
array[23514] <= 16'b0000_0000_0000_0000;
array[23515] <= 16'b0000_0000_0000_0000;
array[23516] <= 16'b0000_0000_0000_0000;
array[23517] <= 16'b0000_0000_0000_0000;
array[23518] <= 16'b0000_0000_0000_0000;
array[23519] <= 16'b0000_0000_0000_0000;
array[23520] <= 16'b0000_0000_0000_0000;
array[23521] <= 16'b0000_0000_0000_0000;
array[23522] <= 16'b0000_0000_0000_0000;
array[23523] <= 16'b0000_0000_0000_0000;
array[23524] <= 16'b0000_0000_0000_0000;
array[23525] <= 16'b0000_0000_0000_0000;
array[23526] <= 16'b0000_0000_0000_0000;
array[23527] <= 16'b0000_0000_0000_0000;
array[23528] <= 16'b0000_0000_0000_0000;
array[23529] <= 16'b0000_0000_0000_0000;
array[23530] <= 16'b0000_0000_0000_0000;
array[23531] <= 16'b0000_0000_0000_0000;
array[23532] <= 16'b0000_0000_0000_0000;
array[23533] <= 16'b0000_0000_0000_0000;
array[23534] <= 16'b0000_0000_0000_0000;
array[23535] <= 16'b0000_0000_0000_0000;
array[23536] <= 16'b0000_0000_0000_0000;
array[23537] <= 16'b0000_0000_0000_0000;
array[23538] <= 16'b0000_0000_0000_0000;
array[23539] <= 16'b0000_0000_0000_0000;
array[23540] <= 16'b0000_0000_0000_0000;
array[23541] <= 16'b0000_0000_0000_0000;
array[23542] <= 16'b0000_0000_0000_0000;
array[23543] <= 16'b0000_0000_0000_0000;
array[23544] <= 16'b0000_0000_0000_0000;
array[23545] <= 16'b0000_0000_0000_0000;
array[23546] <= 16'b0000_0000_0000_0000;
array[23547] <= 16'b0000_0000_0000_0000;
array[23548] <= 16'b0000_0000_0000_0000;
array[23549] <= 16'b0000_0000_0000_0000;
array[23550] <= 16'b0000_0000_0000_0000;
array[23551] <= 16'b0000_0000_0000_0000;
array[23552] <= 16'b0000_0000_0000_0000;
array[23553] <= 16'b0000_0000_0000_0000;
array[23554] <= 16'b0000_0000_0000_0000;
array[23555] <= 16'b0000_0000_0000_0000;
array[23556] <= 16'b0000_0000_0000_0000;
array[23557] <= 16'b0000_0000_0000_0000;
array[23558] <= 16'b0000_0000_0000_0000;
array[23559] <= 16'b0000_0000_0000_0000;
array[23560] <= 16'b0000_0000_0000_0000;
array[23561] <= 16'b0000_0000_0000_0000;
array[23562] <= 16'b0000_0000_0000_0000;
array[23563] <= 16'b0000_0000_0000_0000;
array[23564] <= 16'b0000_0000_0000_0000;
array[23565] <= 16'b0000_0000_0000_0000;
array[23566] <= 16'b0000_0000_0000_0000;
array[23567] <= 16'b0000_0000_0000_0000;
array[23568] <= 16'b0000_0000_0000_0000;
array[23569] <= 16'b0000_0000_0000_0000;
array[23570] <= 16'b0000_0000_0000_0000;
array[23571] <= 16'b0000_0000_0000_0000;
array[23572] <= 16'b0000_0000_0000_0000;
array[23573] <= 16'b0000_0000_0000_0000;
array[23574] <= 16'b0000_0000_0000_0000;
array[23575] <= 16'b0000_0000_0000_0000;
array[23576] <= 16'b0000_0000_0000_0000;
array[23577] <= 16'b0000_0000_0000_0000;
array[23578] <= 16'b0000_0000_0000_0000;
array[23579] <= 16'b0000_0000_0000_0000;
array[23580] <= 16'b0000_0000_0000_0000;
array[23581] <= 16'b0000_0000_0000_0000;
array[23582] <= 16'b0000_0000_0000_0000;
array[23583] <= 16'b0000_0000_0000_0000;
array[23584] <= 16'b0000_0000_0000_0000;
array[23585] <= 16'b0000_0000_0000_0000;
array[23586] <= 16'b0000_0000_0000_0000;
array[23587] <= 16'b0000_0000_0000_0000;
array[23588] <= 16'b0000_0000_0000_0000;
array[23589] <= 16'b0000_0000_0000_0000;
array[23590] <= 16'b0000_0000_0000_0000;
array[23591] <= 16'b0000_0000_0000_0000;
array[23592] <= 16'b0000_0000_0000_0000;
array[23593] <= 16'b0000_0000_0000_0000;
array[23594] <= 16'b0000_0000_0000_0000;
array[23595] <= 16'b0000_0000_0000_0000;
array[23596] <= 16'b0000_0000_0000_0000;
array[23597] <= 16'b0000_0000_0000_0000;
array[23598] <= 16'b0000_0000_0000_0000;
array[23599] <= 16'b0000_0000_0000_0000;
array[23600] <= 16'b0000_0000_0000_0000;
array[23601] <= 16'b0000_0000_0000_0000;
array[23602] <= 16'b0000_0000_0000_0000;
array[23603] <= 16'b0000_0000_0000_0000;
array[23604] <= 16'b0000_0000_0000_0000;
array[23605] <= 16'b0000_0000_0000_0000;
array[23606] <= 16'b0000_0000_0000_0000;
array[23607] <= 16'b0000_0000_0000_0000;
array[23608] <= 16'b0000_0000_0000_0000;
array[23609] <= 16'b0000_0000_0000_0000;
array[23610] <= 16'b0000_0000_0000_0000;
array[23611] <= 16'b0000_0000_0000_0000;
array[23612] <= 16'b0000_0000_0000_0000;
array[23613] <= 16'b0000_0000_0000_0000;
array[23614] <= 16'b0000_0000_0000_0000;
array[23615] <= 16'b0000_0000_0000_0000;
array[23616] <= 16'b0000_0000_0000_0000;
array[23617] <= 16'b0000_0000_0000_0000;
array[23618] <= 16'b0000_0000_0000_0000;
array[23619] <= 16'b0000_0000_0000_0000;
array[23620] <= 16'b0000_0000_0000_0000;
array[23621] <= 16'b0000_0000_0000_0000;
array[23622] <= 16'b0000_0000_0000_0000;
array[23623] <= 16'b0000_0000_0000_0000;
array[23624] <= 16'b0000_0000_0000_0000;
array[23625] <= 16'b0000_0000_0000_0000;
array[23626] <= 16'b0000_0000_0000_0000;
array[23627] <= 16'b0000_0000_0000_0000;
array[23628] <= 16'b0000_0000_0000_0000;
array[23629] <= 16'b0000_0000_0000_0000;
array[23630] <= 16'b0000_0000_0000_0000;
array[23631] <= 16'b0000_0000_0000_0000;
array[23632] <= 16'b0000_0000_0000_0000;
array[23633] <= 16'b0000_0000_0000_0000;
array[23634] <= 16'b0000_0000_0000_0000;
array[23635] <= 16'b0000_0000_0000_0000;
array[23636] <= 16'b0000_0000_0000_0000;
array[23637] <= 16'b0000_0000_0000_0000;
array[23638] <= 16'b0000_0000_0000_0000;
array[23639] <= 16'b0000_0000_0000_0000;
array[23640] <= 16'b0000_0000_0000_0000;
array[23641] <= 16'b0000_0000_0000_0000;
array[23642] <= 16'b0000_0000_0000_0000;
array[23643] <= 16'b0000_0000_0000_0000;
array[23644] <= 16'b0000_0000_0000_0000;
array[23645] <= 16'b0000_0000_0000_0000;
array[23646] <= 16'b0000_0000_0000_0000;
array[23647] <= 16'b0000_0000_0000_0000;
array[23648] <= 16'b0000_0000_0000_0000;
array[23649] <= 16'b0000_0000_0000_0000;
array[23650] <= 16'b0000_0000_0000_0000;
array[23651] <= 16'b0000_0000_0000_0000;
array[23652] <= 16'b0000_0000_0000_0000;
array[23653] <= 16'b0000_0000_0000_0000;
array[23654] <= 16'b0000_0000_0000_0000;
array[23655] <= 16'b0000_0000_0000_0000;
array[23656] <= 16'b0000_0000_0000_0000;
array[23657] <= 16'b0000_0000_0000_0000;
array[23658] <= 16'b0000_0000_0000_0000;
array[23659] <= 16'b0000_0000_0000_0000;
array[23660] <= 16'b0000_0000_0000_0000;
array[23661] <= 16'b0000_0000_0000_0000;
array[23662] <= 16'b0000_0000_0000_0000;
array[23663] <= 16'b0000_0000_0000_0000;
array[23664] <= 16'b0000_0000_0000_0000;
array[23665] <= 16'b0000_0000_0000_0000;
array[23666] <= 16'b0000_0000_0000_0000;
array[23667] <= 16'b0000_0000_0000_0000;
array[23668] <= 16'b0000_0000_0000_0000;
array[23669] <= 16'b0000_0000_0000_0000;
array[23670] <= 16'b0000_0000_0000_0000;
array[23671] <= 16'b0000_0000_0000_0000;
array[23672] <= 16'b0000_0000_0000_0000;
array[23673] <= 16'b0000_0000_0000_0000;
array[23674] <= 16'b0000_0000_0000_0000;
array[23675] <= 16'b0000_0000_0000_0000;
array[23676] <= 16'b0000_0000_0000_0000;
array[23677] <= 16'b0000_0000_0000_0000;
array[23678] <= 16'b0000_0000_0000_0000;
array[23679] <= 16'b0000_0000_0000_0000;
array[23680] <= 16'b0000_0000_0000_0000;
array[23681] <= 16'b0000_0000_0000_0000;
array[23682] <= 16'b0000_0000_0000_0000;
array[23683] <= 16'b0000_0000_0000_0000;
array[23684] <= 16'b0000_0000_0000_0000;
array[23685] <= 16'b0000_0000_0000_0000;
array[23686] <= 16'b0000_0000_0000_0000;
array[23687] <= 16'b0000_0000_0000_0000;
array[23688] <= 16'b0000_0000_0000_0000;
array[23689] <= 16'b0000_0000_0000_0000;
array[23690] <= 16'b0000_0000_0000_0000;
array[23691] <= 16'b0000_0000_0000_0000;
array[23692] <= 16'b0000_0000_0000_0000;
array[23693] <= 16'b0000_0000_0000_0000;
array[23694] <= 16'b0000_0000_0000_0000;
array[23695] <= 16'b0000_0000_0000_0000;
array[23696] <= 16'b0000_0000_0000_0000;
array[23697] <= 16'b0000_0000_0000_0000;
array[23698] <= 16'b0000_0000_0000_0000;
array[23699] <= 16'b0000_0000_0000_0000;
array[23700] <= 16'b0000_0000_0000_0000;
array[23701] <= 16'b0000_0000_0000_0000;
array[23702] <= 16'b0000_0000_0000_0000;
array[23703] <= 16'b0000_0000_0000_0000;
array[23704] <= 16'b0000_0000_0000_0000;
array[23705] <= 16'b0000_0000_0000_0000;
array[23706] <= 16'b0000_0000_0000_0000;
array[23707] <= 16'b0000_0000_0000_0000;
array[23708] <= 16'b0000_0000_0000_0000;
array[23709] <= 16'b0000_0000_0000_0000;
array[23710] <= 16'b0000_0000_0000_0000;
array[23711] <= 16'b0000_0000_0000_0000;
array[23712] <= 16'b0000_0000_0000_0000;
array[23713] <= 16'b0000_0000_0000_0000;
array[23714] <= 16'b0000_0000_0000_0000;
array[23715] <= 16'b0000_0000_0000_0000;
array[23716] <= 16'b0000_0000_0000_0000;
array[23717] <= 16'b0000_0000_0000_0000;
array[23718] <= 16'b0000_0000_0000_0000;
array[23719] <= 16'b0000_0000_0000_0000;
array[23720] <= 16'b0000_0000_0000_0000;
array[23721] <= 16'b0000_0000_0000_0000;
array[23722] <= 16'b0000_0000_0000_0000;
array[23723] <= 16'b0000_0000_0000_0000;
array[23724] <= 16'b0000_0000_0000_0000;
array[23725] <= 16'b0000_0000_0000_0000;
array[23726] <= 16'b0000_0000_0000_0000;
array[23727] <= 16'b0000_0000_0000_0000;
array[23728] <= 16'b0000_0000_0000_0000;
array[23729] <= 16'b0000_0000_0000_0000;
array[23730] <= 16'b0000_0000_0000_0000;
array[23731] <= 16'b0000_0000_0000_0000;
array[23732] <= 16'b0000_0000_0000_0000;
array[23733] <= 16'b0000_0000_0000_0000;
array[23734] <= 16'b0000_0000_0000_0000;
array[23735] <= 16'b0000_0000_0000_0000;
array[23736] <= 16'b0000_0000_0000_0000;
array[23737] <= 16'b0000_0000_0000_0000;
array[23738] <= 16'b0000_0000_0000_0000;
array[23739] <= 16'b0000_0000_0000_0000;
array[23740] <= 16'b0000_0000_0000_0000;
array[23741] <= 16'b0000_0000_0000_0000;
array[23742] <= 16'b0000_0000_0000_0000;
array[23743] <= 16'b0000_0000_0000_0000;
array[23744] <= 16'b0000_0000_0000_0000;
array[23745] <= 16'b0000_0000_0000_0000;
array[23746] <= 16'b0000_0000_0000_0000;
array[23747] <= 16'b0000_0000_0000_0000;
array[23748] <= 16'b0000_0000_0000_0000;
array[23749] <= 16'b0000_0000_0000_0000;
array[23750] <= 16'b0000_0000_0000_0000;
array[23751] <= 16'b0000_0000_0000_0000;
array[23752] <= 16'b0000_0000_0000_0000;
array[23753] <= 16'b0000_0000_0000_0000;
array[23754] <= 16'b0000_0000_0000_0000;
array[23755] <= 16'b0000_0000_0000_0000;
array[23756] <= 16'b0000_0000_0000_0000;
array[23757] <= 16'b0000_0000_0000_0000;
array[23758] <= 16'b0000_0000_0000_0000;
array[23759] <= 16'b0000_0000_0000_0000;
array[23760] <= 16'b0000_0000_0000_0000;
array[23761] <= 16'b0000_0000_0000_0000;
array[23762] <= 16'b0000_0000_0000_0000;
array[23763] <= 16'b0000_0000_0000_0000;
array[23764] <= 16'b0000_0000_0000_0000;
array[23765] <= 16'b0000_0000_0000_0000;
array[23766] <= 16'b0000_0000_0000_0000;
array[23767] <= 16'b0000_0000_0000_0000;
array[23768] <= 16'b0000_0000_0000_0000;
array[23769] <= 16'b0000_0000_0000_0000;
array[23770] <= 16'b0000_0000_0000_0000;
array[23771] <= 16'b0000_0000_0000_0000;
array[23772] <= 16'b0000_0000_0000_0000;
array[23773] <= 16'b0000_0000_0000_0000;
array[23774] <= 16'b0000_0000_0000_0000;
array[23775] <= 16'b0000_0000_0000_0000;
array[23776] <= 16'b0000_0000_0000_0000;
array[23777] <= 16'b0000_0000_0000_0000;
array[23778] <= 16'b0000_0000_0000_0000;
array[23779] <= 16'b0000_0000_0000_0000;
array[23780] <= 16'b0000_0000_0000_0000;
array[23781] <= 16'b0000_0000_0000_0000;
array[23782] <= 16'b0000_0000_0000_0000;
array[23783] <= 16'b0000_0000_0000_0000;
array[23784] <= 16'b0000_0000_0000_0000;
array[23785] <= 16'b0000_0000_0000_0000;
array[23786] <= 16'b0000_0000_0000_0000;
array[23787] <= 16'b0000_0000_0000_0000;
array[23788] <= 16'b0000_0000_0000_0000;
array[23789] <= 16'b0000_0000_0000_0000;
array[23790] <= 16'b0000_0000_0000_0000;
array[23791] <= 16'b0000_0000_0000_0000;
array[23792] <= 16'b0000_0000_0000_0000;
array[23793] <= 16'b0000_0000_0000_0000;
array[23794] <= 16'b0000_0000_0000_0000;
array[23795] <= 16'b0000_0000_0000_0000;
array[23796] <= 16'b0000_0000_0000_0000;
array[23797] <= 16'b0000_0000_0000_0000;
array[23798] <= 16'b0000_0000_0000_0000;
array[23799] <= 16'b0000_0000_0000_0000;
array[23800] <= 16'b0000_0000_0000_0000;
array[23801] <= 16'b0000_0000_0000_0000;
array[23802] <= 16'b0000_0000_0000_0000;
array[23803] <= 16'b0000_0000_0000_0000;
array[23804] <= 16'b0000_0000_0000_0000;
array[23805] <= 16'b0000_0000_0000_0000;
array[23806] <= 16'b0000_0000_0000_0000;
array[23807] <= 16'b0000_0000_0000_0000;
array[23808] <= 16'b0000_0000_0000_0000;
array[23809] <= 16'b0000_0000_0000_0000;
array[23810] <= 16'b0000_0000_0000_0000;
array[23811] <= 16'b0000_0000_0000_0000;
array[23812] <= 16'b0000_0000_0000_0000;
array[23813] <= 16'b0000_0000_0000_0000;
array[23814] <= 16'b0000_0000_0000_0000;
array[23815] <= 16'b0000_0000_0000_0000;
array[23816] <= 16'b0000_0000_0000_0000;
array[23817] <= 16'b0000_0000_0000_0000;
array[23818] <= 16'b0000_0000_0000_0000;
array[23819] <= 16'b0000_0000_0000_0000;
array[23820] <= 16'b0000_0000_0000_0000;
array[23821] <= 16'b0000_0000_0000_0000;
array[23822] <= 16'b0000_0000_0000_0000;
array[23823] <= 16'b0000_0000_0000_0000;
array[23824] <= 16'b0000_0000_0000_0000;
array[23825] <= 16'b0000_0000_0000_0000;
array[23826] <= 16'b0000_0000_0000_0000;
array[23827] <= 16'b0000_0000_0000_0000;
array[23828] <= 16'b0000_0000_0000_0000;
array[23829] <= 16'b0000_0000_0000_0000;
array[23830] <= 16'b0000_0000_0000_0000;
array[23831] <= 16'b0000_0000_0000_0000;
array[23832] <= 16'b0000_0000_0000_0000;
array[23833] <= 16'b0000_0000_0000_0000;
array[23834] <= 16'b0000_0000_0000_0000;
array[23835] <= 16'b0000_0000_0000_0000;
array[23836] <= 16'b0000_0000_0000_0000;
array[23837] <= 16'b0000_0000_0000_0000;
array[23838] <= 16'b0000_0000_0000_0000;
array[23839] <= 16'b0000_0000_0000_0000;
array[23840] <= 16'b0000_0000_0000_0000;
array[23841] <= 16'b0000_0000_0000_0000;
array[23842] <= 16'b0000_0000_0000_0000;
array[23843] <= 16'b0000_0000_0000_0000;
array[23844] <= 16'b0000_0000_0000_0000;
array[23845] <= 16'b0000_0000_0000_0000;
array[23846] <= 16'b0000_0000_0000_0000;
array[23847] <= 16'b0000_0000_0000_0000;
array[23848] <= 16'b0000_0000_0000_0000;
array[23849] <= 16'b0000_0000_0000_0000;
array[23850] <= 16'b0000_0000_0000_0000;
array[23851] <= 16'b0000_0000_0000_0000;
array[23852] <= 16'b0000_0000_0000_0000;
array[23853] <= 16'b0000_0000_0000_0000;
array[23854] <= 16'b0000_0000_0000_0000;
array[23855] <= 16'b0000_0000_0000_0000;
array[23856] <= 16'b0000_0000_0000_0000;
array[23857] <= 16'b0000_0000_0000_0000;
array[23858] <= 16'b0000_0000_0000_0000;
array[23859] <= 16'b0000_0000_0000_0000;
array[23860] <= 16'b0000_0000_0000_0000;
array[23861] <= 16'b0000_0000_0000_0000;
array[23862] <= 16'b0000_0000_0000_0000;
array[23863] <= 16'b0000_0000_0000_0000;
array[23864] <= 16'b0000_0000_0000_0000;
array[23865] <= 16'b0000_0000_0000_0000;
array[23866] <= 16'b0000_0000_0000_0000;
array[23867] <= 16'b0000_0000_0000_0000;
array[23868] <= 16'b0000_0000_0000_0000;
array[23869] <= 16'b0000_0000_0000_0000;
array[23870] <= 16'b0000_0000_0000_0000;
array[23871] <= 16'b0000_0000_0000_0000;
array[23872] <= 16'b0000_0000_0000_0000;
array[23873] <= 16'b0000_0000_0000_0000;
array[23874] <= 16'b0000_0000_0000_0000;
array[23875] <= 16'b0000_0000_0000_0000;
array[23876] <= 16'b0000_0000_0000_0000;
array[23877] <= 16'b0000_0000_0000_0000;
array[23878] <= 16'b0000_0000_0000_0000;
array[23879] <= 16'b0000_0000_0000_0000;
array[23880] <= 16'b0000_0000_0000_0000;
array[23881] <= 16'b0000_0000_0000_0000;
array[23882] <= 16'b0000_0000_0000_0000;
array[23883] <= 16'b0000_0000_0000_0000;
array[23884] <= 16'b0000_0000_0000_0000;
array[23885] <= 16'b0000_0000_0000_0000;
array[23886] <= 16'b0000_0000_0000_0000;
array[23887] <= 16'b0000_0000_0000_0000;
array[23888] <= 16'b0000_0000_0000_0000;
array[23889] <= 16'b0000_0000_0000_0000;
array[23890] <= 16'b0000_0000_0000_0000;
array[23891] <= 16'b0000_0000_0000_0000;
array[23892] <= 16'b0000_0000_0000_0000;
array[23893] <= 16'b0000_0000_0000_0000;
array[23894] <= 16'b0000_0000_0000_0000;
array[23895] <= 16'b0000_0000_0000_0000;
array[23896] <= 16'b0000_0000_0000_0000;
array[23897] <= 16'b0000_0000_0000_0000;
array[23898] <= 16'b0000_0000_0000_0000;
array[23899] <= 16'b0000_0000_0000_0000;
array[23900] <= 16'b0000_0000_0000_0000;
array[23901] <= 16'b0000_0000_0000_0000;
array[23902] <= 16'b0000_0000_0000_0000;
array[23903] <= 16'b0000_0000_0000_0000;
array[23904] <= 16'b0000_0000_0000_0000;
array[23905] <= 16'b0000_0000_0000_0000;
array[23906] <= 16'b0000_0000_0000_0000;
array[23907] <= 16'b0000_0000_0000_0000;
array[23908] <= 16'b0000_0000_0000_0000;
array[23909] <= 16'b0000_0000_0000_0000;
array[23910] <= 16'b0000_0000_0000_0000;
array[23911] <= 16'b0000_0000_0000_0000;
array[23912] <= 16'b0000_0000_0000_0000;
array[23913] <= 16'b0000_0000_0000_0000;
array[23914] <= 16'b0000_0000_0000_0000;
array[23915] <= 16'b0000_0000_0000_0000;
array[23916] <= 16'b0000_0000_0000_0000;
array[23917] <= 16'b0000_0000_0000_0000;
array[23918] <= 16'b0000_0000_0000_0000;
array[23919] <= 16'b0000_0000_0000_0000;
array[23920] <= 16'b0000_0000_0000_0000;
array[23921] <= 16'b0000_0000_0000_0000;
array[23922] <= 16'b0000_0000_0000_0000;
array[23923] <= 16'b0000_0000_0000_0000;
array[23924] <= 16'b0000_0000_0000_0000;
array[23925] <= 16'b0000_0000_0000_0000;
array[23926] <= 16'b0000_0000_0000_0000;
array[23927] <= 16'b0000_0000_0000_0000;
array[23928] <= 16'b0000_0000_0000_0000;
array[23929] <= 16'b0000_0000_0000_0000;
array[23930] <= 16'b0000_0000_0000_0000;
array[23931] <= 16'b0000_0000_0000_0000;
array[23932] <= 16'b0000_0000_0000_0000;
array[23933] <= 16'b0000_0000_0000_0000;
array[23934] <= 16'b0000_0000_0000_0000;
array[23935] <= 16'b0000_0000_0000_0000;
array[23936] <= 16'b0000_0000_0000_0000;
array[23937] <= 16'b0000_0000_0000_0000;
array[23938] <= 16'b0000_0000_0000_0000;
array[23939] <= 16'b0000_0000_0000_0000;
array[23940] <= 16'b0000_0000_0000_0000;
array[23941] <= 16'b0000_0000_0000_0000;
array[23942] <= 16'b0000_0000_0000_0000;
array[23943] <= 16'b0000_0000_0000_0000;
array[23944] <= 16'b0000_0000_0000_0000;
array[23945] <= 16'b0000_0000_0000_0000;
array[23946] <= 16'b0000_0000_0000_0000;
array[23947] <= 16'b0000_0000_0000_0000;
array[23948] <= 16'b0000_0000_0000_0000;
array[23949] <= 16'b0000_0000_0000_0000;
array[23950] <= 16'b0000_0000_0000_0000;
array[23951] <= 16'b0000_0000_0000_0000;
array[23952] <= 16'b0000_0000_0000_0000;
array[23953] <= 16'b0000_0000_0000_0000;
array[23954] <= 16'b0000_0000_0000_0000;
array[23955] <= 16'b0000_0000_0000_0000;
array[23956] <= 16'b0000_0000_0000_0000;
array[23957] <= 16'b0000_0000_0000_0000;
array[23958] <= 16'b0000_0000_0000_0000;
array[23959] <= 16'b0000_0000_0000_0000;
array[23960] <= 16'b0000_0000_0000_0000;
array[23961] <= 16'b0000_0000_0000_0000;
array[23962] <= 16'b0000_0000_0000_0000;
array[23963] <= 16'b0000_0000_0000_0000;
array[23964] <= 16'b0000_0000_0000_0000;
array[23965] <= 16'b0000_0000_0000_0000;
array[23966] <= 16'b0000_0000_0000_0000;
array[23967] <= 16'b0000_0000_0000_0000;
array[23968] <= 16'b0000_0000_0000_0000;
array[23969] <= 16'b0000_0000_0000_0000;
array[23970] <= 16'b0000_0000_0000_0000;
array[23971] <= 16'b0000_0000_0000_0000;
array[23972] <= 16'b0000_0000_0000_0000;
array[23973] <= 16'b0000_0000_0000_0000;
array[23974] <= 16'b0000_0000_0000_0000;
array[23975] <= 16'b0000_0000_0000_0000;
array[23976] <= 16'b0000_0000_0000_0000;
array[23977] <= 16'b0000_0000_0000_0000;
array[23978] <= 16'b0000_0000_0000_0000;
array[23979] <= 16'b0000_0000_0000_0000;
array[23980] <= 16'b0000_0000_0000_0000;
array[23981] <= 16'b0000_0000_0000_0000;
array[23982] <= 16'b0000_0000_0000_0000;
array[23983] <= 16'b0000_0000_0000_0000;
array[23984] <= 16'b0000_0000_0000_0000;
array[23985] <= 16'b0000_0000_0000_0000;
array[23986] <= 16'b0000_0000_0000_0000;
array[23987] <= 16'b0000_0000_0000_0000;
array[23988] <= 16'b0000_0000_0000_0000;
array[23989] <= 16'b0000_0000_0000_0000;
array[23990] <= 16'b0000_0000_0000_0000;
array[23991] <= 16'b0000_0000_0000_0000;
array[23992] <= 16'b0000_0000_0000_0000;
array[23993] <= 16'b0000_0000_0000_0000;
array[23994] <= 16'b0000_0000_0000_0000;
array[23995] <= 16'b0000_0000_0000_0000;
array[23996] <= 16'b0000_0000_0000_0000;
array[23997] <= 16'b0000_0000_0000_0000;
array[23998] <= 16'b0000_0000_0000_0000;
array[23999] <= 16'b0000_0000_0000_0000;
array[24000] <= 16'b0000_0000_0000_0000;
array[24001] <= 16'b0000_0000_0000_0000;
array[24002] <= 16'b0000_0000_0000_0000;
array[24003] <= 16'b0000_0000_0000_0000;
array[24004] <= 16'b0000_0000_0000_0000;
array[24005] <= 16'b0000_0000_0000_0000;
array[24006] <= 16'b0000_0000_0000_0000;
array[24007] <= 16'b0000_0000_0000_0000;
array[24008] <= 16'b0000_0000_0000_0000;
array[24009] <= 16'b0000_0000_0000_0000;
array[24010] <= 16'b0000_0000_0000_0000;
array[24011] <= 16'b0000_0000_0000_0000;
array[24012] <= 16'b0000_0000_0000_0000;
array[24013] <= 16'b0000_0000_0000_0000;
array[24014] <= 16'b0000_0000_0000_0000;
array[24015] <= 16'b0000_0000_0000_0000;
array[24016] <= 16'b0000_0000_0000_0000;
array[24017] <= 16'b0000_0000_0000_0000;
array[24018] <= 16'b0000_0000_0000_0000;
array[24019] <= 16'b0000_0000_0000_0000;
array[24020] <= 16'b0000_0000_0000_0000;
array[24021] <= 16'b0000_0000_0000_0000;
array[24022] <= 16'b0000_0000_0000_0000;
array[24023] <= 16'b0000_0000_0000_0000;
array[24024] <= 16'b0000_0000_0000_0000;
array[24025] <= 16'b0000_0000_0000_0000;
array[24026] <= 16'b0000_0000_0000_0000;
array[24027] <= 16'b0000_0000_0000_0000;
array[24028] <= 16'b0000_0000_0000_0000;
array[24029] <= 16'b0000_0000_0000_0000;
array[24030] <= 16'b0000_0000_0000_0000;
array[24031] <= 16'b0000_0000_0000_0000;
array[24032] <= 16'b0000_0000_0000_0000;
array[24033] <= 16'b0000_0000_0000_0000;
array[24034] <= 16'b0000_0000_0000_0000;
array[24035] <= 16'b0000_0000_0000_0000;
array[24036] <= 16'b0000_0000_0000_0000;
array[24037] <= 16'b0000_0000_0000_0000;
array[24038] <= 16'b0000_0000_0000_0000;
array[24039] <= 16'b0000_0000_0000_0000;
array[24040] <= 16'b0000_0000_0000_0000;
array[24041] <= 16'b0000_0000_0000_0000;
array[24042] <= 16'b0000_0000_0000_0000;
array[24043] <= 16'b0000_0000_0000_0000;
array[24044] <= 16'b0000_0000_0000_0000;
array[24045] <= 16'b0000_0000_0000_0000;
array[24046] <= 16'b0000_0000_0000_0000;
array[24047] <= 16'b0000_0000_0000_0000;
array[24048] <= 16'b0000_0000_0000_0000;
array[24049] <= 16'b0000_0000_0000_0000;
array[24050] <= 16'b0000_0000_0000_0000;
array[24051] <= 16'b0000_0000_0000_0000;
array[24052] <= 16'b0000_0000_0000_0000;
array[24053] <= 16'b0000_0000_0000_0000;
array[24054] <= 16'b0000_0000_0000_0000;
array[24055] <= 16'b0000_0000_0000_0000;
array[24056] <= 16'b0000_0000_0000_0000;
array[24057] <= 16'b0000_0000_0000_0000;
array[24058] <= 16'b0000_0000_0000_0000;
array[24059] <= 16'b0000_0000_0000_0000;
array[24060] <= 16'b0000_0000_0000_0000;
array[24061] <= 16'b0000_0000_0000_0000;
array[24062] <= 16'b0000_0000_0000_0000;
array[24063] <= 16'b0000_0000_0000_0000;
array[24064] <= 16'b0000_0000_0000_0000;
array[24065] <= 16'b0000_0000_0000_0000;
array[24066] <= 16'b0000_0000_0000_0000;
array[24067] <= 16'b0000_0000_0000_0000;
array[24068] <= 16'b0000_0000_0000_0000;
array[24069] <= 16'b0000_0000_0000_0000;
array[24070] <= 16'b0000_0000_0000_0000;
array[24071] <= 16'b0000_0000_0000_0000;
array[24072] <= 16'b0000_0000_0000_0000;
array[24073] <= 16'b0000_0000_0000_0000;
array[24074] <= 16'b0000_0000_0000_0000;
array[24075] <= 16'b0000_0000_0000_0000;
array[24076] <= 16'b0000_0000_0000_0000;
array[24077] <= 16'b0000_0000_0000_0000;
array[24078] <= 16'b0000_0000_0000_0000;
array[24079] <= 16'b0000_0000_0000_0000;
array[24080] <= 16'b0000_0000_0000_0000;
array[24081] <= 16'b0000_0000_0000_0000;
array[24082] <= 16'b0000_0000_0000_0000;
array[24083] <= 16'b0000_0000_0000_0000;
array[24084] <= 16'b0000_0000_0000_0000;
array[24085] <= 16'b0000_0000_0000_0000;
array[24086] <= 16'b0000_0000_0000_0000;
array[24087] <= 16'b0000_0000_0000_0000;
array[24088] <= 16'b0000_0000_0000_0000;
array[24089] <= 16'b0000_0000_0000_0000;
array[24090] <= 16'b0000_0000_0000_0000;
array[24091] <= 16'b0000_0000_0000_0000;
array[24092] <= 16'b0000_0000_0000_0000;
array[24093] <= 16'b0000_0000_0000_0000;
array[24094] <= 16'b0000_0000_0000_0000;
array[24095] <= 16'b0000_0000_0000_0000;
array[24096] <= 16'b0000_0000_0000_0000;
array[24097] <= 16'b0000_0000_0000_0000;
array[24098] <= 16'b0000_0000_0000_0000;
array[24099] <= 16'b0000_0000_0000_0000;
array[24100] <= 16'b0000_0000_0000_0000;
array[24101] <= 16'b0000_0000_0000_0000;
array[24102] <= 16'b0000_0000_0000_0000;
array[24103] <= 16'b0000_0000_0000_0000;
array[24104] <= 16'b0000_0000_0000_0000;
array[24105] <= 16'b0000_0000_0000_0000;
array[24106] <= 16'b0000_0000_0000_0000;
array[24107] <= 16'b0000_0000_0000_0000;
array[24108] <= 16'b0000_0000_0000_0000;
array[24109] <= 16'b0000_0000_0000_0000;
array[24110] <= 16'b0000_0000_0000_0000;
array[24111] <= 16'b0000_0000_0000_0000;
array[24112] <= 16'b0000_0000_0000_0000;
array[24113] <= 16'b0000_0000_0000_0000;
array[24114] <= 16'b0000_0000_0000_0000;
array[24115] <= 16'b0000_0000_0000_0000;
array[24116] <= 16'b0000_0000_0000_0000;
array[24117] <= 16'b0000_0000_0000_0000;
array[24118] <= 16'b0000_0000_0000_0000;
array[24119] <= 16'b0000_0000_0000_0000;
array[24120] <= 16'b0000_0000_0000_0000;
array[24121] <= 16'b0000_0000_0000_0000;
array[24122] <= 16'b0000_0000_0000_0000;
array[24123] <= 16'b0000_0000_0000_0000;
array[24124] <= 16'b0000_0000_0000_0000;
array[24125] <= 16'b0000_0000_0000_0000;
array[24126] <= 16'b0000_0000_0000_0000;
array[24127] <= 16'b0000_0000_0000_0000;
array[24128] <= 16'b0000_0000_0000_0000;
array[24129] <= 16'b0000_0000_0000_0000;
array[24130] <= 16'b0000_0000_0000_0000;
array[24131] <= 16'b0000_0000_0000_0000;
array[24132] <= 16'b0000_0000_0000_0000;
array[24133] <= 16'b0000_0000_0000_0000;
array[24134] <= 16'b0000_0000_0000_0000;
array[24135] <= 16'b0000_0000_0000_0000;
array[24136] <= 16'b0000_0000_0000_0000;
array[24137] <= 16'b0000_0000_0000_0000;
array[24138] <= 16'b0000_0000_0000_0000;
array[24139] <= 16'b0000_0000_0000_0000;
array[24140] <= 16'b0000_0000_0000_0000;
array[24141] <= 16'b0000_0000_0000_0000;
array[24142] <= 16'b0000_0000_0000_0000;
array[24143] <= 16'b0000_0000_0000_0000;
array[24144] <= 16'b0000_0000_0000_0000;
array[24145] <= 16'b0000_0000_0000_0000;
array[24146] <= 16'b0000_0000_0000_0000;
array[24147] <= 16'b0000_0000_0000_0000;
array[24148] <= 16'b0000_0000_0000_0000;
array[24149] <= 16'b0000_0000_0000_0000;
array[24150] <= 16'b0000_0000_0000_0000;
array[24151] <= 16'b0000_0000_0000_0000;
array[24152] <= 16'b0000_0000_0000_0000;
array[24153] <= 16'b0000_0000_0000_0000;
array[24154] <= 16'b0000_0000_0000_0000;
array[24155] <= 16'b0000_0000_0000_0000;
array[24156] <= 16'b0000_0000_0000_0000;
array[24157] <= 16'b0000_0000_0000_0000;
array[24158] <= 16'b0000_0000_0000_0000;
array[24159] <= 16'b0000_0000_0000_0000;
array[24160] <= 16'b0000_0000_0000_0000;
array[24161] <= 16'b0000_0000_0000_0000;
array[24162] <= 16'b0000_0000_0000_0000;
array[24163] <= 16'b0000_0000_0000_0000;
array[24164] <= 16'b0000_0000_0000_0000;
array[24165] <= 16'b0000_0000_0000_0000;
array[24166] <= 16'b0000_0000_0000_0000;
array[24167] <= 16'b0000_0000_0000_0000;
array[24168] <= 16'b0000_0000_0000_0000;
array[24169] <= 16'b0000_0000_0000_0000;
array[24170] <= 16'b0000_0000_0000_0000;
array[24171] <= 16'b0000_0000_0000_0000;
array[24172] <= 16'b0000_0000_0000_0000;
array[24173] <= 16'b0000_0000_0000_0000;
array[24174] <= 16'b0000_0000_0000_0000;
array[24175] <= 16'b0000_0000_0000_0000;
array[24176] <= 16'b0000_0000_0000_0000;
array[24177] <= 16'b0000_0000_0000_0000;
array[24178] <= 16'b0000_0000_0000_0000;
array[24179] <= 16'b0000_0000_0000_0000;
array[24180] <= 16'b0000_0000_0000_0000;
array[24181] <= 16'b0000_0000_0000_0000;
array[24182] <= 16'b0000_0000_0000_0000;
array[24183] <= 16'b0000_0000_0000_0000;
array[24184] <= 16'b0000_0000_0000_0000;
array[24185] <= 16'b0000_0000_0000_0000;
array[24186] <= 16'b0000_0000_0000_0000;
array[24187] <= 16'b0000_0000_0000_0000;
array[24188] <= 16'b0000_0000_0000_0000;
array[24189] <= 16'b0000_0000_0000_0000;
array[24190] <= 16'b0000_0000_0000_0000;
array[24191] <= 16'b0000_0000_0000_0000;
array[24192] <= 16'b0000_0000_0000_0000;
array[24193] <= 16'b0000_0000_0000_0000;
array[24194] <= 16'b0000_0000_0000_0000;
array[24195] <= 16'b0000_0000_0000_0000;
array[24196] <= 16'b0000_0000_0000_0000;
array[24197] <= 16'b0000_0000_0000_0000;
array[24198] <= 16'b0000_0000_0000_0000;
array[24199] <= 16'b0000_0000_0000_0000;
array[24200] <= 16'b0000_0000_0000_0000;
array[24201] <= 16'b0000_0000_0000_0000;
array[24202] <= 16'b0000_0000_0000_0000;
array[24203] <= 16'b0000_0000_0000_0000;
array[24204] <= 16'b0000_0000_0000_0000;
array[24205] <= 16'b0000_0000_0000_0000;
array[24206] <= 16'b0000_0000_0000_0000;
array[24207] <= 16'b0000_0000_0000_0000;
array[24208] <= 16'b0000_0000_0000_0000;
array[24209] <= 16'b0000_0000_0000_0000;
array[24210] <= 16'b0000_0000_0000_0000;
array[24211] <= 16'b0000_0000_0000_0000;
array[24212] <= 16'b0000_0000_0000_0000;
array[24213] <= 16'b0000_0000_0000_0000;
array[24214] <= 16'b0000_0000_0000_0000;
array[24215] <= 16'b0000_0000_0000_0000;
array[24216] <= 16'b0000_0000_0000_0000;
array[24217] <= 16'b0000_0000_0000_0000;
array[24218] <= 16'b0000_0000_0000_0000;
array[24219] <= 16'b0000_0000_0000_0000;
array[24220] <= 16'b0000_0000_0000_0000;
array[24221] <= 16'b0000_0000_0000_0000;
array[24222] <= 16'b0000_0000_0000_0000;
array[24223] <= 16'b0000_0000_0000_0000;
array[24224] <= 16'b0000_0000_0000_0000;
array[24225] <= 16'b0000_0000_0000_0000;
array[24226] <= 16'b0000_0000_0000_0000;
array[24227] <= 16'b0000_0000_0000_0000;
array[24228] <= 16'b0000_0000_0000_0000;
array[24229] <= 16'b0000_0000_0000_0000;
array[24230] <= 16'b0000_0000_0000_0000;
array[24231] <= 16'b0000_0000_0000_0000;
array[24232] <= 16'b0000_0000_0000_0000;
array[24233] <= 16'b0000_0000_0000_0000;
array[24234] <= 16'b0000_0000_0000_0000;
array[24235] <= 16'b0000_0000_0000_0000;
array[24236] <= 16'b0000_0000_0000_0000;
array[24237] <= 16'b0000_0000_0000_0000;
array[24238] <= 16'b0000_0000_0000_0000;
array[24239] <= 16'b0000_0000_0000_0000;
array[24240] <= 16'b0000_0000_0000_0000;
array[24241] <= 16'b0000_0000_0000_0000;
array[24242] <= 16'b0000_0000_0000_0000;
array[24243] <= 16'b0000_0000_0000_0000;
array[24244] <= 16'b0000_0000_0000_0000;
array[24245] <= 16'b0000_0000_0000_0000;
array[24246] <= 16'b0000_0000_0000_0000;
array[24247] <= 16'b0000_0000_0000_0000;
array[24248] <= 16'b0000_0000_0000_0000;
array[24249] <= 16'b0000_0000_0000_0000;
array[24250] <= 16'b0000_0000_0000_0000;
array[24251] <= 16'b0000_0000_0000_0000;
array[24252] <= 16'b0000_0000_0000_0000;
array[24253] <= 16'b0000_0000_0000_0000;
array[24254] <= 16'b0000_0000_0000_0000;
array[24255] <= 16'b0000_0000_0000_0000;
array[24256] <= 16'b0000_0000_0000_0000;
array[24257] <= 16'b0000_0000_0000_0000;
array[24258] <= 16'b0000_0000_0000_0000;
array[24259] <= 16'b0000_0000_0000_0000;
array[24260] <= 16'b0000_0000_0000_0000;
array[24261] <= 16'b0000_0000_0000_0000;
array[24262] <= 16'b0000_0000_0000_0000;
array[24263] <= 16'b0000_0000_0000_0000;
array[24264] <= 16'b0000_0000_0000_0000;
array[24265] <= 16'b0000_0000_0000_0000;
array[24266] <= 16'b0000_0000_0000_0000;
array[24267] <= 16'b0000_0000_0000_0000;
array[24268] <= 16'b0000_0000_0000_0000;
array[24269] <= 16'b0000_0000_0000_0000;
array[24270] <= 16'b0000_0000_0000_0000;
array[24271] <= 16'b0000_0000_0000_0000;
array[24272] <= 16'b0000_0000_0000_0000;
array[24273] <= 16'b0000_0000_0000_0000;
array[24274] <= 16'b0000_0000_0000_0000;
array[24275] <= 16'b0000_0000_0000_0000;
array[24276] <= 16'b0000_0000_0000_0000;
array[24277] <= 16'b0000_0000_0000_0000;
array[24278] <= 16'b0000_0000_0000_0000;
array[24279] <= 16'b0000_0000_0000_0000;
array[24280] <= 16'b0000_0000_0000_0000;
array[24281] <= 16'b0000_0000_0000_0000;
array[24282] <= 16'b0000_0000_0000_0000;
array[24283] <= 16'b0000_0000_0000_0000;
array[24284] <= 16'b0000_0000_0000_0000;
array[24285] <= 16'b0000_0000_0000_0000;
array[24286] <= 16'b0000_0000_0000_0000;
array[24287] <= 16'b0000_0000_0000_0000;
array[24288] <= 16'b0000_0000_0000_0000;
array[24289] <= 16'b0000_0000_0000_0000;
array[24290] <= 16'b0000_0000_0000_0000;
array[24291] <= 16'b0000_0000_0000_0000;
array[24292] <= 16'b0000_0000_0000_0000;
array[24293] <= 16'b0000_0000_0000_0000;
array[24294] <= 16'b0000_0000_0000_0000;
array[24295] <= 16'b0000_0000_0000_0000;
array[24296] <= 16'b0000_0000_0000_0000;
array[24297] <= 16'b0000_0000_0000_0000;
array[24298] <= 16'b0000_0000_0000_0000;
array[24299] <= 16'b0000_0000_0000_0000;
array[24300] <= 16'b0000_0000_0000_0000;
array[24301] <= 16'b0000_0000_0000_0000;
array[24302] <= 16'b0000_0000_0000_0000;
array[24303] <= 16'b0000_0000_0000_0000;
array[24304] <= 16'b0000_0000_0000_0000;
array[24305] <= 16'b0000_0000_0000_0000;
array[24306] <= 16'b0000_0000_0000_0000;
array[24307] <= 16'b0000_0000_0000_0000;
array[24308] <= 16'b0000_0000_0000_0000;
array[24309] <= 16'b0000_0000_0000_0000;
array[24310] <= 16'b0000_0000_0000_0000;
array[24311] <= 16'b0000_0000_0000_0000;
array[24312] <= 16'b0000_0000_0000_0000;
array[24313] <= 16'b0000_0000_0000_0000;
array[24314] <= 16'b0000_0000_0000_0000;
array[24315] <= 16'b0000_0000_0000_0000;
array[24316] <= 16'b0000_0000_0000_0000;
array[24317] <= 16'b0000_0000_0000_0000;
array[24318] <= 16'b0000_0000_0000_0000;
array[24319] <= 16'b0000_0000_0000_0000;
array[24320] <= 16'b0000_0000_0000_0000;
array[24321] <= 16'b0000_0000_0000_0000;
array[24322] <= 16'b0000_0000_0000_0000;
array[24323] <= 16'b0000_0000_0000_0000;
array[24324] <= 16'b0000_0000_0000_0000;
array[24325] <= 16'b0000_0000_0000_0000;
array[24326] <= 16'b0000_0000_0000_0000;
array[24327] <= 16'b0000_0000_0000_0000;
array[24328] <= 16'b0000_0000_0000_0000;
array[24329] <= 16'b0000_0000_0000_0000;
array[24330] <= 16'b0000_0000_0000_0000;
array[24331] <= 16'b0000_0000_0000_0000;
array[24332] <= 16'b0000_0000_0000_0000;
array[24333] <= 16'b0000_0000_0000_0000;
array[24334] <= 16'b0000_0000_0000_0000;
array[24335] <= 16'b0000_0000_0000_0000;
array[24336] <= 16'b0000_0000_0000_0000;
array[24337] <= 16'b0000_0000_0000_0000;
array[24338] <= 16'b0000_0000_0000_0000;
array[24339] <= 16'b0000_0000_0000_0000;
array[24340] <= 16'b0000_0000_0000_0000;
array[24341] <= 16'b0000_0000_0000_0000;
array[24342] <= 16'b0000_0000_0000_0000;
array[24343] <= 16'b0000_0000_0000_0000;
array[24344] <= 16'b0000_0000_0000_0000;
array[24345] <= 16'b0000_0000_0000_0000;
array[24346] <= 16'b0000_0000_0000_0000;
array[24347] <= 16'b0000_0000_0000_0000;
array[24348] <= 16'b0000_0000_0000_0000;
array[24349] <= 16'b0000_0000_0000_0000;
array[24350] <= 16'b0000_0000_0000_0000;
array[24351] <= 16'b0000_0000_0000_0000;
array[24352] <= 16'b0000_0000_0000_0000;
array[24353] <= 16'b0000_0000_0000_0000;
array[24354] <= 16'b0000_0000_0000_0000;
array[24355] <= 16'b0000_0000_0000_0000;
array[24356] <= 16'b0000_0000_0000_0000;
array[24357] <= 16'b0000_0000_0000_0000;
array[24358] <= 16'b0000_0000_0000_0000;
array[24359] <= 16'b0000_0000_0000_0000;
array[24360] <= 16'b0000_0000_0000_0000;
array[24361] <= 16'b0000_0000_0000_0000;
array[24362] <= 16'b0000_0000_0000_0000;
array[24363] <= 16'b0000_0000_0000_0000;
array[24364] <= 16'b0000_0000_0000_0000;
array[24365] <= 16'b0000_0000_0000_0000;
array[24366] <= 16'b0000_0000_0000_0000;
array[24367] <= 16'b0000_0000_0000_0000;
array[24368] <= 16'b0000_0000_0000_0000;
array[24369] <= 16'b0000_0000_0000_0000;
array[24370] <= 16'b0000_0000_0000_0000;
array[24371] <= 16'b0000_0000_0000_0000;
array[24372] <= 16'b0000_0000_0000_0000;
array[24373] <= 16'b0000_0000_0000_0000;
array[24374] <= 16'b0000_0000_0000_0000;
array[24375] <= 16'b0000_0000_0000_0000;
array[24376] <= 16'b0000_0000_0000_0000;
array[24377] <= 16'b0000_0000_0000_0000;
array[24378] <= 16'b0000_0000_0000_0000;
array[24379] <= 16'b0000_0000_0000_0000;
array[24380] <= 16'b0000_0000_0000_0000;
array[24381] <= 16'b0000_0000_0000_0000;
array[24382] <= 16'b0000_0000_0000_0000;
array[24383] <= 16'b0000_0000_0000_0000;
array[24384] <= 16'b0000_0000_0000_0000;
array[24385] <= 16'b0000_0000_0000_0000;
array[24386] <= 16'b0000_0000_0000_0000;
array[24387] <= 16'b0000_0000_0000_0000;
array[24388] <= 16'b0000_0000_0000_0000;
array[24389] <= 16'b0000_0000_0000_0000;
array[24390] <= 16'b0000_0000_0000_0000;
array[24391] <= 16'b0000_0000_0000_0000;
array[24392] <= 16'b0000_0000_0000_0000;
array[24393] <= 16'b0000_0000_0000_0000;
array[24394] <= 16'b0000_0000_0000_0000;
array[24395] <= 16'b0000_0000_0000_0000;
array[24396] <= 16'b0000_0000_0000_0000;
array[24397] <= 16'b0000_0000_0000_0000;
array[24398] <= 16'b0000_0000_0000_0000;
array[24399] <= 16'b0000_0000_0000_0000;
array[24400] <= 16'b0000_0000_0000_0000;
array[24401] <= 16'b0000_0000_0000_0000;
array[24402] <= 16'b0000_0000_0000_0000;
array[24403] <= 16'b0000_0000_0000_0000;
array[24404] <= 16'b0000_0000_0000_0000;
array[24405] <= 16'b0000_0000_0000_0000;
array[24406] <= 16'b0000_0000_0000_0000;
array[24407] <= 16'b0000_0000_0000_0000;
array[24408] <= 16'b0000_0000_0000_0000;
array[24409] <= 16'b0000_0000_0000_0000;
array[24410] <= 16'b0000_0000_0000_0000;
array[24411] <= 16'b0000_0000_0000_0000;
array[24412] <= 16'b0000_0000_0000_0000;
array[24413] <= 16'b0000_0000_0000_0000;
array[24414] <= 16'b0000_0000_0000_0000;
array[24415] <= 16'b0000_0000_0000_0000;
array[24416] <= 16'b0000_0000_0000_0000;
array[24417] <= 16'b0000_0000_0000_0000;
array[24418] <= 16'b0000_0000_0000_0000;
array[24419] <= 16'b0000_0000_0000_0000;
array[24420] <= 16'b0000_0000_0000_0000;
array[24421] <= 16'b0000_0000_0000_0000;
array[24422] <= 16'b0000_0000_0000_0000;
array[24423] <= 16'b0000_0000_0000_0000;
array[24424] <= 16'b0000_0000_0000_0000;
array[24425] <= 16'b0000_0000_0000_0000;
array[24426] <= 16'b0000_0000_0000_0000;
array[24427] <= 16'b0000_0000_0000_0000;
array[24428] <= 16'b0000_0000_0000_0000;
array[24429] <= 16'b0000_0000_0000_0000;
array[24430] <= 16'b0000_0000_0000_0000;
array[24431] <= 16'b0000_0000_0000_0000;
array[24432] <= 16'b0000_0000_0000_0000;
array[24433] <= 16'b0000_0000_0000_0000;
array[24434] <= 16'b0000_0000_0000_0000;
array[24435] <= 16'b0000_0000_0000_0000;
array[24436] <= 16'b0000_0000_0000_0000;
array[24437] <= 16'b0000_0000_0000_0000;
array[24438] <= 16'b0000_0000_0000_0000;
array[24439] <= 16'b0000_0000_0000_0000;
array[24440] <= 16'b0000_0000_0000_0000;
array[24441] <= 16'b0000_0000_0000_0000;
array[24442] <= 16'b0000_0000_0000_0000;
array[24443] <= 16'b0000_0000_0000_0000;
array[24444] <= 16'b0000_0000_0000_0000;
array[24445] <= 16'b0000_0000_0000_0000;
array[24446] <= 16'b0000_0000_0000_0000;
array[24447] <= 16'b0000_0000_0000_0000;
array[24448] <= 16'b0000_0000_0000_0000;
array[24449] <= 16'b0000_0000_0000_0000;
array[24450] <= 16'b0000_0000_0000_0000;
array[24451] <= 16'b0000_0000_0000_0000;
array[24452] <= 16'b0000_0000_0000_0000;
array[24453] <= 16'b0000_0000_0000_0000;
array[24454] <= 16'b0000_0000_0000_0000;
array[24455] <= 16'b0000_0000_0000_0000;
array[24456] <= 16'b0000_0000_0000_0000;
array[24457] <= 16'b0000_0000_0000_0000;
array[24458] <= 16'b0000_0000_0000_0000;
array[24459] <= 16'b0000_0000_0000_0000;
array[24460] <= 16'b0000_0000_0000_0000;
array[24461] <= 16'b0000_0000_0000_0000;
array[24462] <= 16'b0000_0000_0000_0000;
array[24463] <= 16'b0000_0000_0000_0000;
array[24464] <= 16'b0000_0000_0000_0000;
array[24465] <= 16'b0000_0000_0000_0000;
array[24466] <= 16'b0000_0000_0000_0000;
array[24467] <= 16'b0000_0000_0000_0000;
array[24468] <= 16'b0000_0000_0000_0000;
array[24469] <= 16'b0000_0000_0000_0000;
array[24470] <= 16'b0000_0000_0000_0000;
array[24471] <= 16'b0000_0000_0000_0000;
array[24472] <= 16'b0000_0000_0000_0000;
array[24473] <= 16'b0000_0000_0000_0000;
array[24474] <= 16'b0000_0000_0000_0000;
array[24475] <= 16'b0000_0000_0000_0000;
array[24476] <= 16'b0000_0000_0000_0000;
array[24477] <= 16'b0000_0000_0000_0000;
array[24478] <= 16'b0000_0000_0000_0000;
array[24479] <= 16'b0000_0000_0000_0000;
array[24480] <= 16'b0000_0000_0000_0000;
array[24481] <= 16'b0000_0000_0000_0000;
array[24482] <= 16'b0000_0000_0000_0000;
array[24483] <= 16'b0000_0000_0000_0000;
array[24484] <= 16'b0000_0000_0000_0000;
array[24485] <= 16'b0000_0000_0000_0000;
array[24486] <= 16'b0000_0000_0000_0000;
array[24487] <= 16'b0000_0000_0000_0000;
array[24488] <= 16'b0000_0000_0000_0000;
array[24489] <= 16'b0000_0000_0000_0000;
array[24490] <= 16'b0000_0000_0000_0000;
array[24491] <= 16'b0000_0000_0000_0000;
array[24492] <= 16'b0000_0000_0000_0000;
array[24493] <= 16'b0000_0000_0000_0000;
array[24494] <= 16'b0000_0000_0000_0000;
array[24495] <= 16'b0000_0000_0000_0000;
array[24496] <= 16'b0000_0000_0000_0000;
array[24497] <= 16'b0000_0000_0000_0000;
array[24498] <= 16'b0000_0000_0000_0000;
array[24499] <= 16'b0000_0000_0000_0000;
array[24500] <= 16'b0000_0000_0000_0000;
array[24501] <= 16'b0000_0000_0000_0000;
array[24502] <= 16'b0000_0000_0000_0000;
array[24503] <= 16'b0000_0000_0000_0000;
array[24504] <= 16'b0000_0000_0000_0000;
array[24505] <= 16'b0000_0000_0000_0000;
array[24506] <= 16'b0000_0000_0000_0000;
array[24507] <= 16'b0000_0000_0000_0000;
array[24508] <= 16'b0000_0000_0000_0000;
array[24509] <= 16'b0000_0000_0000_0000;
array[24510] <= 16'b0000_0000_0000_0000;
array[24511] <= 16'b0000_0000_0000_0000;
array[24512] <= 16'b0000_0000_0000_0000;
array[24513] <= 16'b0000_0000_0000_0000;
array[24514] <= 16'b0000_0000_0000_0000;
array[24515] <= 16'b0000_0000_0000_0000;
array[24516] <= 16'b0000_0000_0000_0000;
array[24517] <= 16'b0000_0000_0000_0000;
array[24518] <= 16'b0000_0000_0000_0000;
array[24519] <= 16'b0000_0000_0000_0000;
array[24520] <= 16'b0000_0000_0000_0000;
array[24521] <= 16'b0000_0000_0000_0000;
array[24522] <= 16'b0000_0000_0000_0000;
array[24523] <= 16'b0000_0000_0000_0000;
array[24524] <= 16'b0000_0000_0000_0000;
array[24525] <= 16'b0000_0000_0000_0000;
array[24526] <= 16'b0000_0000_0000_0000;
array[24527] <= 16'b0000_0000_0000_0000;
array[24528] <= 16'b0000_0000_0000_0000;
array[24529] <= 16'b0000_0000_0000_0000;
array[24530] <= 16'b0000_0000_0000_0000;
array[24531] <= 16'b0000_0000_0000_0000;
array[24532] <= 16'b0000_0000_0000_0000;
array[24533] <= 16'b0000_0000_0000_0000;
array[24534] <= 16'b0000_0000_0000_0000;
array[24535] <= 16'b0000_0000_0000_0000;
array[24536] <= 16'b0000_0000_0000_0000;
array[24537] <= 16'b0000_0000_0000_0000;
array[24538] <= 16'b0000_0000_0000_0000;
array[24539] <= 16'b0000_0000_0000_0000;
array[24540] <= 16'b0000_0000_0000_0000;
array[24541] <= 16'b0000_0000_0000_0000;
array[24542] <= 16'b0000_0000_0000_0000;
array[24543] <= 16'b0000_0000_0000_0000;
array[24544] <= 16'b0000_0000_0000_0000;
array[24545] <= 16'b0000_0000_0000_0000;
array[24546] <= 16'b0000_0000_0000_0000;
array[24547] <= 16'b0000_0000_0000_0000;
array[24548] <= 16'b0000_0000_0000_0000;
array[24549] <= 16'b0000_0000_0000_0000;
array[24550] <= 16'b0000_0000_0000_0000;
array[24551] <= 16'b0000_0000_0000_0000;
array[24552] <= 16'b0000_0000_0000_0000;
array[24553] <= 16'b0000_0000_0000_0000;
array[24554] <= 16'b0000_0000_0000_0000;
array[24555] <= 16'b0000_0000_0000_0000;
array[24556] <= 16'b0000_0000_0000_0000;
array[24557] <= 16'b0000_0000_0000_0000;
array[24558] <= 16'b0000_0000_0000_0000;
array[24559] <= 16'b0000_0000_0000_0000;
array[24560] <= 16'b0000_0000_0000_0000;
array[24561] <= 16'b0000_0000_0000_0000;
array[24562] <= 16'b0000_0000_0000_0000;
array[24563] <= 16'b0000_0000_0000_0000;
array[24564] <= 16'b0000_0000_0000_0000;
array[24565] <= 16'b0000_0000_0000_0000;
array[24566] <= 16'b0000_0000_0000_0000;
array[24567] <= 16'b0000_0000_0000_0000;
array[24568] <= 16'b0000_0000_0000_0000;
array[24569] <= 16'b0000_0000_0000_0000;
array[24570] <= 16'b0000_0000_0000_0000;
array[24571] <= 16'b0000_0000_0000_0000;
array[24572] <= 16'b0000_0000_0000_0000;
array[24573] <= 16'b0000_0000_0000_0000;
array[24574] <= 16'b0000_0000_0000_0000;
array[24575] <= 16'b0000_0000_0000_0000;
array[24576] <= 16'b0000_0000_0000_0000;
array[24577] <= 16'b0000_0000_0000_0000;
array[24578] <= 16'b0000_0000_0000_0000;
array[24579] <= 16'b0000_0000_0000_0000;
array[24580] <= 16'b0000_0000_0000_0000;
array[24581] <= 16'b0000_0000_0000_0000;
array[24582] <= 16'b0000_0000_0000_0000;
array[24583] <= 16'b0000_0000_0000_0000;
array[24584] <= 16'b0000_0000_0000_0000;
array[24585] <= 16'b0000_0000_0000_0000;
array[24586] <= 16'b0000_0000_0000_0000;
array[24587] <= 16'b0000_0000_0000_0000;
array[24588] <= 16'b0000_0000_0000_0000;
array[24589] <= 16'b0000_0000_0000_0000;
array[24590] <= 16'b0000_0000_0000_0000;
array[24591] <= 16'b0000_0000_0000_0000;
array[24592] <= 16'b0000_0000_0000_0000;
array[24593] <= 16'b0000_0000_0000_0000;
array[24594] <= 16'b0000_0000_0000_0000;
array[24595] <= 16'b0000_0000_0000_0000;
array[24596] <= 16'b0000_0000_0000_0000;
array[24597] <= 16'b0000_0000_0000_0000;
array[24598] <= 16'b0000_0000_0000_0000;
array[24599] <= 16'b0000_0000_0000_0000;
array[24600] <= 16'b0000_0000_0000_0000;
array[24601] <= 16'b0000_0000_0000_0000;
array[24602] <= 16'b0000_0000_0000_0000;
array[24603] <= 16'b0000_0000_0000_0000;
array[24604] <= 16'b0000_0000_0000_0000;
array[24605] <= 16'b0000_0000_0000_0000;
array[24606] <= 16'b0000_0000_0000_0000;
array[24607] <= 16'b0000_0000_0000_0000;
array[24608] <= 16'b0000_0000_0000_0000;
array[24609] <= 16'b0000_0000_0000_0000;
array[24610] <= 16'b0000_0000_0000_0000;
array[24611] <= 16'b0000_0000_0000_0000;
array[24612] <= 16'b0000_0000_0000_0000;
array[24613] <= 16'b0000_0000_0000_0000;
array[24614] <= 16'b0000_0000_0000_0000;
array[24615] <= 16'b0000_0000_0000_0000;
array[24616] <= 16'b0000_0000_0000_0000;
array[24617] <= 16'b0000_0000_0000_0000;
array[24618] <= 16'b0000_0000_0000_0000;
array[24619] <= 16'b0000_0000_0000_0000;
array[24620] <= 16'b0000_0000_0000_0000;
array[24621] <= 16'b0000_0000_0000_0000;
array[24622] <= 16'b0000_0000_0000_0000;
array[24623] <= 16'b0000_0000_0000_0000;
array[24624] <= 16'b0000_0000_0000_0000;
array[24625] <= 16'b0000_0000_0000_0000;
array[24626] <= 16'b0000_0000_0000_0000;
array[24627] <= 16'b0000_0000_0000_0000;
array[24628] <= 16'b0000_0000_0000_0000;
array[24629] <= 16'b0000_0000_0000_0000;
array[24630] <= 16'b0000_0000_0000_0000;
array[24631] <= 16'b0000_0000_0000_0000;
array[24632] <= 16'b0000_0000_0000_0000;
array[24633] <= 16'b0000_0000_0000_0000;
array[24634] <= 16'b0000_0000_0000_0000;
array[24635] <= 16'b0000_0000_0000_0000;
array[24636] <= 16'b0000_0000_0000_0000;
array[24637] <= 16'b0000_0000_0000_0000;
array[24638] <= 16'b0000_0000_0000_0000;
array[24639] <= 16'b0000_0000_0000_0000;
array[24640] <= 16'b0000_0000_0000_0000;
array[24641] <= 16'b0000_0000_0000_0000;
array[24642] <= 16'b0000_0000_0000_0000;
array[24643] <= 16'b0000_0000_0000_0000;
array[24644] <= 16'b0000_0000_0000_0000;
array[24645] <= 16'b0000_0000_0000_0000;
array[24646] <= 16'b0000_0000_0000_0000;
array[24647] <= 16'b0000_0000_0000_0000;
array[24648] <= 16'b0000_0000_0000_0000;
array[24649] <= 16'b0000_0000_0000_0000;
array[24650] <= 16'b0000_0000_0000_0000;
array[24651] <= 16'b0000_0000_0000_0000;
array[24652] <= 16'b0000_0000_0000_0000;
array[24653] <= 16'b0000_0000_0000_0000;
array[24654] <= 16'b0000_0000_0000_0000;
array[24655] <= 16'b0000_0000_0000_0000;
array[24656] <= 16'b0000_0000_0000_0000;
array[24657] <= 16'b0000_0000_0000_0000;
array[24658] <= 16'b0000_0000_0000_0000;
array[24659] <= 16'b0000_0000_0000_0000;
array[24660] <= 16'b0000_0000_0000_0000;
array[24661] <= 16'b0000_0000_0000_0000;
array[24662] <= 16'b0000_0000_0000_0000;
array[24663] <= 16'b0000_0000_0000_0000;
array[24664] <= 16'b0000_0000_0000_0000;
array[24665] <= 16'b0000_0000_0000_0000;
array[24666] <= 16'b0000_0000_0000_0000;
array[24667] <= 16'b0000_0000_0000_0000;
array[24668] <= 16'b0000_0000_0000_0000;
array[24669] <= 16'b0000_0000_0000_0000;
array[24670] <= 16'b0000_0000_0000_0000;
array[24671] <= 16'b0000_0000_0000_0000;
array[24672] <= 16'b0000_0000_0000_0000;
array[24673] <= 16'b0000_0000_0000_0000;
array[24674] <= 16'b0000_0000_0000_0000;
array[24675] <= 16'b0000_0000_0000_0000;
array[24676] <= 16'b0000_0000_0000_0000;
array[24677] <= 16'b0000_0000_0000_0000;
array[24678] <= 16'b0000_0000_0000_0000;
array[24679] <= 16'b0000_0000_0000_0000;
array[24680] <= 16'b0000_0000_0000_0000;
array[24681] <= 16'b0000_0000_0000_0000;
array[24682] <= 16'b0000_0000_0000_0000;
array[24683] <= 16'b0000_0000_0000_0000;
array[24684] <= 16'b0000_0000_0000_0000;
array[24685] <= 16'b0000_0000_0000_0000;
array[24686] <= 16'b0000_0000_0000_0000;
array[24687] <= 16'b0000_0000_0000_0000;
array[24688] <= 16'b0000_0000_0000_0000;
array[24689] <= 16'b0000_0000_0000_0000;
array[24690] <= 16'b0000_0000_0000_0000;
array[24691] <= 16'b0000_0000_0000_0000;
array[24692] <= 16'b0000_0000_0000_0000;
array[24693] <= 16'b0000_0000_0000_0000;
array[24694] <= 16'b0000_0000_0000_0000;
array[24695] <= 16'b0000_0000_0000_0000;
array[24696] <= 16'b0000_0000_0000_0000;
array[24697] <= 16'b0000_0000_0000_0000;
array[24698] <= 16'b0000_0000_0000_0000;
array[24699] <= 16'b0000_0000_0000_0000;
array[24700] <= 16'b0000_0000_0000_0000;
array[24701] <= 16'b0000_0000_0000_0000;
array[24702] <= 16'b0000_0000_0000_0000;
array[24703] <= 16'b0000_0000_0000_0000;
array[24704] <= 16'b0000_0000_0000_0000;
array[24705] <= 16'b0000_0000_0000_0000;
array[24706] <= 16'b0000_0000_0000_0000;
array[24707] <= 16'b0000_0000_0000_0000;
array[24708] <= 16'b0000_0000_0000_0000;
array[24709] <= 16'b0000_0000_0000_0000;
array[24710] <= 16'b0000_0000_0000_0000;
array[24711] <= 16'b0000_0000_0000_0000;
array[24712] <= 16'b0000_0000_0000_0000;
array[24713] <= 16'b0000_0000_0000_0000;
array[24714] <= 16'b0000_0000_0000_0000;
array[24715] <= 16'b0000_0000_0000_0000;
array[24716] <= 16'b0000_0000_0000_0000;
array[24717] <= 16'b0000_0000_0000_0000;
array[24718] <= 16'b0000_0000_0000_0000;
array[24719] <= 16'b0000_0000_0000_0000;
array[24720] <= 16'b0000_0000_0000_0000;
array[24721] <= 16'b0000_0000_0000_0000;
array[24722] <= 16'b0000_0000_0000_0000;
array[24723] <= 16'b0000_0000_0000_0000;
array[24724] <= 16'b0000_0000_0000_0000;
array[24725] <= 16'b0000_0000_0000_0000;
array[24726] <= 16'b0000_0000_0000_0000;
array[24727] <= 16'b0000_0000_0000_0000;
array[24728] <= 16'b0000_0000_0000_0000;
array[24729] <= 16'b0000_0000_0000_0000;
array[24730] <= 16'b0000_0000_0000_0000;
array[24731] <= 16'b0000_0000_0000_0000;
array[24732] <= 16'b0000_0000_0000_0000;
array[24733] <= 16'b0000_0000_0000_0000;
array[24734] <= 16'b0000_0000_0000_0000;
array[24735] <= 16'b0000_0000_0000_0000;
array[24736] <= 16'b0000_0000_0000_0000;
array[24737] <= 16'b0000_0000_0000_0000;
array[24738] <= 16'b0000_0000_0000_0000;
array[24739] <= 16'b0000_0000_0000_0000;
array[24740] <= 16'b0000_0000_0000_0000;
array[24741] <= 16'b0000_0000_0000_0000;
array[24742] <= 16'b0000_0000_0000_0000;
array[24743] <= 16'b0000_0000_0000_0000;
array[24744] <= 16'b0000_0000_0000_0000;
array[24745] <= 16'b0000_0000_0000_0000;
array[24746] <= 16'b0000_0000_0000_0000;
array[24747] <= 16'b0000_0000_0000_0000;
array[24748] <= 16'b0000_0000_0000_0000;
array[24749] <= 16'b0000_0000_0000_0000;
array[24750] <= 16'b0000_0000_0000_0000;
array[24751] <= 16'b0000_0000_0000_0000;
array[24752] <= 16'b0000_0000_0000_0000;
array[24753] <= 16'b0000_0000_0000_0000;
array[24754] <= 16'b0000_0000_0000_0000;
array[24755] <= 16'b0000_0000_0000_0000;
array[24756] <= 16'b0000_0000_0000_0000;
array[24757] <= 16'b0000_0000_0000_0000;
array[24758] <= 16'b0000_0000_0000_0000;
array[24759] <= 16'b0000_0000_0000_0000;
array[24760] <= 16'b0000_0000_0000_0000;
array[24761] <= 16'b0000_0000_0000_0000;
array[24762] <= 16'b0000_0000_0000_0000;
array[24763] <= 16'b0000_0000_0000_0000;
array[24764] <= 16'b0000_0000_0000_0000;
array[24765] <= 16'b0000_0000_0000_0000;
array[24766] <= 16'b0000_0000_0000_0000;
array[24767] <= 16'b0000_0000_0000_0000;
array[24768] <= 16'b0000_0000_0000_0000;
array[24769] <= 16'b0000_0000_0000_0000;
array[24770] <= 16'b0000_0000_0000_0000;
array[24771] <= 16'b0000_0000_0000_0000;
array[24772] <= 16'b0000_0000_0000_0000;
array[24773] <= 16'b0000_0000_0000_0000;
array[24774] <= 16'b0000_0000_0000_0000;
array[24775] <= 16'b0000_0000_0000_0000;
array[24776] <= 16'b0000_0000_0000_0000;
array[24777] <= 16'b0000_0000_0000_0000;
array[24778] <= 16'b0000_0000_0000_0000;
array[24779] <= 16'b0000_0000_0000_0000;
array[24780] <= 16'b0000_0000_0000_0000;
array[24781] <= 16'b0000_0000_0000_0000;
array[24782] <= 16'b0000_0000_0000_0000;
array[24783] <= 16'b0000_0000_0000_0000;
array[24784] <= 16'b0000_0000_0000_0000;
array[24785] <= 16'b0000_0000_0000_0000;
array[24786] <= 16'b0000_0000_0000_0000;
array[24787] <= 16'b0000_0000_0000_0000;
array[24788] <= 16'b0000_0000_0000_0000;
array[24789] <= 16'b0000_0000_0000_0000;
array[24790] <= 16'b0000_0000_0000_0000;
array[24791] <= 16'b0000_0000_0000_0000;
array[24792] <= 16'b0000_0000_0000_0000;
array[24793] <= 16'b0000_0000_0000_0000;
array[24794] <= 16'b0000_0000_0000_0000;
array[24795] <= 16'b0000_0000_0000_0000;
array[24796] <= 16'b0000_0000_0000_0000;
array[24797] <= 16'b0000_0000_0000_0000;
array[24798] <= 16'b0000_0000_0000_0000;
array[24799] <= 16'b0000_0000_0000_0000;
array[24800] <= 16'b0000_0000_0000_0000;
array[24801] <= 16'b0000_0000_0000_0000;
array[24802] <= 16'b0000_0000_0000_0000;
array[24803] <= 16'b0000_0000_0000_0000;
array[24804] <= 16'b0000_0000_0000_0000;
array[24805] <= 16'b0000_0000_0000_0000;
array[24806] <= 16'b0000_0000_0000_0000;
array[24807] <= 16'b0000_0000_0000_0000;
array[24808] <= 16'b0000_0000_0000_0000;
array[24809] <= 16'b0000_0000_0000_0000;
array[24810] <= 16'b0000_0000_0000_0000;
array[24811] <= 16'b0000_0000_0000_0000;
array[24812] <= 16'b0000_0000_0000_0000;
array[24813] <= 16'b0000_0000_0000_0000;
array[24814] <= 16'b0000_0000_0000_0000;
array[24815] <= 16'b0000_0000_0000_0000;
array[24816] <= 16'b0000_0000_0000_0000;
array[24817] <= 16'b0000_0000_0000_0000;
array[24818] <= 16'b0000_0000_0000_0000;
array[24819] <= 16'b0000_0000_0000_0000;
array[24820] <= 16'b0000_0000_0000_0000;
array[24821] <= 16'b0000_0000_0000_0000;
array[24822] <= 16'b0000_0000_0000_0000;
array[24823] <= 16'b0000_0000_0000_0000;
array[24824] <= 16'b0000_0000_0000_0000;
array[24825] <= 16'b0000_0000_0000_0000;
array[24826] <= 16'b0000_0000_0000_0000;
array[24827] <= 16'b0000_0000_0000_0000;
array[24828] <= 16'b0000_0000_0000_0000;
array[24829] <= 16'b0000_0000_0000_0000;
array[24830] <= 16'b0000_0000_0000_0000;
array[24831] <= 16'b0000_0000_0000_0000;
array[24832] <= 16'b0000_0000_0000_0000;
array[24833] <= 16'b0000_0000_0000_0000;
array[24834] <= 16'b0000_0000_0000_0000;
array[24835] <= 16'b0000_0000_0000_0000;
array[24836] <= 16'b0000_0000_0000_0000;
array[24837] <= 16'b0000_0000_0000_0000;
array[24838] <= 16'b0000_0000_0000_0000;
array[24839] <= 16'b0000_0000_0000_0000;
array[24840] <= 16'b0000_0000_0000_0000;
array[24841] <= 16'b0000_0000_0000_0000;
array[24842] <= 16'b0000_0000_0000_0000;
array[24843] <= 16'b0000_0000_0000_0000;
array[24844] <= 16'b0000_0000_0000_0000;
array[24845] <= 16'b0000_0000_0000_0000;
array[24846] <= 16'b0000_0000_0000_0000;
array[24847] <= 16'b0000_0000_0000_0000;
array[24848] <= 16'b0000_0000_0000_0000;
array[24849] <= 16'b0000_0000_0000_0000;
array[24850] <= 16'b0000_0000_0000_0000;
array[24851] <= 16'b0000_0000_0000_0000;
array[24852] <= 16'b0000_0000_0000_0000;
array[24853] <= 16'b0000_0000_0000_0000;
array[24854] <= 16'b0000_0000_0000_0000;
array[24855] <= 16'b0000_0000_0000_0000;
array[24856] <= 16'b0000_0000_0000_0000;
array[24857] <= 16'b0000_0000_0000_0000;
array[24858] <= 16'b0000_0000_0000_0000;
array[24859] <= 16'b0000_0000_0000_0000;
array[24860] <= 16'b0000_0000_0000_0000;
array[24861] <= 16'b0000_0000_0000_0000;
array[24862] <= 16'b0000_0000_0000_0000;
array[24863] <= 16'b0000_0000_0000_0000;
array[24864] <= 16'b0000_0000_0000_0000;
array[24865] <= 16'b0000_0000_0000_0000;
array[24866] <= 16'b0000_0000_0000_0000;
array[24867] <= 16'b0000_0000_0000_0000;
array[24868] <= 16'b0000_0000_0000_0000;
array[24869] <= 16'b0000_0000_0000_0000;
array[24870] <= 16'b0000_0000_0000_0000;
array[24871] <= 16'b0000_0000_0000_0000;
array[24872] <= 16'b0000_0000_0000_0000;
array[24873] <= 16'b0000_0000_0000_0000;
array[24874] <= 16'b0000_0000_0000_0000;
array[24875] <= 16'b0000_0000_0000_0000;
array[24876] <= 16'b0000_0000_0000_0000;
array[24877] <= 16'b0000_0000_0000_0000;
array[24878] <= 16'b0000_0000_0000_0000;
array[24879] <= 16'b0000_0000_0000_0000;
array[24880] <= 16'b0000_0000_0000_0000;
array[24881] <= 16'b0000_0000_0000_0000;
array[24882] <= 16'b0000_0000_0000_0000;
array[24883] <= 16'b0000_0000_0000_0000;
array[24884] <= 16'b0000_0000_0000_0000;
array[24885] <= 16'b0000_0000_0000_0000;
array[24886] <= 16'b0000_0000_0000_0000;
array[24887] <= 16'b0000_0000_0000_0000;
array[24888] <= 16'b0000_0000_0000_0000;
array[24889] <= 16'b0000_0000_0000_0000;
array[24890] <= 16'b0000_0000_0000_0000;
array[24891] <= 16'b0000_0000_0000_0000;
array[24892] <= 16'b0000_0000_0000_0000;
array[24893] <= 16'b0000_0000_0000_0000;
array[24894] <= 16'b0000_0000_0000_0000;
array[24895] <= 16'b0000_0000_0000_0000;
array[24896] <= 16'b0000_0000_0000_0000;
array[24897] <= 16'b0000_0000_0000_0000;
array[24898] <= 16'b0000_0000_0000_0000;
array[24899] <= 16'b0000_0000_0000_0000;
array[24900] <= 16'b0000_0000_0000_0000;
array[24901] <= 16'b0000_0000_0000_0000;
array[24902] <= 16'b0000_0000_0000_0000;
array[24903] <= 16'b0000_0000_0000_0000;
array[24904] <= 16'b0000_0000_0000_0000;
array[24905] <= 16'b0000_0000_0000_0000;
array[24906] <= 16'b0000_0000_0000_0000;
array[24907] <= 16'b0000_0000_0000_0000;
array[24908] <= 16'b0000_0000_0000_0000;
array[24909] <= 16'b0000_0000_0000_0000;
array[24910] <= 16'b0000_0000_0000_0000;
array[24911] <= 16'b0000_0000_0000_0000;
array[24912] <= 16'b0000_0000_0000_0000;
array[24913] <= 16'b0000_0000_0000_0000;
array[24914] <= 16'b0000_0000_0000_0000;
array[24915] <= 16'b0000_0000_0000_0000;
array[24916] <= 16'b0000_0000_0000_0000;
array[24917] <= 16'b0000_0000_0000_0000;
array[24918] <= 16'b0000_0000_0000_0000;
array[24919] <= 16'b0000_0000_0000_0000;
array[24920] <= 16'b0000_0000_0000_0000;
array[24921] <= 16'b0000_0000_0000_0000;
array[24922] <= 16'b0000_0000_0000_0000;
array[24923] <= 16'b0000_0000_0000_0000;
array[24924] <= 16'b0000_0000_0000_0000;
array[24925] <= 16'b0000_0000_0000_0000;
array[24926] <= 16'b0000_0000_0000_0000;
array[24927] <= 16'b0000_0000_0000_0000;
array[24928] <= 16'b0000_0000_0000_0000;
array[24929] <= 16'b0000_0000_0000_0000;
array[24930] <= 16'b0000_0000_0000_0000;
array[24931] <= 16'b0000_0000_0000_0000;
array[24932] <= 16'b0000_0000_0000_0000;
array[24933] <= 16'b0000_0000_0000_0000;
array[24934] <= 16'b0000_0000_0000_0000;
array[24935] <= 16'b0000_0000_0000_0000;
array[24936] <= 16'b0000_0000_0000_0000;
array[24937] <= 16'b0000_0000_0000_0000;
array[24938] <= 16'b0000_0000_0000_0000;
array[24939] <= 16'b0000_0000_0000_0000;
array[24940] <= 16'b0000_0000_0000_0000;
array[24941] <= 16'b0000_0000_0000_0000;
array[24942] <= 16'b0000_0000_0000_0000;
array[24943] <= 16'b0000_0000_0000_0000;
array[24944] <= 16'b0000_0000_0000_0000;
array[24945] <= 16'b0000_0000_0000_0000;
array[24946] <= 16'b0000_0000_0000_0000;
array[24947] <= 16'b0000_0000_0000_0000;
array[24948] <= 16'b0000_0000_0000_0000;
array[24949] <= 16'b0000_0000_0000_0000;
array[24950] <= 16'b0000_0000_0000_0000;
array[24951] <= 16'b0000_0000_0000_0000;
array[24952] <= 16'b0000_0000_0000_0000;
array[24953] <= 16'b0000_0000_0000_0000;
array[24954] <= 16'b0000_0000_0000_0000;
array[24955] <= 16'b0000_0000_0000_0000;
array[24956] <= 16'b0000_0000_0000_0000;
array[24957] <= 16'b0000_0000_0000_0000;
array[24958] <= 16'b0000_0000_0000_0000;
array[24959] <= 16'b0000_0000_0000_0000;
array[24960] <= 16'b0000_0000_0000_0000;
array[24961] <= 16'b0000_0000_0000_0000;
array[24962] <= 16'b0000_0000_0000_0000;
array[24963] <= 16'b0000_0000_0000_0000;
array[24964] <= 16'b0000_0000_0000_0000;
array[24965] <= 16'b0000_0000_0000_0000;
array[24966] <= 16'b0000_0000_0000_0000;
array[24967] <= 16'b0000_0000_0000_0000;
array[24968] <= 16'b0000_0000_0000_0000;
array[24969] <= 16'b0000_0000_0000_0000;
array[24970] <= 16'b0000_0000_0000_0000;
array[24971] <= 16'b0000_0000_0000_0000;
array[24972] <= 16'b0000_0000_0000_0000;
array[24973] <= 16'b0000_0000_0000_0000;
array[24974] <= 16'b0000_0000_0000_0000;
array[24975] <= 16'b0000_0000_0000_0000;
array[24976] <= 16'b0000_0000_0000_0000;
array[24977] <= 16'b0000_0000_0000_0000;
array[24978] <= 16'b0000_0000_0000_0000;
array[24979] <= 16'b0000_0000_0000_0000;
array[24980] <= 16'b0000_0000_0000_0000;
array[24981] <= 16'b0000_0000_0000_0000;
array[24982] <= 16'b0000_0000_0000_0000;
array[24983] <= 16'b0000_0000_0000_0000;
array[24984] <= 16'b0000_0000_0000_0000;
array[24985] <= 16'b0000_0000_0000_0000;
array[24986] <= 16'b0000_0000_0000_0000;
array[24987] <= 16'b0000_0000_0000_0000;
array[24988] <= 16'b0000_0000_0000_0000;
array[24989] <= 16'b0000_0000_0000_0000;
array[24990] <= 16'b0000_0000_0000_0000;
array[24991] <= 16'b0000_0000_0000_0000;
array[24992] <= 16'b0000_0000_0000_0000;
array[24993] <= 16'b0000_0000_0000_0000;
array[24994] <= 16'b0000_0000_0000_0000;
array[24995] <= 16'b0000_0000_0000_0000;
array[24996] <= 16'b0000_0000_0000_0000;
array[24997] <= 16'b0000_0000_0000_0000;
array[24998] <= 16'b0000_0000_0000_0000;
array[24999] <= 16'b0000_0000_0000_0000;
array[25000] <= 16'b0000_0000_0000_0000;
array[25001] <= 16'b0000_0000_0000_0000;
array[25002] <= 16'b0000_0000_0000_0000;
array[25003] <= 16'b0000_0000_0000_0000;
array[25004] <= 16'b0000_0000_0000_0000;
array[25005] <= 16'b0000_0000_0000_0000;
array[25006] <= 16'b0000_0000_0000_0000;
array[25007] <= 16'b0000_0000_0000_0000;
array[25008] <= 16'b0000_0000_0000_0000;
array[25009] <= 16'b0000_0000_0000_0000;
array[25010] <= 16'b0000_0000_0000_0000;
array[25011] <= 16'b0000_0000_0000_0000;
array[25012] <= 16'b0000_0000_0000_0000;
array[25013] <= 16'b0000_0000_0000_0000;
array[25014] <= 16'b0000_0000_0000_0000;
array[25015] <= 16'b0000_0000_0000_0000;
array[25016] <= 16'b0000_0000_0000_0000;
array[25017] <= 16'b0000_0000_0000_0000;
array[25018] <= 16'b0000_0000_0000_0000;
array[25019] <= 16'b0000_0000_0000_0000;
array[25020] <= 16'b0000_0000_0000_0000;
array[25021] <= 16'b0000_0000_0000_0000;
array[25022] <= 16'b0000_0000_0000_0000;
array[25023] <= 16'b0000_0000_0000_0000;
array[25024] <= 16'b0000_0000_0000_0000;
array[25025] <= 16'b0000_0000_0000_0000;
array[25026] <= 16'b0000_0000_0000_0000;
array[25027] <= 16'b0000_0000_0000_0000;
array[25028] <= 16'b0000_0000_0000_0000;
array[25029] <= 16'b0000_0000_0000_0000;
array[25030] <= 16'b0000_0000_0000_0000;
array[25031] <= 16'b0000_0000_0000_0000;
array[25032] <= 16'b0000_0000_0000_0000;
array[25033] <= 16'b0000_0000_0000_0000;
array[25034] <= 16'b0000_0000_0000_0000;
array[25035] <= 16'b0000_0000_0000_0000;
array[25036] <= 16'b0000_0000_0000_0000;
array[25037] <= 16'b0000_0000_0000_0000;
array[25038] <= 16'b0000_0000_0000_0000;
array[25039] <= 16'b0000_0000_0000_0000;
array[25040] <= 16'b0000_0000_0000_0000;
array[25041] <= 16'b0000_0000_0000_0000;
array[25042] <= 16'b0000_0000_0000_0000;
array[25043] <= 16'b0000_0000_0000_0000;
array[25044] <= 16'b0000_0000_0000_0000;
array[25045] <= 16'b0000_0000_0000_0000;
array[25046] <= 16'b0000_0000_0000_0000;
array[25047] <= 16'b0000_0000_0000_0000;
array[25048] <= 16'b0000_0000_0000_0000;
array[25049] <= 16'b0000_0000_0000_0000;
array[25050] <= 16'b0000_0000_0000_0000;
array[25051] <= 16'b0000_0000_0000_0000;
array[25052] <= 16'b0000_0000_0000_0000;
array[25053] <= 16'b0000_0000_0000_0000;
array[25054] <= 16'b0000_0000_0000_0000;
array[25055] <= 16'b0000_0000_0000_0000;
array[25056] <= 16'b0000_0000_0000_0000;
array[25057] <= 16'b0000_0000_0000_0000;
array[25058] <= 16'b0000_0000_0000_0000;
array[25059] <= 16'b0000_0000_0000_0000;
array[25060] <= 16'b0000_0000_0000_0000;
array[25061] <= 16'b0000_0000_0000_0000;
array[25062] <= 16'b0000_0000_0000_0000;
array[25063] <= 16'b0000_0000_0000_0000;
array[25064] <= 16'b0000_0000_0000_0000;
array[25065] <= 16'b0000_0000_0000_0000;
array[25066] <= 16'b0000_0000_0000_0000;
array[25067] <= 16'b0000_0000_0000_0000;
array[25068] <= 16'b0000_0000_0000_0000;
array[25069] <= 16'b0000_0000_0000_0000;
array[25070] <= 16'b0000_0000_0000_0000;
array[25071] <= 16'b0000_0000_0000_0000;
array[25072] <= 16'b0000_0000_0000_0000;
array[25073] <= 16'b0000_0000_0000_0000;
array[25074] <= 16'b0000_0000_0000_0000;
array[25075] <= 16'b0000_0000_0000_0000;
array[25076] <= 16'b0000_0000_0000_0000;
array[25077] <= 16'b0000_0000_0000_0000;
array[25078] <= 16'b0000_0000_0000_0000;
array[25079] <= 16'b0000_0000_0000_0000;
array[25080] <= 16'b0000_0000_0000_0000;
array[25081] <= 16'b0000_0000_0000_0000;
array[25082] <= 16'b0000_0000_0000_0000;
array[25083] <= 16'b0000_0000_0000_0000;
array[25084] <= 16'b0000_0000_0000_0000;
array[25085] <= 16'b0000_0000_0000_0000;
array[25086] <= 16'b0000_0000_0000_0000;
array[25087] <= 16'b0000_0000_0000_0000;
array[25088] <= 16'b0000_0000_0000_0000;
array[25089] <= 16'b0000_0000_0000_0000;
array[25090] <= 16'b0000_0000_0000_0000;
array[25091] <= 16'b0000_0000_0000_0000;
array[25092] <= 16'b0000_0000_0000_0000;
array[25093] <= 16'b0000_0000_0000_0000;
array[25094] <= 16'b0000_0000_0000_0000;
array[25095] <= 16'b0000_0000_0000_0000;
array[25096] <= 16'b0000_0000_0000_0000;
array[25097] <= 16'b0000_0000_0000_0000;
array[25098] <= 16'b0000_0000_0000_0000;
array[25099] <= 16'b0000_0000_0000_0000;
array[25100] <= 16'b0000_0000_0000_0000;
array[25101] <= 16'b0000_0000_0000_0000;
array[25102] <= 16'b0000_0000_0000_0000;
array[25103] <= 16'b0000_0000_0000_0000;
array[25104] <= 16'b0000_0000_0000_0000;
array[25105] <= 16'b0000_0000_0000_0000;
array[25106] <= 16'b0000_0000_0000_0000;
array[25107] <= 16'b0000_0000_0000_0000;
array[25108] <= 16'b0000_0000_0000_0000;
array[25109] <= 16'b0000_0000_0000_0000;
array[25110] <= 16'b0000_0000_0000_0000;
array[25111] <= 16'b0000_0000_0000_0000;
array[25112] <= 16'b0000_0000_0000_0000;
array[25113] <= 16'b0000_0000_0000_0000;
array[25114] <= 16'b0000_0000_0000_0000;
array[25115] <= 16'b0000_0000_0000_0000;
array[25116] <= 16'b0000_0000_0000_0000;
array[25117] <= 16'b0000_0000_0000_0000;
array[25118] <= 16'b0000_0000_0000_0000;
array[25119] <= 16'b0000_0000_0000_0000;
array[25120] <= 16'b0000_0000_0000_0000;
array[25121] <= 16'b0000_0000_0000_0000;
array[25122] <= 16'b0000_0000_0000_0000;
array[25123] <= 16'b0000_0000_0000_0000;
array[25124] <= 16'b0000_0000_0000_0000;
array[25125] <= 16'b0000_0000_0000_0000;
array[25126] <= 16'b0000_0000_0000_0000;
array[25127] <= 16'b0000_0000_0000_0000;
array[25128] <= 16'b0000_0000_0000_0000;
array[25129] <= 16'b0000_0000_0000_0000;
array[25130] <= 16'b0000_0000_0000_0000;
array[25131] <= 16'b0000_0000_0000_0000;
array[25132] <= 16'b0000_0000_0000_0000;
array[25133] <= 16'b0000_0000_0000_0000;
array[25134] <= 16'b0000_0000_0000_0000;
array[25135] <= 16'b0000_0000_0000_0000;
array[25136] <= 16'b0000_0000_0000_0000;
array[25137] <= 16'b0000_0000_0000_0000;
array[25138] <= 16'b0000_0000_0000_0000;
array[25139] <= 16'b0000_0000_0000_0000;
array[25140] <= 16'b0000_0000_0000_0000;
array[25141] <= 16'b0000_0000_0000_0000;
array[25142] <= 16'b0000_0000_0000_0000;
array[25143] <= 16'b0000_0000_0000_0000;
array[25144] <= 16'b0000_0000_0000_0000;
array[25145] <= 16'b0000_0000_0000_0000;
array[25146] <= 16'b0000_0000_0000_0000;
array[25147] <= 16'b0000_0000_0000_0000;
array[25148] <= 16'b0000_0000_0000_0000;
array[25149] <= 16'b0000_0000_0000_0000;
array[25150] <= 16'b0000_0000_0000_0000;
array[25151] <= 16'b0000_0000_0000_0000;
array[25152] <= 16'b0000_0000_0000_0000;
array[25153] <= 16'b0000_0000_0000_0000;
array[25154] <= 16'b0000_0000_0000_0000;
array[25155] <= 16'b0000_0000_0000_0000;
array[25156] <= 16'b0000_0000_0000_0000;
array[25157] <= 16'b0000_0000_0000_0000;
array[25158] <= 16'b0000_0000_0000_0000;
array[25159] <= 16'b0000_0000_0000_0000;
array[25160] <= 16'b0000_0000_0000_0000;
array[25161] <= 16'b0000_0000_0000_0000;
array[25162] <= 16'b0000_0000_0000_0000;
array[25163] <= 16'b0000_0000_0000_0000;
array[25164] <= 16'b0000_0000_0000_0000;
array[25165] <= 16'b0000_0000_0000_0000;
array[25166] <= 16'b0000_0000_0000_0000;
array[25167] <= 16'b0000_0000_0000_0000;
array[25168] <= 16'b0000_0000_0000_0000;
array[25169] <= 16'b0000_0000_0000_0000;
array[25170] <= 16'b0000_0000_0000_0000;
array[25171] <= 16'b0000_0000_0000_0000;
array[25172] <= 16'b0000_0000_0000_0000;
array[25173] <= 16'b0000_0000_0000_0000;
array[25174] <= 16'b0000_0000_0000_0000;
array[25175] <= 16'b0000_0000_0000_0000;
array[25176] <= 16'b0000_0000_0000_0000;
array[25177] <= 16'b0000_0000_0000_0000;
array[25178] <= 16'b0000_0000_0000_0000;
array[25179] <= 16'b0000_0000_0000_0000;
array[25180] <= 16'b0000_0000_0000_0000;
array[25181] <= 16'b0000_0000_0000_0000;
array[25182] <= 16'b0000_0000_0000_0000;
array[25183] <= 16'b0000_0000_0000_0000;
array[25184] <= 16'b0000_0000_0000_0000;
array[25185] <= 16'b0000_0000_0000_0000;
array[25186] <= 16'b0000_0000_0000_0000;
array[25187] <= 16'b0000_0000_0000_0000;
array[25188] <= 16'b0000_0000_0000_0000;
array[25189] <= 16'b0000_0000_0000_0000;
array[25190] <= 16'b0000_0000_0000_0000;
array[25191] <= 16'b0000_0000_0000_0000;
array[25192] <= 16'b0000_0000_0000_0000;
array[25193] <= 16'b0000_0000_0000_0000;
array[25194] <= 16'b0000_0000_0000_0000;
array[25195] <= 16'b0000_0000_0000_0000;
array[25196] <= 16'b0000_0000_0000_0000;
array[25197] <= 16'b0000_0000_0000_0000;
array[25198] <= 16'b0000_0000_0000_0000;
array[25199] <= 16'b0000_0000_0000_0000;
array[25200] <= 16'b0000_0000_0000_0000;
array[25201] <= 16'b0000_0000_0000_0000;
array[25202] <= 16'b0000_0000_0000_0000;
array[25203] <= 16'b0000_0000_0000_0000;
array[25204] <= 16'b0000_0000_0000_0000;
array[25205] <= 16'b0000_0000_0000_0000;
array[25206] <= 16'b0000_0000_0000_0000;
array[25207] <= 16'b0000_0000_0000_0000;
array[25208] <= 16'b0000_0000_0000_0000;
array[25209] <= 16'b0000_0000_0000_0000;
array[25210] <= 16'b0000_0000_0000_0000;
array[25211] <= 16'b0000_0000_0000_0000;
array[25212] <= 16'b0000_0000_0000_0000;
array[25213] <= 16'b0000_0000_0000_0000;
array[25214] <= 16'b0000_0000_0000_0000;
array[25215] <= 16'b0000_0000_0000_0000;
array[25216] <= 16'b0000_0000_0000_0000;
array[25217] <= 16'b0000_0000_0000_0000;
array[25218] <= 16'b0000_0000_0000_0000;
array[25219] <= 16'b0000_0000_0000_0000;
array[25220] <= 16'b0000_0000_0000_0000;
array[25221] <= 16'b0000_0000_0000_0000;
array[25222] <= 16'b0000_0000_0000_0000;
array[25223] <= 16'b0000_0000_0000_0000;
array[25224] <= 16'b0000_0000_0000_0000;
array[25225] <= 16'b0000_0000_0000_0000;
array[25226] <= 16'b0000_0000_0000_0000;
array[25227] <= 16'b0000_0000_0000_0000;
array[25228] <= 16'b0000_0000_0000_0000;
array[25229] <= 16'b0000_0000_0000_0000;
array[25230] <= 16'b0000_0000_0000_0000;
array[25231] <= 16'b0000_0000_0000_0000;
array[25232] <= 16'b0000_0000_0000_0000;
array[25233] <= 16'b0000_0000_0000_0000;
array[25234] <= 16'b0000_0000_0000_0000;
array[25235] <= 16'b0000_0000_0000_0000;
array[25236] <= 16'b0000_0000_0000_0000;
array[25237] <= 16'b0000_0000_0000_0000;
array[25238] <= 16'b0000_0000_0000_0000;
array[25239] <= 16'b0000_0000_0000_0000;
array[25240] <= 16'b0000_0000_0000_0000;
array[25241] <= 16'b0000_0000_0000_0000;
array[25242] <= 16'b0000_0000_0000_0000;
array[25243] <= 16'b0000_0000_0000_0000;
array[25244] <= 16'b0000_0000_0000_0000;
array[25245] <= 16'b0000_0000_0000_0000;
array[25246] <= 16'b0000_0000_0000_0000;
array[25247] <= 16'b0000_0000_0000_0000;
array[25248] <= 16'b0000_0000_0000_0000;
array[25249] <= 16'b0000_0000_0000_0000;
array[25250] <= 16'b0000_0000_0000_0000;
array[25251] <= 16'b0000_0000_0000_0000;
array[25252] <= 16'b0000_0000_0000_0000;
array[25253] <= 16'b0000_0000_0000_0000;
array[25254] <= 16'b0000_0000_0000_0000;
array[25255] <= 16'b0000_0000_0000_0000;
array[25256] <= 16'b0000_0000_0000_0000;
array[25257] <= 16'b0000_0000_0000_0000;
array[25258] <= 16'b0000_0000_0000_0000;
array[25259] <= 16'b0000_0000_0000_0000;
array[25260] <= 16'b0000_0000_0000_0000;
array[25261] <= 16'b0000_0000_0000_0000;
array[25262] <= 16'b0000_0000_0000_0000;
array[25263] <= 16'b0000_0000_0000_0000;
array[25264] <= 16'b0000_0000_0000_0000;
array[25265] <= 16'b0000_0000_0000_0000;
array[25266] <= 16'b0000_0000_0000_0000;
array[25267] <= 16'b0000_0000_0000_0000;
array[25268] <= 16'b0000_0000_0000_0000;
array[25269] <= 16'b0000_0000_0000_0000;
array[25270] <= 16'b0000_0000_0000_0000;
array[25271] <= 16'b0000_0000_0000_0000;
array[25272] <= 16'b0000_0000_0000_0000;
array[25273] <= 16'b0000_0000_0000_0000;
array[25274] <= 16'b0000_0000_0000_0000;
array[25275] <= 16'b0000_0000_0000_0000;
array[25276] <= 16'b0000_0000_0000_0000;
array[25277] <= 16'b0000_0000_0000_0000;
array[25278] <= 16'b0000_0000_0000_0000;
array[25279] <= 16'b0000_0000_0000_0000;
array[25280] <= 16'b0000_0000_0000_0000;
array[25281] <= 16'b0000_0000_0000_0000;
array[25282] <= 16'b0000_0000_0000_0000;
array[25283] <= 16'b0000_0000_0000_0000;
array[25284] <= 16'b0000_0000_0000_0000;
array[25285] <= 16'b0000_0000_0000_0000;
array[25286] <= 16'b0000_0000_0000_0000;
array[25287] <= 16'b0000_0000_0000_0000;
array[25288] <= 16'b0000_0000_0000_0000;
array[25289] <= 16'b0000_0000_0000_0000;
array[25290] <= 16'b0000_0000_0000_0000;
array[25291] <= 16'b0000_0000_0000_0000;
array[25292] <= 16'b0000_0000_0000_0000;
array[25293] <= 16'b0000_0000_0000_0000;
array[25294] <= 16'b0000_0000_0000_0000;
array[25295] <= 16'b0000_0000_0000_0000;
array[25296] <= 16'b0000_0000_0000_0000;
array[25297] <= 16'b0000_0000_0000_0000;
array[25298] <= 16'b0000_0000_0000_0000;
array[25299] <= 16'b0000_0000_0000_0000;
array[25300] <= 16'b0000_0000_0000_0000;
array[25301] <= 16'b0000_0000_0000_0000;
array[25302] <= 16'b0000_0000_0000_0000;
array[25303] <= 16'b0000_0000_0000_0000;
array[25304] <= 16'b0000_0000_0000_0000;
array[25305] <= 16'b0000_0000_0000_0000;
array[25306] <= 16'b0000_0000_0000_0000;
array[25307] <= 16'b0000_0000_0000_0000;
array[25308] <= 16'b0000_0000_0000_0000;
array[25309] <= 16'b0000_0000_0000_0000;
array[25310] <= 16'b0000_0000_0000_0000;
array[25311] <= 16'b0000_0000_0000_0000;
array[25312] <= 16'b0000_0000_0000_0000;
array[25313] <= 16'b0000_0000_0000_0000;
array[25314] <= 16'b0000_0000_0000_0000;
array[25315] <= 16'b0000_0000_0000_0000;
array[25316] <= 16'b0000_0000_0000_0000;
array[25317] <= 16'b0000_0000_0000_0000;
array[25318] <= 16'b0000_0000_0000_0000;
array[25319] <= 16'b0000_0000_0000_0000;
array[25320] <= 16'b0000_0000_0000_0000;
array[25321] <= 16'b0000_0000_0000_0000;
array[25322] <= 16'b0000_0000_0000_0000;
array[25323] <= 16'b0000_0000_0000_0000;
array[25324] <= 16'b0000_0000_0000_0000;
array[25325] <= 16'b0000_0000_0000_0000;
array[25326] <= 16'b0000_0000_0000_0000;
array[25327] <= 16'b0000_0000_0000_0000;
array[25328] <= 16'b0000_0000_0000_0000;
array[25329] <= 16'b0000_0000_0000_0000;
array[25330] <= 16'b0000_0000_0000_0000;
array[25331] <= 16'b0000_0000_0000_0000;
array[25332] <= 16'b0000_0000_0000_0000;
array[25333] <= 16'b0000_0000_0000_0000;
array[25334] <= 16'b0000_0000_0000_0000;
array[25335] <= 16'b0000_0000_0000_0000;
array[25336] <= 16'b0000_0000_0000_0000;
array[25337] <= 16'b0000_0000_0000_0000;
array[25338] <= 16'b0000_0000_0000_0000;
array[25339] <= 16'b0000_0000_0000_0000;
array[25340] <= 16'b0000_0000_0000_0000;
array[25341] <= 16'b0000_0000_0000_0000;
array[25342] <= 16'b0000_0000_0000_0000;
array[25343] <= 16'b0000_0000_0000_0000;
array[25344] <= 16'b0000_0000_0000_0000;
array[25345] <= 16'b0000_0000_0000_0000;
array[25346] <= 16'b0000_0000_0000_0000;
array[25347] <= 16'b0000_0000_0000_0000;
array[25348] <= 16'b0000_0000_0000_0000;
array[25349] <= 16'b0000_0000_0000_0000;
array[25350] <= 16'b0000_0000_0000_0000;
array[25351] <= 16'b0000_0000_0000_0000;
array[25352] <= 16'b0000_0000_0000_0000;
array[25353] <= 16'b0000_0000_0000_0000;
array[25354] <= 16'b0000_0000_0000_0000;
array[25355] <= 16'b0000_0000_0000_0000;
array[25356] <= 16'b0000_0000_0000_0000;
array[25357] <= 16'b0000_0000_0000_0000;
array[25358] <= 16'b0000_0000_0000_0000;
array[25359] <= 16'b0000_0000_0000_0000;
array[25360] <= 16'b0000_0000_0000_0000;
array[25361] <= 16'b0000_0000_0000_0000;
array[25362] <= 16'b0000_0000_0000_0000;
array[25363] <= 16'b0000_0000_0000_0000;
array[25364] <= 16'b0000_0000_0000_0000;
array[25365] <= 16'b0000_0000_0000_0000;
array[25366] <= 16'b0000_0000_0000_0000;
array[25367] <= 16'b0000_0000_0000_0000;
array[25368] <= 16'b0000_0000_0000_0000;
array[25369] <= 16'b0000_0000_0000_0000;
array[25370] <= 16'b0000_0000_0000_0000;
array[25371] <= 16'b0000_0000_0000_0000;
array[25372] <= 16'b0000_0000_0000_0000;
array[25373] <= 16'b0000_0000_0000_0000;
array[25374] <= 16'b0000_0000_0000_0000;
array[25375] <= 16'b0000_0000_0000_0000;
array[25376] <= 16'b0000_0000_0000_0000;
array[25377] <= 16'b0000_0000_0000_0000;
array[25378] <= 16'b0000_0000_0000_0000;
array[25379] <= 16'b0000_0000_0000_0000;
array[25380] <= 16'b0000_0000_0000_0000;
array[25381] <= 16'b0000_0000_0000_0000;
array[25382] <= 16'b0000_0000_0000_0000;
array[25383] <= 16'b0000_0000_0000_0000;
array[25384] <= 16'b0000_0000_0000_0000;
array[25385] <= 16'b0000_0000_0000_0000;
array[25386] <= 16'b0000_0000_0000_0000;
array[25387] <= 16'b0000_0000_0000_0000;
array[25388] <= 16'b0000_0000_0000_0000;
array[25389] <= 16'b0000_0000_0000_0000;
array[25390] <= 16'b0000_0000_0000_0000;
array[25391] <= 16'b0000_0000_0000_0000;
array[25392] <= 16'b0000_0000_0000_0000;
array[25393] <= 16'b0000_0000_0000_0000;
array[25394] <= 16'b0000_0000_0000_0000;
array[25395] <= 16'b0000_0000_0000_0000;
array[25396] <= 16'b0000_0000_0000_0000;
array[25397] <= 16'b0000_0000_0000_0000;
array[25398] <= 16'b0000_0000_0000_0000;
array[25399] <= 16'b0000_0000_0000_0000;
array[25400] <= 16'b0000_0000_0000_0000;
array[25401] <= 16'b0000_0000_0000_0000;
array[25402] <= 16'b0000_0000_0000_0000;
array[25403] <= 16'b0000_0000_0000_0000;
array[25404] <= 16'b0000_0000_0000_0000;
array[25405] <= 16'b0000_0000_0000_0000;
array[25406] <= 16'b0000_0000_0000_0000;
array[25407] <= 16'b0000_0000_0000_0000;
array[25408] <= 16'b0000_0000_0000_0000;
array[25409] <= 16'b0000_0000_0000_0000;
array[25410] <= 16'b0000_0000_0000_0000;
array[25411] <= 16'b0000_0000_0000_0000;
array[25412] <= 16'b0000_0000_0000_0000;
array[25413] <= 16'b0000_0000_0000_0000;
array[25414] <= 16'b0000_0000_0000_0000;
array[25415] <= 16'b0000_0000_0000_0000;
array[25416] <= 16'b0000_0000_0000_0000;
array[25417] <= 16'b0000_0000_0000_0000;
array[25418] <= 16'b0000_0000_0000_0000;
array[25419] <= 16'b0000_0000_0000_0000;
array[25420] <= 16'b0000_0000_0000_0000;
array[25421] <= 16'b0000_0000_0000_0000;
array[25422] <= 16'b0000_0000_0000_0000;
array[25423] <= 16'b0000_0000_0000_0000;
array[25424] <= 16'b0000_0000_0000_0000;
array[25425] <= 16'b0000_0000_0000_0000;
array[25426] <= 16'b0000_0000_0000_0000;
array[25427] <= 16'b0000_0000_0000_0000;
array[25428] <= 16'b0000_0000_0000_0000;
array[25429] <= 16'b0000_0000_0000_0000;
array[25430] <= 16'b0000_0000_0000_0000;
array[25431] <= 16'b0000_0000_0000_0000;
array[25432] <= 16'b0000_0000_0000_0000;
array[25433] <= 16'b0000_0000_0000_0000;
array[25434] <= 16'b0000_0000_0000_0000;
array[25435] <= 16'b0000_0000_0000_0000;
array[25436] <= 16'b0000_0000_0000_0000;
array[25437] <= 16'b0000_0000_0000_0000;
array[25438] <= 16'b0000_0000_0000_0000;
array[25439] <= 16'b0000_0000_0000_0000;
array[25440] <= 16'b0000_0000_0000_0000;
array[25441] <= 16'b0000_0000_0000_0000;
array[25442] <= 16'b0000_0000_0000_0000;
array[25443] <= 16'b0000_0000_0000_0000;
array[25444] <= 16'b0000_0000_0000_0000;
array[25445] <= 16'b0000_0000_0000_0000;
array[25446] <= 16'b0000_0000_0000_0000;
array[25447] <= 16'b0000_0000_0000_0000;
array[25448] <= 16'b0000_0000_0000_0000;
array[25449] <= 16'b0000_0000_0000_0000;
array[25450] <= 16'b0000_0000_0000_0000;
array[25451] <= 16'b0000_0000_0000_0000;
array[25452] <= 16'b0000_0000_0000_0000;
array[25453] <= 16'b0000_0000_0000_0000;
array[25454] <= 16'b0000_0000_0000_0000;
array[25455] <= 16'b0000_0000_0000_0000;
array[25456] <= 16'b0000_0000_0000_0000;
array[25457] <= 16'b0000_0000_0000_0000;
array[25458] <= 16'b0000_0000_0000_0000;
array[25459] <= 16'b0000_0000_0000_0000;
array[25460] <= 16'b0000_0000_0000_0000;
array[25461] <= 16'b0000_0000_0000_0000;
array[25462] <= 16'b0000_0000_0000_0000;
array[25463] <= 16'b0000_0000_0000_0000;
array[25464] <= 16'b0000_0000_0000_0000;
array[25465] <= 16'b0000_0000_0000_0000;
array[25466] <= 16'b0000_0000_0000_0000;
array[25467] <= 16'b0000_0000_0000_0000;
array[25468] <= 16'b0000_0000_0000_0000;
array[25469] <= 16'b0000_0000_0000_0000;
array[25470] <= 16'b0000_0000_0000_0000;
array[25471] <= 16'b0000_0000_0000_0000;
array[25472] <= 16'b0000_0000_0000_0000;
array[25473] <= 16'b0000_0000_0000_0000;
array[25474] <= 16'b0000_0000_0000_0000;
array[25475] <= 16'b0000_0000_0000_0000;
array[25476] <= 16'b0000_0000_0000_0000;
array[25477] <= 16'b0000_0000_0000_0000;
array[25478] <= 16'b0000_0000_0000_0000;
array[25479] <= 16'b0000_0000_0000_0000;
array[25480] <= 16'b0000_0000_0000_0000;
array[25481] <= 16'b0000_0000_0000_0000;
array[25482] <= 16'b0000_0000_0000_0000;
array[25483] <= 16'b0000_0000_0000_0000;
array[25484] <= 16'b0000_0000_0000_0000;
array[25485] <= 16'b0000_0000_0000_0000;
array[25486] <= 16'b0000_0000_0000_0000;
array[25487] <= 16'b0000_0000_0000_0000;
array[25488] <= 16'b0000_0000_0000_0000;
array[25489] <= 16'b0000_0000_0000_0000;
array[25490] <= 16'b0000_0000_0000_0000;
array[25491] <= 16'b0000_0000_0000_0000;
array[25492] <= 16'b0000_0000_0000_0000;
array[25493] <= 16'b0000_0000_0000_0000;
array[25494] <= 16'b0000_0000_0000_0000;
array[25495] <= 16'b0000_0000_0000_0000;
array[25496] <= 16'b0000_0000_0000_0000;
array[25497] <= 16'b0000_0000_0000_0000;
array[25498] <= 16'b0000_0000_0000_0000;
array[25499] <= 16'b0000_0000_0000_0000;
array[25500] <= 16'b0000_0000_0000_0000;
array[25501] <= 16'b0000_0000_0000_0000;
array[25502] <= 16'b0000_0000_0000_0000;
array[25503] <= 16'b0000_0000_0000_0000;
array[25504] <= 16'b0000_0000_0000_0000;
array[25505] <= 16'b0000_0000_0000_0000;
array[25506] <= 16'b0000_0000_0000_0000;
array[25507] <= 16'b0000_0000_0000_0000;
array[25508] <= 16'b0000_0000_0000_0000;
array[25509] <= 16'b0000_0000_0000_0000;
array[25510] <= 16'b0000_0000_0000_0000;
array[25511] <= 16'b0000_0000_0000_0000;
array[25512] <= 16'b0000_0000_0000_0000;
array[25513] <= 16'b0000_0000_0000_0000;
array[25514] <= 16'b0000_0000_0000_0000;
array[25515] <= 16'b0000_0000_0000_0000;
array[25516] <= 16'b0000_0000_0000_0000;
array[25517] <= 16'b0000_0000_0000_0000;
array[25518] <= 16'b0000_0000_0000_0000;
array[25519] <= 16'b0000_0000_0000_0000;
array[25520] <= 16'b0000_0000_0000_0000;
array[25521] <= 16'b0000_0000_0000_0000;
array[25522] <= 16'b0000_0000_0000_0000;
array[25523] <= 16'b0000_0000_0000_0000;
array[25524] <= 16'b0000_0000_0000_0000;
array[25525] <= 16'b0000_0000_0000_0000;
array[25526] <= 16'b0000_0000_0000_0000;
array[25527] <= 16'b0000_0000_0000_0000;
array[25528] <= 16'b0000_0000_0000_0000;
array[25529] <= 16'b0000_0000_0000_0000;
array[25530] <= 16'b0000_0000_0000_0000;
array[25531] <= 16'b0000_0000_0000_0000;
array[25532] <= 16'b0000_0000_0000_0000;
array[25533] <= 16'b0000_0000_0000_0000;
array[25534] <= 16'b0000_0000_0000_0000;
array[25535] <= 16'b0000_0000_0000_0000;
array[25536] <= 16'b0000_0000_0000_0000;
array[25537] <= 16'b0000_0000_0000_0000;
array[25538] <= 16'b0000_0000_0000_0000;
array[25539] <= 16'b0000_0000_0000_0000;
array[25540] <= 16'b0000_0000_0000_0000;
array[25541] <= 16'b0000_0000_0000_0000;
array[25542] <= 16'b0000_0000_0000_0000;
array[25543] <= 16'b0000_0000_0000_0000;
array[25544] <= 16'b0000_0000_0000_0000;
array[25545] <= 16'b0000_0000_0000_0000;
array[25546] <= 16'b0000_0000_0000_0000;
array[25547] <= 16'b0000_0000_0000_0000;
array[25548] <= 16'b0000_0000_0000_0000;
array[25549] <= 16'b0000_0000_0000_0000;
array[25550] <= 16'b0000_0000_0000_0000;
array[25551] <= 16'b0000_0000_0000_0000;
array[25552] <= 16'b0000_0000_0000_0000;
array[25553] <= 16'b0000_0000_0000_0000;
array[25554] <= 16'b0000_0000_0000_0000;
array[25555] <= 16'b0000_0000_0000_0000;
array[25556] <= 16'b0000_0000_0000_0000;
array[25557] <= 16'b0000_0000_0000_0000;
array[25558] <= 16'b0000_0000_0000_0000;
array[25559] <= 16'b0000_0000_0000_0000;
array[25560] <= 16'b0000_0000_0000_0000;
array[25561] <= 16'b0000_0000_0000_0000;
array[25562] <= 16'b0000_0000_0000_0000;
array[25563] <= 16'b0000_0000_0000_0000;
array[25564] <= 16'b0000_0000_0000_0000;
array[25565] <= 16'b0000_0000_0000_0000;
array[25566] <= 16'b0000_0000_0000_0000;
array[25567] <= 16'b0000_0000_0000_0000;
array[25568] <= 16'b0000_0000_0000_0000;
array[25569] <= 16'b0000_0000_0000_0000;
array[25570] <= 16'b0000_0000_0000_0000;
array[25571] <= 16'b0000_0000_0000_0000;
array[25572] <= 16'b0000_0000_0000_0000;
array[25573] <= 16'b0000_0000_0000_0000;
array[25574] <= 16'b0000_0000_0000_0000;
array[25575] <= 16'b0000_0000_0000_0000;
array[25576] <= 16'b0000_0000_0000_0000;
array[25577] <= 16'b0000_0000_0000_0000;
array[25578] <= 16'b0000_0000_0000_0000;
array[25579] <= 16'b0000_0000_0000_0000;
array[25580] <= 16'b0000_0000_0000_0000;
array[25581] <= 16'b0000_0000_0000_0000;
array[25582] <= 16'b0000_0000_0000_0000;
array[25583] <= 16'b0000_0000_0000_0000;
array[25584] <= 16'b0000_0000_0000_0000;
array[25585] <= 16'b0000_0000_0000_0000;
array[25586] <= 16'b0000_0000_0000_0000;
array[25587] <= 16'b0000_0000_0000_0000;
array[25588] <= 16'b0000_0000_0000_0000;
array[25589] <= 16'b0000_0000_0000_0000;
array[25590] <= 16'b0000_0000_0000_0000;
array[25591] <= 16'b0000_0000_0000_0000;
array[25592] <= 16'b0000_0000_0000_0000;
array[25593] <= 16'b0000_0000_0000_0000;
array[25594] <= 16'b0000_0000_0000_0000;
array[25595] <= 16'b0000_0000_0000_0000;
array[25596] <= 16'b0000_0000_0000_0000;
array[25597] <= 16'b0000_0000_0000_0000;
array[25598] <= 16'b0000_0000_0000_0000;
array[25599] <= 16'b0000_0000_0000_0000;
array[25600] <= 16'b0000_0000_0000_0000;
array[25601] <= 16'b0000_0000_0000_0000;
array[25602] <= 16'b0000_0000_0000_0000;
array[25603] <= 16'b0000_0000_0000_0000;
array[25604] <= 16'b0000_0000_0000_0000;
array[25605] <= 16'b0000_0000_0000_0000;
array[25606] <= 16'b0000_0000_0000_0000;
array[25607] <= 16'b0000_0000_0000_0000;
array[25608] <= 16'b0000_0000_0000_0000;
array[25609] <= 16'b0000_0000_0000_0000;
array[25610] <= 16'b0000_0000_0000_0000;
array[25611] <= 16'b0000_0000_0000_0000;
array[25612] <= 16'b0000_0000_0000_0000;
array[25613] <= 16'b0000_0000_0000_0000;
array[25614] <= 16'b0000_0000_0000_0000;
array[25615] <= 16'b0000_0000_0000_0000;
array[25616] <= 16'b0000_0000_0000_0000;
array[25617] <= 16'b0000_0000_0000_0000;
array[25618] <= 16'b0000_0000_0000_0000;
array[25619] <= 16'b0000_0000_0000_0000;
array[25620] <= 16'b0000_0000_0000_0000;
array[25621] <= 16'b0000_0000_0000_0000;
array[25622] <= 16'b0000_0000_0000_0000;
array[25623] <= 16'b0000_0000_0000_0000;
array[25624] <= 16'b0000_0000_0000_0000;
array[25625] <= 16'b0000_0000_0000_0000;
array[25626] <= 16'b0000_0000_0000_0000;
array[25627] <= 16'b0000_0000_0000_0000;
array[25628] <= 16'b0000_0000_0000_0000;
array[25629] <= 16'b0000_0000_0000_0000;
array[25630] <= 16'b0000_0000_0000_0000;
array[25631] <= 16'b0000_0000_0000_0000;
array[25632] <= 16'b0000_0000_0000_0000;
array[25633] <= 16'b0000_0000_0000_0000;
array[25634] <= 16'b0000_0000_0000_0000;
array[25635] <= 16'b0000_0000_0000_0000;
array[25636] <= 16'b0000_0000_0000_0000;
array[25637] <= 16'b0000_0000_0000_0000;
array[25638] <= 16'b0000_0000_0000_0000;
array[25639] <= 16'b0000_0000_0000_0000;
array[25640] <= 16'b0000_0000_0000_0000;
array[25641] <= 16'b0000_0000_0000_0000;
array[25642] <= 16'b0000_0000_0000_0000;
array[25643] <= 16'b0000_0000_0000_0000;
array[25644] <= 16'b0000_0000_0000_0000;
array[25645] <= 16'b0000_0000_0000_0000;
array[25646] <= 16'b0000_0000_0000_0000;
array[25647] <= 16'b0000_0000_0000_0000;
array[25648] <= 16'b0000_0000_0000_0000;
array[25649] <= 16'b0000_0000_0000_0000;
array[25650] <= 16'b0000_0000_0000_0000;
array[25651] <= 16'b0000_0000_0000_0000;
array[25652] <= 16'b0000_0000_0000_0000;
array[25653] <= 16'b0000_0000_0000_0000;
array[25654] <= 16'b0000_0000_0000_0000;
array[25655] <= 16'b0000_0000_0000_0000;
array[25656] <= 16'b0000_0000_0000_0000;
array[25657] <= 16'b0000_0000_0000_0000;
array[25658] <= 16'b0000_0000_0000_0000;
array[25659] <= 16'b0000_0000_0000_0000;
array[25660] <= 16'b0000_0000_0000_0000;
array[25661] <= 16'b0000_0000_0000_0000;
array[25662] <= 16'b0000_0000_0000_0000;
array[25663] <= 16'b0000_0000_0000_0000;
array[25664] <= 16'b0000_0000_0000_0000;
array[25665] <= 16'b0000_0000_0000_0000;
array[25666] <= 16'b0000_0000_0000_0000;
array[25667] <= 16'b0000_0000_0000_0000;
array[25668] <= 16'b0000_0000_0000_0000;
array[25669] <= 16'b0000_0000_0000_0000;
array[25670] <= 16'b0000_0000_0000_0000;
array[25671] <= 16'b0000_0000_0000_0000;
array[25672] <= 16'b0000_0000_0000_0000;
array[25673] <= 16'b0000_0000_0000_0000;
array[25674] <= 16'b0000_0000_0000_0000;
array[25675] <= 16'b0000_0000_0000_0000;
array[25676] <= 16'b0000_0000_0000_0000;
array[25677] <= 16'b0000_0000_0000_0000;
array[25678] <= 16'b0000_0000_0000_0000;
array[25679] <= 16'b0000_0000_0000_0000;
array[25680] <= 16'b0000_0000_0000_0000;
array[25681] <= 16'b0000_0000_0000_0000;
array[25682] <= 16'b0000_0000_0000_0000;
array[25683] <= 16'b0000_0000_0000_0000;
array[25684] <= 16'b0000_0000_0000_0000;
array[25685] <= 16'b0000_0000_0000_0000;
array[25686] <= 16'b0000_0000_0000_0000;
array[25687] <= 16'b0000_0000_0000_0000;
array[25688] <= 16'b0000_0000_0000_0000;
array[25689] <= 16'b0000_0000_0000_0000;
array[25690] <= 16'b0000_0000_0000_0000;
array[25691] <= 16'b0000_0000_0000_0000;
array[25692] <= 16'b0000_0000_0000_0000;
array[25693] <= 16'b0000_0000_0000_0000;
array[25694] <= 16'b0000_0000_0000_0000;
array[25695] <= 16'b0000_0000_0000_0000;
array[25696] <= 16'b0000_0000_0000_0000;
array[25697] <= 16'b0000_0000_0000_0000;
array[25698] <= 16'b0000_0000_0000_0000;
array[25699] <= 16'b0000_0000_0000_0000;
array[25700] <= 16'b0000_0000_0000_0000;
array[25701] <= 16'b0000_0000_0000_0000;
array[25702] <= 16'b0000_0000_0000_0000;
array[25703] <= 16'b0000_0000_0000_0000;
array[25704] <= 16'b0000_0000_0000_0000;
array[25705] <= 16'b0000_0000_0000_0000;
array[25706] <= 16'b0000_0000_0000_0000;
array[25707] <= 16'b0000_0000_0000_0000;
array[25708] <= 16'b0000_0000_0000_0000;
array[25709] <= 16'b0000_0000_0000_0000;
array[25710] <= 16'b0000_0000_0000_0000;
array[25711] <= 16'b0000_0000_0000_0000;
array[25712] <= 16'b0000_0000_0000_0000;
array[25713] <= 16'b0000_0000_0000_0000;
array[25714] <= 16'b0000_0000_0000_0000;
array[25715] <= 16'b0000_0000_0000_0000;
array[25716] <= 16'b0000_0000_0000_0000;
array[25717] <= 16'b0000_0000_0000_0000;
array[25718] <= 16'b0000_0000_0000_0000;
array[25719] <= 16'b0000_0000_0000_0000;
array[25720] <= 16'b0000_0000_0000_0000;
array[25721] <= 16'b0000_0000_0000_0000;
array[25722] <= 16'b0000_0000_0000_0000;
array[25723] <= 16'b0000_0000_0000_0000;
array[25724] <= 16'b0000_0000_0000_0000;
array[25725] <= 16'b0000_0000_0000_0000;
array[25726] <= 16'b0000_0000_0000_0000;
array[25727] <= 16'b0000_0000_0000_0000;
array[25728] <= 16'b0000_0000_0000_0000;
array[25729] <= 16'b0000_0000_0000_0000;
array[25730] <= 16'b0000_0000_0000_0000;
array[25731] <= 16'b0000_0000_0000_0000;
array[25732] <= 16'b0000_0000_0000_0000;
array[25733] <= 16'b0000_0000_0000_0000;
array[25734] <= 16'b0000_0000_0000_0000;
array[25735] <= 16'b0000_0000_0000_0000;
array[25736] <= 16'b0000_0000_0000_0000;
array[25737] <= 16'b0000_0000_0000_0000;
array[25738] <= 16'b0000_0000_0000_0000;
array[25739] <= 16'b0000_0000_0000_0000;
array[25740] <= 16'b0000_0000_0000_0000;
array[25741] <= 16'b0000_0000_0000_0000;
array[25742] <= 16'b0000_0000_0000_0000;
array[25743] <= 16'b0000_0000_0000_0000;
array[25744] <= 16'b0000_0000_0000_0000;
array[25745] <= 16'b0000_0000_0000_0000;
array[25746] <= 16'b0000_0000_0000_0000;
array[25747] <= 16'b0000_0000_0000_0000;
array[25748] <= 16'b0000_0000_0000_0000;
array[25749] <= 16'b0000_0000_0000_0000;
array[25750] <= 16'b0000_0000_0000_0000;
array[25751] <= 16'b0000_0000_0000_0000;
array[25752] <= 16'b0000_0000_0000_0000;
array[25753] <= 16'b0000_0000_0000_0000;
array[25754] <= 16'b0000_0000_0000_0000;
array[25755] <= 16'b0000_0000_0000_0000;
array[25756] <= 16'b0000_0000_0000_0000;
array[25757] <= 16'b0000_0000_0000_0000;
array[25758] <= 16'b0000_0000_0000_0000;
array[25759] <= 16'b0000_0000_0000_0000;
array[25760] <= 16'b0000_0000_0000_0000;
array[25761] <= 16'b0000_0000_0000_0000;
array[25762] <= 16'b0000_0000_0000_0000;
array[25763] <= 16'b0000_0000_0000_0000;
array[25764] <= 16'b0000_0000_0000_0000;
array[25765] <= 16'b0000_0000_0000_0000;
array[25766] <= 16'b0000_0000_0000_0000;
array[25767] <= 16'b0000_0000_0000_0000;
array[25768] <= 16'b0000_0000_0000_0000;
array[25769] <= 16'b0000_0000_0000_0000;
array[25770] <= 16'b0000_0000_0000_0000;
array[25771] <= 16'b0000_0000_0000_0000;
array[25772] <= 16'b0000_0000_0000_0000;
array[25773] <= 16'b0000_0000_0000_0000;
array[25774] <= 16'b0000_0000_0000_0000;
array[25775] <= 16'b0000_0000_0000_0000;
array[25776] <= 16'b0000_0000_0000_0000;
array[25777] <= 16'b0000_0000_0000_0000;
array[25778] <= 16'b0000_0000_0000_0000;
array[25779] <= 16'b0000_0000_0000_0000;
array[25780] <= 16'b0000_0000_0000_0000;
array[25781] <= 16'b0000_0000_0000_0000;
array[25782] <= 16'b0000_0000_0000_0000;
array[25783] <= 16'b0000_0000_0000_0000;
array[25784] <= 16'b0000_0000_0000_0000;
array[25785] <= 16'b0000_0000_0000_0000;
array[25786] <= 16'b0000_0000_0000_0000;
array[25787] <= 16'b0000_0000_0000_0000;
array[25788] <= 16'b0000_0000_0000_0000;
array[25789] <= 16'b0000_0000_0000_0000;
array[25790] <= 16'b0000_0000_0000_0000;
array[25791] <= 16'b0000_0000_0000_0000;
array[25792] <= 16'b0000_0000_0000_0000;
array[25793] <= 16'b0000_0000_0000_0000;
array[25794] <= 16'b0000_0000_0000_0000;
array[25795] <= 16'b0000_0000_0000_0000;
array[25796] <= 16'b0000_0000_0000_0000;
array[25797] <= 16'b0000_0000_0000_0000;
array[25798] <= 16'b0000_0000_0000_0000;
array[25799] <= 16'b0000_0000_0000_0000;
array[25800] <= 16'b0000_0000_0000_0000;
array[25801] <= 16'b0000_0000_0000_0000;
array[25802] <= 16'b0000_0000_0000_0000;
array[25803] <= 16'b0000_0000_0000_0000;
array[25804] <= 16'b0000_0000_0000_0000;
array[25805] <= 16'b0000_0000_0000_0000;
array[25806] <= 16'b0000_0000_0000_0000;
array[25807] <= 16'b0000_0000_0000_0000;
array[25808] <= 16'b0000_0000_0000_0000;
array[25809] <= 16'b0000_0000_0000_0000;
array[25810] <= 16'b0000_0000_0000_0000;
array[25811] <= 16'b0000_0000_0000_0000;
array[25812] <= 16'b0000_0000_0000_0000;
array[25813] <= 16'b0000_0000_0000_0000;
array[25814] <= 16'b0000_0000_0000_0000;
array[25815] <= 16'b0000_0000_0000_0000;
array[25816] <= 16'b0000_0000_0000_0000;
array[25817] <= 16'b0000_0000_0000_0000;
array[25818] <= 16'b0000_0000_0000_0000;
array[25819] <= 16'b0000_0000_0000_0000;
array[25820] <= 16'b0000_0000_0000_0000;
array[25821] <= 16'b0000_0000_0000_0000;
array[25822] <= 16'b0000_0000_0000_0000;
array[25823] <= 16'b0000_0000_0000_0000;
array[25824] <= 16'b0000_0000_0000_0000;
array[25825] <= 16'b0000_0000_0000_0000;
array[25826] <= 16'b0000_0000_0000_0000;
array[25827] <= 16'b0000_0000_0000_0000;
array[25828] <= 16'b0000_0000_0000_0000;
array[25829] <= 16'b0000_0000_0000_0000;
array[25830] <= 16'b0000_0000_0000_0000;
array[25831] <= 16'b0000_0000_0000_0000;
array[25832] <= 16'b0000_0000_0000_0000;
array[25833] <= 16'b0000_0000_0000_0000;
array[25834] <= 16'b0000_0000_0000_0000;
array[25835] <= 16'b0000_0000_0000_0000;
array[25836] <= 16'b0000_0000_0000_0000;
array[25837] <= 16'b0000_0000_0000_0000;
array[25838] <= 16'b0000_0000_0000_0000;
array[25839] <= 16'b0000_0000_0000_0000;
array[25840] <= 16'b0000_0000_0000_0000;
array[25841] <= 16'b0000_0000_0000_0000;
array[25842] <= 16'b0000_0000_0000_0000;
array[25843] <= 16'b0000_0000_0000_0000;
array[25844] <= 16'b0000_0000_0000_0000;
array[25845] <= 16'b0000_0000_0000_0000;
array[25846] <= 16'b0000_0000_0000_0000;
array[25847] <= 16'b0000_0000_0000_0000;
array[25848] <= 16'b0000_0000_0000_0000;
array[25849] <= 16'b0000_0000_0000_0000;
array[25850] <= 16'b0000_0000_0000_0000;
array[25851] <= 16'b0000_0000_0000_0000;
array[25852] <= 16'b0000_0000_0000_0000;
array[25853] <= 16'b0000_0000_0000_0000;
array[25854] <= 16'b0000_0000_0000_0000;
array[25855] <= 16'b0000_0000_0000_0000;
array[25856] <= 16'b0000_0000_0000_0000;
array[25857] <= 16'b0000_0000_0000_0000;
array[25858] <= 16'b0000_0000_0000_0000;
array[25859] <= 16'b0000_0000_0000_0000;
array[25860] <= 16'b0000_0000_0000_0000;
array[25861] <= 16'b0000_0000_0000_0000;
array[25862] <= 16'b0000_0000_0000_0000;
array[25863] <= 16'b0000_0000_0000_0000;
array[25864] <= 16'b0000_0000_0000_0000;
array[25865] <= 16'b0000_0000_0000_0000;
array[25866] <= 16'b0000_0000_0000_0000;
array[25867] <= 16'b0000_0000_0000_0000;
array[25868] <= 16'b0000_0000_0000_0000;
array[25869] <= 16'b0000_0000_0000_0000;
array[25870] <= 16'b0000_0000_0000_0000;
array[25871] <= 16'b0000_0000_0000_0000;
array[25872] <= 16'b0000_0000_0000_0000;
array[25873] <= 16'b0000_0000_0000_0000;
array[25874] <= 16'b0000_0000_0000_0000;
array[25875] <= 16'b0000_0000_0000_0000;
array[25876] <= 16'b0000_0000_0000_0000;
array[25877] <= 16'b0000_0000_0000_0000;
array[25878] <= 16'b0000_0000_0000_0000;
array[25879] <= 16'b0000_0000_0000_0000;
array[25880] <= 16'b0000_0000_0000_0000;
array[25881] <= 16'b0000_0000_0000_0000;
array[25882] <= 16'b0000_0000_0000_0000;
array[25883] <= 16'b0000_0000_0000_0000;
array[25884] <= 16'b0000_0000_0000_0000;
array[25885] <= 16'b0000_0000_0000_0000;
array[25886] <= 16'b0000_0000_0000_0000;
array[25887] <= 16'b0000_0000_0000_0000;
array[25888] <= 16'b0000_0000_0000_0000;
array[25889] <= 16'b0000_0000_0000_0000;
array[25890] <= 16'b0000_0000_0000_0000;
array[25891] <= 16'b0000_0000_0000_0000;
array[25892] <= 16'b0000_0000_0000_0000;
array[25893] <= 16'b0000_0000_0000_0000;
array[25894] <= 16'b0000_0000_0000_0000;
array[25895] <= 16'b0000_0000_0000_0000;
array[25896] <= 16'b0000_0000_0000_0000;
array[25897] <= 16'b0000_0000_0000_0000;
array[25898] <= 16'b0000_0000_0000_0000;
array[25899] <= 16'b0000_0000_0000_0000;
array[25900] <= 16'b0000_0000_0000_0000;
array[25901] <= 16'b0000_0000_0000_0000;
array[25902] <= 16'b0000_0000_0000_0000;
array[25903] <= 16'b0000_0000_0000_0000;
array[25904] <= 16'b0000_0000_0000_0000;
array[25905] <= 16'b0000_0000_0000_0000;
array[25906] <= 16'b0000_0000_0000_0000;
array[25907] <= 16'b0000_0000_0000_0000;
array[25908] <= 16'b0000_0000_0000_0000;
array[25909] <= 16'b0000_0000_0000_0000;
array[25910] <= 16'b0000_0000_0000_0000;
array[25911] <= 16'b0000_0000_0000_0000;
array[25912] <= 16'b0000_0000_0000_0000;
array[25913] <= 16'b0000_0000_0000_0000;
array[25914] <= 16'b0000_0000_0000_0000;
array[25915] <= 16'b0000_0000_0000_0000;
array[25916] <= 16'b0000_0000_0000_0000;
array[25917] <= 16'b0000_0000_0000_0000;
array[25918] <= 16'b0000_0000_0000_0000;
array[25919] <= 16'b0000_0000_0000_0000;
array[25920] <= 16'b0000_0000_0000_0000;
array[25921] <= 16'b0000_0000_0000_0000;
array[25922] <= 16'b0000_0000_0000_0000;
array[25923] <= 16'b0000_0000_0000_0000;
array[25924] <= 16'b0000_0000_0000_0000;
array[25925] <= 16'b0000_0000_0000_0000;
array[25926] <= 16'b0000_0000_0000_0000;
array[25927] <= 16'b0000_0000_0000_0000;
array[25928] <= 16'b0000_0000_0000_0000;
array[25929] <= 16'b0000_0000_0000_0000;
array[25930] <= 16'b0000_0000_0000_0000;
array[25931] <= 16'b0000_0000_0000_0000;
array[25932] <= 16'b0000_0000_0000_0000;
array[25933] <= 16'b0000_0000_0000_0000;
array[25934] <= 16'b0000_0000_0000_0000;
array[25935] <= 16'b0000_0000_0000_0000;
array[25936] <= 16'b0000_0000_0000_0000;
array[25937] <= 16'b0000_0000_0000_0000;
array[25938] <= 16'b0000_0000_0000_0000;
array[25939] <= 16'b0000_0000_0000_0000;
array[25940] <= 16'b0000_0000_0000_0000;
array[25941] <= 16'b0000_0000_0000_0000;
array[25942] <= 16'b0000_0000_0000_0000;
array[25943] <= 16'b0000_0000_0000_0000;
array[25944] <= 16'b0000_0000_0000_0000;
array[25945] <= 16'b0000_0000_0000_0000;
array[25946] <= 16'b0000_0000_0000_0000;
array[25947] <= 16'b0000_0000_0000_0000;
array[25948] <= 16'b0000_0000_0000_0000;
array[25949] <= 16'b0000_0000_0000_0000;
array[25950] <= 16'b0000_0000_0000_0000;
array[25951] <= 16'b0000_0000_0000_0000;
array[25952] <= 16'b0000_0000_0000_0000;
array[25953] <= 16'b0000_0000_0000_0000;
array[25954] <= 16'b0000_0000_0000_0000;
array[25955] <= 16'b0000_0000_0000_0000;
array[25956] <= 16'b0000_0000_0000_0000;
array[25957] <= 16'b0000_0000_0000_0000;
array[25958] <= 16'b0000_0000_0000_0000;
array[25959] <= 16'b0000_0000_0000_0000;
array[25960] <= 16'b0000_0000_0000_0000;
array[25961] <= 16'b0000_0000_0000_0000;
array[25962] <= 16'b0000_0000_0000_0000;
array[25963] <= 16'b0000_0000_0000_0000;
array[25964] <= 16'b0000_0000_0000_0000;
array[25965] <= 16'b0000_0000_0000_0000;
array[25966] <= 16'b0000_0000_0000_0000;
array[25967] <= 16'b0000_0000_0000_0000;
array[25968] <= 16'b0000_0000_0000_0000;
array[25969] <= 16'b0000_0000_0000_0000;
array[25970] <= 16'b0000_0000_0000_0000;
array[25971] <= 16'b0000_0000_0000_0000;
array[25972] <= 16'b0000_0000_0000_0000;
array[25973] <= 16'b0000_0000_0000_0000;
array[25974] <= 16'b0000_0000_0000_0000;
array[25975] <= 16'b0000_0000_0000_0000;
array[25976] <= 16'b0000_0000_0000_0000;
array[25977] <= 16'b0000_0000_0000_0000;
array[25978] <= 16'b0000_0000_0000_0000;
array[25979] <= 16'b0000_0000_0000_0000;
array[25980] <= 16'b0000_0000_0000_0000;
array[25981] <= 16'b0000_0000_0000_0000;
array[25982] <= 16'b0000_0000_0000_0000;
array[25983] <= 16'b0000_0000_0000_0000;
array[25984] <= 16'b0000_0000_0000_0000;
array[25985] <= 16'b0000_0000_0000_0000;
array[25986] <= 16'b0000_0000_0000_0000;
array[25987] <= 16'b0000_0000_0000_0000;
array[25988] <= 16'b0000_0000_0000_0000;
array[25989] <= 16'b0000_0000_0000_0000;
array[25990] <= 16'b0000_0000_0000_0000;
array[25991] <= 16'b0000_0000_0000_0000;
array[25992] <= 16'b0000_0000_0000_0000;
array[25993] <= 16'b0000_0000_0000_0000;
array[25994] <= 16'b0000_0000_0000_0000;
array[25995] <= 16'b0000_0000_0000_0000;
array[25996] <= 16'b0000_0000_0000_0000;
array[25997] <= 16'b0000_0000_0000_0000;
array[25998] <= 16'b0000_0000_0000_0000;
array[25999] <= 16'b0000_0000_0000_0000;
array[26000] <= 16'b0000_0000_0000_0000;
array[26001] <= 16'b0000_0000_0000_0000;
array[26002] <= 16'b0000_0000_0000_0000;
array[26003] <= 16'b0000_0000_0000_0000;
array[26004] <= 16'b0000_0000_0000_0000;
array[26005] <= 16'b0000_0000_0000_0000;
array[26006] <= 16'b0000_0000_0000_0000;
array[26007] <= 16'b0000_0000_0000_0000;
array[26008] <= 16'b0000_0000_0000_0000;
array[26009] <= 16'b0000_0000_0000_0000;
array[26010] <= 16'b0000_0000_0000_0000;
array[26011] <= 16'b0000_0000_0000_0000;
array[26012] <= 16'b0000_0000_0000_0000;
array[26013] <= 16'b0000_0000_0000_0000;
array[26014] <= 16'b0000_0000_0000_0000;
array[26015] <= 16'b0000_0000_0000_0000;
array[26016] <= 16'b0000_0000_0000_0000;
array[26017] <= 16'b0000_0000_0000_0000;
array[26018] <= 16'b0000_0000_0000_0000;
array[26019] <= 16'b0000_0000_0000_0000;
array[26020] <= 16'b0000_0000_0000_0000;
array[26021] <= 16'b0000_0000_0000_0000;
array[26022] <= 16'b0000_0000_0000_0000;
array[26023] <= 16'b0000_0000_0000_0000;
array[26024] <= 16'b0000_0000_0000_0000;
array[26025] <= 16'b0000_0000_0000_0000;
array[26026] <= 16'b0000_0000_0000_0000;
array[26027] <= 16'b0000_0000_0000_0000;
array[26028] <= 16'b0000_0000_0000_0000;
array[26029] <= 16'b0000_0000_0000_0000;
array[26030] <= 16'b0000_0000_0000_0000;
array[26031] <= 16'b0000_0000_0000_0000;
array[26032] <= 16'b0000_0000_0000_0000;
array[26033] <= 16'b0000_0000_0000_0000;
array[26034] <= 16'b0000_0000_0000_0000;
array[26035] <= 16'b0000_0000_0000_0000;
array[26036] <= 16'b0000_0000_0000_0000;
array[26037] <= 16'b0000_0000_0000_0000;
array[26038] <= 16'b0000_0000_0000_0000;
array[26039] <= 16'b0000_0000_0000_0000;
array[26040] <= 16'b0000_0000_0000_0000;
array[26041] <= 16'b0000_0000_0000_0000;
array[26042] <= 16'b0000_0000_0000_0000;
array[26043] <= 16'b0000_0000_0000_0000;
array[26044] <= 16'b0000_0000_0000_0000;
array[26045] <= 16'b0000_0000_0000_0000;
array[26046] <= 16'b0000_0000_0000_0000;
array[26047] <= 16'b0000_0000_0000_0000;
array[26048] <= 16'b0000_0000_0000_0000;
array[26049] <= 16'b0000_0000_0000_0000;
array[26050] <= 16'b0000_0000_0000_0000;
array[26051] <= 16'b0000_0000_0000_0000;
array[26052] <= 16'b0000_0000_0000_0000;
array[26053] <= 16'b0000_0000_0000_0000;
array[26054] <= 16'b0000_0000_0000_0000;
array[26055] <= 16'b0000_0000_0000_0000;
array[26056] <= 16'b0000_0000_0000_0000;
array[26057] <= 16'b0000_0000_0000_0000;
array[26058] <= 16'b0000_0000_0000_0000;
array[26059] <= 16'b0000_0000_0000_0000;
array[26060] <= 16'b0000_0000_0000_0000;
array[26061] <= 16'b0000_0000_0000_0000;
array[26062] <= 16'b0000_0000_0000_0000;
array[26063] <= 16'b0000_0000_0000_0000;
array[26064] <= 16'b0000_0000_0000_0000;
array[26065] <= 16'b0000_0000_0000_0000;
array[26066] <= 16'b0000_0000_0000_0000;
array[26067] <= 16'b0000_0000_0000_0000;
array[26068] <= 16'b0000_0000_0000_0000;
array[26069] <= 16'b0000_0000_0000_0000;
array[26070] <= 16'b0000_0000_0000_0000;
array[26071] <= 16'b0000_0000_0000_0000;
array[26072] <= 16'b0000_0000_0000_0000;
array[26073] <= 16'b0000_0000_0000_0000;
array[26074] <= 16'b0000_0000_0000_0000;
array[26075] <= 16'b0000_0000_0000_0000;
array[26076] <= 16'b0000_0000_0000_0000;
array[26077] <= 16'b0000_0000_0000_0000;
array[26078] <= 16'b0000_0000_0000_0000;
array[26079] <= 16'b0000_0000_0000_0000;
array[26080] <= 16'b0000_0000_0000_0000;
array[26081] <= 16'b0000_0000_0000_0000;
array[26082] <= 16'b0000_0000_0000_0000;
array[26083] <= 16'b0000_0000_0000_0000;
array[26084] <= 16'b0000_0000_0000_0000;
array[26085] <= 16'b0000_0000_0000_0000;
array[26086] <= 16'b0000_0000_0000_0000;
array[26087] <= 16'b0000_0000_0000_0000;
array[26088] <= 16'b0000_0000_0000_0000;
array[26089] <= 16'b0000_0000_0000_0000;
array[26090] <= 16'b0000_0000_0000_0000;
array[26091] <= 16'b0000_0000_0000_0000;
array[26092] <= 16'b0000_0000_0000_0000;
array[26093] <= 16'b0000_0000_0000_0000;
array[26094] <= 16'b0000_0000_0000_0000;
array[26095] <= 16'b0000_0000_0000_0000;
array[26096] <= 16'b0000_0000_0000_0000;
array[26097] <= 16'b0000_0000_0000_0000;
array[26098] <= 16'b0000_0000_0000_0000;
array[26099] <= 16'b0000_0000_0000_0000;
array[26100] <= 16'b0000_0000_0000_0000;
array[26101] <= 16'b0000_0000_0000_0000;
array[26102] <= 16'b0000_0000_0000_0000;
array[26103] <= 16'b0000_0000_0000_0000;
array[26104] <= 16'b0000_0000_0000_0000;
array[26105] <= 16'b0000_0000_0000_0000;
array[26106] <= 16'b0000_0000_0000_0000;
array[26107] <= 16'b0000_0000_0000_0000;
array[26108] <= 16'b0000_0000_0000_0000;
array[26109] <= 16'b0000_0000_0000_0000;
array[26110] <= 16'b0000_0000_0000_0000;
array[26111] <= 16'b0000_0000_0000_0000;
array[26112] <= 16'b0000_0000_0000_0000;
array[26113] <= 16'b0000_0000_0000_0000;
array[26114] <= 16'b0000_0000_0000_0000;
array[26115] <= 16'b0000_0000_0000_0000;
array[26116] <= 16'b0000_0000_0000_0000;
array[26117] <= 16'b0000_0000_0000_0000;
array[26118] <= 16'b0000_0000_0000_0000;
array[26119] <= 16'b0000_0000_0000_0000;
array[26120] <= 16'b0000_0000_0000_0000;
array[26121] <= 16'b0000_0000_0000_0000;
array[26122] <= 16'b0000_0000_0000_0000;
array[26123] <= 16'b0000_0000_0000_0000;
array[26124] <= 16'b0000_0000_0000_0000;
array[26125] <= 16'b0000_0000_0000_0000;
array[26126] <= 16'b0000_0000_0000_0000;
array[26127] <= 16'b0000_0000_0000_0000;
array[26128] <= 16'b0000_0000_0000_0000;
array[26129] <= 16'b0000_0000_0000_0000;
array[26130] <= 16'b0000_0000_0000_0000;
array[26131] <= 16'b0000_0000_0000_0000;
array[26132] <= 16'b0000_0000_0000_0000;
array[26133] <= 16'b0000_0000_0000_0000;
array[26134] <= 16'b0000_0000_0000_0000;
array[26135] <= 16'b0000_0000_0000_0000;
array[26136] <= 16'b0000_0000_0000_0000;
array[26137] <= 16'b0000_0000_0000_0000;
array[26138] <= 16'b0000_0000_0000_0000;
array[26139] <= 16'b0000_0000_0000_0000;
array[26140] <= 16'b0000_0000_0000_0000;
array[26141] <= 16'b0000_0000_0000_0000;
array[26142] <= 16'b0000_0000_0000_0000;
array[26143] <= 16'b0000_0000_0000_0000;
array[26144] <= 16'b0000_0000_0000_0000;
array[26145] <= 16'b0000_0000_0000_0000;
array[26146] <= 16'b0000_0000_0000_0000;
array[26147] <= 16'b0000_0000_0000_0000;
array[26148] <= 16'b0000_0000_0000_0000;
array[26149] <= 16'b0000_0000_0000_0000;
array[26150] <= 16'b0000_0000_0000_0000;
array[26151] <= 16'b0000_0000_0000_0000;
array[26152] <= 16'b0000_0000_0000_0000;
array[26153] <= 16'b0000_0000_0000_0000;
array[26154] <= 16'b0000_0000_0000_0000;
array[26155] <= 16'b0000_0000_0000_0000;
array[26156] <= 16'b0000_0000_0000_0000;
array[26157] <= 16'b0000_0000_0000_0000;
array[26158] <= 16'b0000_0000_0000_0000;
array[26159] <= 16'b0000_0000_0000_0000;
array[26160] <= 16'b0000_0000_0000_0000;
array[26161] <= 16'b0000_0000_0000_0000;
array[26162] <= 16'b0000_0000_0000_0000;
array[26163] <= 16'b0000_0000_0000_0000;
array[26164] <= 16'b0000_0000_0000_0000;
array[26165] <= 16'b0000_0000_0000_0000;
array[26166] <= 16'b0000_0000_0000_0000;
array[26167] <= 16'b0000_0000_0000_0000;
array[26168] <= 16'b0000_0000_0000_0000;
array[26169] <= 16'b0000_0000_0000_0000;
array[26170] <= 16'b0000_0000_0000_0000;
array[26171] <= 16'b0000_0000_0000_0000;
array[26172] <= 16'b0000_0000_0000_0000;
array[26173] <= 16'b0000_0000_0000_0000;
array[26174] <= 16'b0000_0000_0000_0000;
array[26175] <= 16'b0000_0000_0000_0000;
array[26176] <= 16'b0000_0000_0000_0000;
array[26177] <= 16'b0000_0000_0000_0000;
array[26178] <= 16'b0000_0000_0000_0000;
array[26179] <= 16'b0000_0000_0000_0000;
array[26180] <= 16'b0000_0000_0000_0000;
array[26181] <= 16'b0000_0000_0000_0000;
array[26182] <= 16'b0000_0000_0000_0000;
array[26183] <= 16'b0000_0000_0000_0000;
array[26184] <= 16'b0000_0000_0000_0000;
array[26185] <= 16'b0000_0000_0000_0000;
array[26186] <= 16'b0000_0000_0000_0000;
array[26187] <= 16'b0000_0000_0000_0000;
array[26188] <= 16'b0000_0000_0000_0000;
array[26189] <= 16'b0000_0000_0000_0000;
array[26190] <= 16'b0000_0000_0000_0000;
array[26191] <= 16'b0000_0000_0000_0000;
array[26192] <= 16'b0000_0000_0000_0000;
array[26193] <= 16'b0000_0000_0000_0000;
array[26194] <= 16'b0000_0000_0000_0000;
array[26195] <= 16'b0000_0000_0000_0000;
array[26196] <= 16'b0000_0000_0000_0000;
array[26197] <= 16'b0000_0000_0000_0000;
array[26198] <= 16'b0000_0000_0000_0000;
array[26199] <= 16'b0000_0000_0000_0000;
array[26200] <= 16'b0000_0000_0000_0000;
array[26201] <= 16'b0000_0000_0000_0000;
array[26202] <= 16'b0000_0000_0000_0000;
array[26203] <= 16'b0000_0000_0000_0000;
array[26204] <= 16'b0000_0000_0000_0000;
array[26205] <= 16'b0000_0000_0000_0000;
array[26206] <= 16'b0000_0000_0000_0000;
array[26207] <= 16'b0000_0000_0000_0000;
array[26208] <= 16'b0000_0000_0000_0000;
array[26209] <= 16'b0000_0000_0000_0000;
array[26210] <= 16'b0000_0000_0000_0000;
array[26211] <= 16'b0000_0000_0000_0000;
array[26212] <= 16'b0000_0000_0000_0000;
array[26213] <= 16'b0000_0000_0000_0000;
array[26214] <= 16'b0000_0000_0000_0000;
array[26215] <= 16'b0000_0000_0000_0000;
array[26216] <= 16'b0000_0000_0000_0000;
array[26217] <= 16'b0000_0000_0000_0000;
array[26218] <= 16'b0000_0000_0000_0000;
array[26219] <= 16'b0000_0000_0000_0000;
array[26220] <= 16'b0000_0000_0000_0000;
array[26221] <= 16'b0000_0000_0000_0000;
array[26222] <= 16'b0000_0000_0000_0000;
array[26223] <= 16'b0000_0000_0000_0000;
array[26224] <= 16'b0000_0000_0000_0000;
array[26225] <= 16'b0000_0000_0000_0000;
array[26226] <= 16'b0000_0000_0000_0000;
array[26227] <= 16'b0000_0000_0000_0000;
array[26228] <= 16'b0000_0000_0000_0000;
array[26229] <= 16'b0000_0000_0000_0000;
array[26230] <= 16'b0000_0000_0000_0000;
array[26231] <= 16'b0000_0000_0000_0000;
array[26232] <= 16'b0000_0000_0000_0000;
array[26233] <= 16'b0000_0000_0000_0000;
array[26234] <= 16'b0000_0000_0000_0000;
array[26235] <= 16'b0000_0000_0000_0000;
array[26236] <= 16'b0000_0000_0000_0000;
array[26237] <= 16'b0000_0000_0000_0000;
array[26238] <= 16'b0000_0000_0000_0000;
array[26239] <= 16'b0000_0000_0000_0000;
array[26240] <= 16'b0000_0000_0000_0000;
array[26241] <= 16'b0000_0000_0000_0000;
array[26242] <= 16'b0000_0000_0000_0000;
array[26243] <= 16'b0000_0000_0000_0000;
array[26244] <= 16'b0000_0000_0000_0000;
array[26245] <= 16'b0000_0000_0000_0000;
array[26246] <= 16'b0000_0000_0000_0000;
array[26247] <= 16'b0000_0000_0000_0000;
array[26248] <= 16'b0000_0000_0000_0000;
array[26249] <= 16'b0000_0000_0000_0000;
array[26250] <= 16'b0000_0000_0000_0000;
array[26251] <= 16'b0000_0000_0000_0000;
array[26252] <= 16'b0000_0000_0000_0000;
array[26253] <= 16'b0000_0000_0000_0000;
array[26254] <= 16'b0000_0000_0000_0000;
array[26255] <= 16'b0000_0000_0000_0000;
array[26256] <= 16'b0000_0000_0000_0000;
array[26257] <= 16'b0000_0000_0000_0000;
array[26258] <= 16'b0000_0000_0000_0000;
array[26259] <= 16'b0000_0000_0000_0000;
array[26260] <= 16'b0000_0000_0000_0000;
array[26261] <= 16'b0000_0000_0000_0000;
array[26262] <= 16'b0000_0000_0000_0000;
array[26263] <= 16'b0000_0000_0000_0000;
array[26264] <= 16'b0000_0000_0000_0000;
array[26265] <= 16'b0000_0000_0000_0000;
array[26266] <= 16'b0000_0000_0000_0000;
array[26267] <= 16'b0000_0000_0000_0000;
array[26268] <= 16'b0000_0000_0000_0000;
array[26269] <= 16'b0000_0000_0000_0000;
array[26270] <= 16'b0000_0000_0000_0000;
array[26271] <= 16'b0000_0000_0000_0000;
array[26272] <= 16'b0000_0000_0000_0000;
array[26273] <= 16'b0000_0000_0000_0000;
array[26274] <= 16'b0000_0000_0000_0000;
array[26275] <= 16'b0000_0000_0000_0000;
array[26276] <= 16'b0000_0000_0000_0000;
array[26277] <= 16'b0000_0000_0000_0000;
array[26278] <= 16'b0000_0000_0000_0000;
array[26279] <= 16'b0000_0000_0000_0000;
array[26280] <= 16'b0000_0000_0000_0000;
array[26281] <= 16'b0000_0000_0000_0000;
array[26282] <= 16'b0000_0000_0000_0000;
array[26283] <= 16'b0000_0000_0000_0000;
array[26284] <= 16'b0000_0000_0000_0000;
array[26285] <= 16'b0000_0000_0000_0000;
array[26286] <= 16'b0000_0000_0000_0000;
array[26287] <= 16'b0000_0000_0000_0000;
array[26288] <= 16'b0000_0000_0000_0000;
array[26289] <= 16'b0000_0000_0000_0000;
array[26290] <= 16'b0000_0000_0000_0000;
array[26291] <= 16'b0000_0000_0000_0000;
array[26292] <= 16'b0000_0000_0000_0000;
array[26293] <= 16'b0000_0000_0000_0000;
array[26294] <= 16'b0000_0000_0000_0000;
array[26295] <= 16'b0000_0000_0000_0000;
array[26296] <= 16'b0000_0000_0000_0000;
array[26297] <= 16'b0000_0000_0000_0000;
array[26298] <= 16'b0000_0000_0000_0000;
array[26299] <= 16'b0000_0000_0000_0000;
array[26300] <= 16'b0000_0000_0000_0000;
array[26301] <= 16'b0000_0000_0000_0000;
array[26302] <= 16'b0000_0000_0000_0000;
array[26303] <= 16'b0000_0000_0000_0000;
array[26304] <= 16'b0000_0000_0000_0000;
array[26305] <= 16'b0000_0000_0000_0000;
array[26306] <= 16'b0000_0000_0000_0000;
array[26307] <= 16'b0000_0000_0000_0000;
array[26308] <= 16'b0000_0000_0000_0000;
array[26309] <= 16'b0000_0000_0000_0000;
array[26310] <= 16'b0000_0000_0000_0000;
array[26311] <= 16'b0000_0000_0000_0000;
array[26312] <= 16'b0000_0000_0000_0000;
array[26313] <= 16'b0000_0000_0000_0000;
array[26314] <= 16'b0000_0000_0000_0000;
array[26315] <= 16'b0000_0000_0000_0000;
array[26316] <= 16'b0000_0000_0000_0000;
array[26317] <= 16'b0000_0000_0000_0000;
array[26318] <= 16'b0000_0000_0000_0000;
array[26319] <= 16'b0000_0000_0000_0000;
array[26320] <= 16'b0000_0000_0000_0000;
array[26321] <= 16'b0000_0000_0000_0000;
array[26322] <= 16'b0000_0000_0000_0000;
array[26323] <= 16'b0000_0000_0000_0000;
array[26324] <= 16'b0000_0000_0000_0000;
array[26325] <= 16'b0000_0000_0000_0000;
array[26326] <= 16'b0000_0000_0000_0000;
array[26327] <= 16'b0000_0000_0000_0000;
array[26328] <= 16'b0000_0000_0000_0000;
array[26329] <= 16'b0000_0000_0000_0000;
array[26330] <= 16'b0000_0000_0000_0000;
array[26331] <= 16'b0000_0000_0000_0000;
array[26332] <= 16'b0000_0000_0000_0000;
array[26333] <= 16'b0000_0000_0000_0000;
array[26334] <= 16'b0000_0000_0000_0000;
array[26335] <= 16'b0000_0000_0000_0000;
array[26336] <= 16'b0000_0000_0000_0000;
array[26337] <= 16'b0000_0000_0000_0000;
array[26338] <= 16'b0000_0000_0000_0000;
array[26339] <= 16'b0000_0000_0000_0000;
array[26340] <= 16'b0000_0000_0000_0000;
array[26341] <= 16'b0000_0000_0000_0000;
array[26342] <= 16'b0000_0000_0000_0000;
array[26343] <= 16'b0000_0000_0000_0000;
array[26344] <= 16'b0000_0000_0000_0000;
array[26345] <= 16'b0000_0000_0000_0000;
array[26346] <= 16'b0000_0000_0000_0000;
array[26347] <= 16'b0000_0000_0000_0000;
array[26348] <= 16'b0000_0000_0000_0000;
array[26349] <= 16'b0000_0000_0000_0000;
array[26350] <= 16'b0000_0000_0000_0000;
array[26351] <= 16'b0000_0000_0000_0000;
array[26352] <= 16'b0000_0000_0000_0000;
array[26353] <= 16'b0000_0000_0000_0000;
array[26354] <= 16'b0000_0000_0000_0000;
array[26355] <= 16'b0000_0000_0000_0000;
array[26356] <= 16'b0000_0000_0000_0000;
array[26357] <= 16'b0000_0000_0000_0000;
array[26358] <= 16'b0000_0000_0000_0000;
array[26359] <= 16'b0000_0000_0000_0000;
array[26360] <= 16'b0000_0000_0000_0000;
array[26361] <= 16'b0000_0000_0000_0000;
array[26362] <= 16'b0000_0000_0000_0000;
array[26363] <= 16'b0000_0000_0000_0000;
array[26364] <= 16'b0000_0000_0000_0000;
array[26365] <= 16'b0000_0000_0000_0000;
array[26366] <= 16'b0000_0000_0000_0000;
array[26367] <= 16'b0000_0000_0000_0000;
array[26368] <= 16'b0000_0000_0000_0000;
array[26369] <= 16'b0000_0000_0000_0000;
array[26370] <= 16'b0000_0000_0000_0000;
array[26371] <= 16'b0000_0000_0000_0000;
array[26372] <= 16'b0000_0000_0000_0000;
array[26373] <= 16'b0000_0000_0000_0000;
array[26374] <= 16'b0000_0000_0000_0000;
array[26375] <= 16'b0000_0000_0000_0000;
array[26376] <= 16'b0000_0000_0000_0000;
array[26377] <= 16'b0000_0000_0000_0000;
array[26378] <= 16'b0000_0000_0000_0000;
array[26379] <= 16'b0000_0000_0000_0000;
array[26380] <= 16'b0000_0000_0000_0000;
array[26381] <= 16'b0000_0000_0000_0000;
array[26382] <= 16'b0000_0000_0000_0000;
array[26383] <= 16'b0000_0000_0000_0000;
array[26384] <= 16'b0000_0000_0000_0000;
array[26385] <= 16'b0000_0000_0000_0000;
array[26386] <= 16'b0000_0000_0000_0000;
array[26387] <= 16'b0000_0000_0000_0000;
array[26388] <= 16'b0000_0000_0000_0000;
array[26389] <= 16'b0000_0000_0000_0000;
array[26390] <= 16'b0000_0000_0000_0000;
array[26391] <= 16'b0000_0000_0000_0000;
array[26392] <= 16'b0000_0000_0000_0000;
array[26393] <= 16'b0000_0000_0000_0000;
array[26394] <= 16'b0000_0000_0000_0000;
array[26395] <= 16'b0000_0000_0000_0000;
array[26396] <= 16'b0000_0000_0000_0000;
array[26397] <= 16'b0000_0000_0000_0000;
array[26398] <= 16'b0000_0000_0000_0000;
array[26399] <= 16'b0000_0000_0000_0000;
array[26400] <= 16'b0000_0000_0000_0000;
array[26401] <= 16'b0000_0000_0000_0000;
array[26402] <= 16'b0000_0000_0000_0000;
array[26403] <= 16'b0000_0000_0000_0000;
array[26404] <= 16'b0000_0000_0000_0000;
array[26405] <= 16'b0000_0000_0000_0000;
array[26406] <= 16'b0000_0000_0000_0000;
array[26407] <= 16'b0000_0000_0000_0000;
array[26408] <= 16'b0000_0000_0000_0000;
array[26409] <= 16'b0000_0000_0000_0000;
array[26410] <= 16'b0000_0000_0000_0000;
array[26411] <= 16'b0000_0000_0000_0000;
array[26412] <= 16'b0000_0000_0000_0000;
array[26413] <= 16'b0000_0000_0000_0000;
array[26414] <= 16'b0000_0000_0000_0000;
array[26415] <= 16'b0000_0000_0000_0000;
array[26416] <= 16'b0000_0000_0000_0000;
array[26417] <= 16'b0000_0000_0000_0000;
array[26418] <= 16'b0000_0000_0000_0000;
array[26419] <= 16'b0000_0000_0000_0000;
array[26420] <= 16'b0000_0000_0000_0000;
array[26421] <= 16'b0000_0000_0000_0000;
array[26422] <= 16'b0000_0000_0000_0000;
array[26423] <= 16'b0000_0000_0000_0000;
array[26424] <= 16'b0000_0000_0000_0000;
array[26425] <= 16'b0000_0000_0000_0000;
array[26426] <= 16'b0000_0000_0000_0000;
array[26427] <= 16'b0000_0000_0000_0000;
array[26428] <= 16'b0000_0000_0000_0000;
array[26429] <= 16'b0000_0000_0000_0000;
array[26430] <= 16'b0000_0000_0000_0000;
array[26431] <= 16'b0000_0000_0000_0000;
array[26432] <= 16'b0000_0000_0000_0000;
array[26433] <= 16'b0000_0000_0000_0000;
array[26434] <= 16'b0000_0000_0000_0000;
array[26435] <= 16'b0000_0000_0000_0000;
array[26436] <= 16'b0000_0000_0000_0000;
array[26437] <= 16'b0000_0000_0000_0000;
array[26438] <= 16'b0000_0000_0000_0000;
array[26439] <= 16'b0000_0000_0000_0000;
array[26440] <= 16'b0000_0000_0000_0000;
array[26441] <= 16'b0000_0000_0000_0000;
array[26442] <= 16'b0000_0000_0000_0000;
array[26443] <= 16'b0000_0000_0000_0000;
array[26444] <= 16'b0000_0000_0000_0000;
array[26445] <= 16'b0000_0000_0000_0000;
array[26446] <= 16'b0000_0000_0000_0000;
array[26447] <= 16'b0000_0000_0000_0000;
array[26448] <= 16'b0000_0000_0000_0000;
array[26449] <= 16'b0000_0000_0000_0000;
array[26450] <= 16'b0000_0000_0000_0000;
array[26451] <= 16'b0000_0000_0000_0000;
array[26452] <= 16'b0000_0000_0000_0000;
array[26453] <= 16'b0000_0000_0000_0000;
array[26454] <= 16'b0000_0000_0000_0000;
array[26455] <= 16'b0000_0000_0000_0000;
array[26456] <= 16'b0000_0000_0000_0000;
array[26457] <= 16'b0000_0000_0000_0000;
array[26458] <= 16'b0000_0000_0000_0000;
array[26459] <= 16'b0000_0000_0000_0000;
array[26460] <= 16'b0000_0000_0000_0000;
array[26461] <= 16'b0000_0000_0000_0000;
array[26462] <= 16'b0000_0000_0000_0000;
array[26463] <= 16'b0000_0000_0000_0000;
array[26464] <= 16'b0000_0000_0000_0000;
array[26465] <= 16'b0000_0000_0000_0000;
array[26466] <= 16'b0000_0000_0000_0000;
array[26467] <= 16'b0000_0000_0000_0000;
array[26468] <= 16'b0000_0000_0000_0000;
array[26469] <= 16'b0000_0000_0000_0000;
array[26470] <= 16'b0000_0000_0000_0000;
array[26471] <= 16'b0000_0000_0000_0000;
array[26472] <= 16'b0000_0000_0000_0000;
array[26473] <= 16'b0000_0000_0000_0000;
array[26474] <= 16'b0000_0000_0000_0000;
array[26475] <= 16'b0000_0000_0000_0000;
array[26476] <= 16'b0000_0000_0000_0000;
array[26477] <= 16'b0000_0000_0000_0000;
array[26478] <= 16'b0000_0000_0000_0000;
array[26479] <= 16'b0000_0000_0000_0000;
array[26480] <= 16'b0000_0000_0000_0000;
array[26481] <= 16'b0000_0000_0000_0000;
array[26482] <= 16'b0000_0000_0000_0000;
array[26483] <= 16'b0000_0000_0000_0000;
array[26484] <= 16'b0000_0000_0000_0000;
array[26485] <= 16'b0000_0000_0000_0000;
array[26486] <= 16'b0000_0000_0000_0000;
array[26487] <= 16'b0000_0000_0000_0000;
array[26488] <= 16'b0000_0000_0000_0000;
array[26489] <= 16'b0000_0000_0000_0000;
array[26490] <= 16'b0000_0000_0000_0000;
array[26491] <= 16'b0000_0000_0000_0000;
array[26492] <= 16'b0000_0000_0000_0000;
array[26493] <= 16'b0000_0000_0000_0000;
array[26494] <= 16'b0000_0000_0000_0000;
array[26495] <= 16'b0000_0000_0000_0000;
array[26496] <= 16'b0000_0000_0000_0000;
array[26497] <= 16'b0000_0000_0000_0000;
array[26498] <= 16'b0000_0000_0000_0000;
array[26499] <= 16'b0000_0000_0000_0000;
array[26500] <= 16'b0000_0000_0000_0000;
array[26501] <= 16'b0000_0000_0000_0000;
array[26502] <= 16'b0000_0000_0000_0000;
array[26503] <= 16'b0000_0000_0000_0000;
array[26504] <= 16'b0000_0000_0000_0000;
array[26505] <= 16'b0000_0000_0000_0000;
array[26506] <= 16'b0000_0000_0000_0000;
array[26507] <= 16'b0000_0000_0000_0000;
array[26508] <= 16'b0000_0000_0000_0000;
array[26509] <= 16'b0000_0000_0000_0000;
array[26510] <= 16'b0000_0000_0000_0000;
array[26511] <= 16'b0000_0000_0000_0000;
array[26512] <= 16'b0000_0000_0000_0000;
array[26513] <= 16'b0000_0000_0000_0000;
array[26514] <= 16'b0000_0000_0000_0000;
array[26515] <= 16'b0000_0000_0000_0000;
array[26516] <= 16'b0000_0000_0000_0000;
array[26517] <= 16'b0000_0000_0000_0000;
array[26518] <= 16'b0000_0000_0000_0000;
array[26519] <= 16'b0000_0000_0000_0000;
array[26520] <= 16'b0000_0000_0000_0000;
array[26521] <= 16'b0000_0000_0000_0000;
array[26522] <= 16'b0000_0000_0000_0000;
array[26523] <= 16'b0000_0000_0000_0000;
array[26524] <= 16'b0000_0000_0000_0000;
array[26525] <= 16'b0000_0000_0000_0000;
array[26526] <= 16'b0000_0000_0000_0000;
array[26527] <= 16'b0000_0000_0000_0000;
array[26528] <= 16'b0000_0000_0000_0000;
array[26529] <= 16'b0000_0000_0000_0000;
array[26530] <= 16'b0000_0000_0000_0000;
array[26531] <= 16'b0000_0000_0000_0000;
array[26532] <= 16'b0000_0000_0000_0000;
array[26533] <= 16'b0000_0000_0000_0000;
array[26534] <= 16'b0000_0000_0000_0000;
array[26535] <= 16'b0000_0000_0000_0000;
array[26536] <= 16'b0000_0000_0000_0000;
array[26537] <= 16'b0000_0000_0000_0000;
array[26538] <= 16'b0000_0000_0000_0000;
array[26539] <= 16'b0000_0000_0000_0000;
array[26540] <= 16'b0000_0000_0000_0000;
array[26541] <= 16'b0000_0000_0000_0000;
array[26542] <= 16'b0000_0000_0000_0000;
array[26543] <= 16'b0000_0000_0000_0000;
array[26544] <= 16'b0000_0000_0000_0000;
array[26545] <= 16'b0000_0000_0000_0000;
array[26546] <= 16'b0000_0000_0000_0000;
array[26547] <= 16'b0000_0000_0000_0000;
array[26548] <= 16'b0000_0000_0000_0000;
array[26549] <= 16'b0000_0000_0000_0000;
array[26550] <= 16'b0000_0000_0000_0000;
array[26551] <= 16'b0000_0000_0000_0000;
array[26552] <= 16'b0000_0000_0000_0000;
array[26553] <= 16'b0000_0000_0000_0000;
array[26554] <= 16'b0000_0000_0000_0000;
array[26555] <= 16'b0000_0000_0000_0000;
array[26556] <= 16'b0000_0000_0000_0000;
array[26557] <= 16'b0000_0000_0000_0000;
array[26558] <= 16'b0000_0000_0000_0000;
array[26559] <= 16'b0000_0000_0000_0000;
array[26560] <= 16'b0000_0000_0000_0000;
array[26561] <= 16'b0000_0000_0000_0000;
array[26562] <= 16'b0000_0000_0000_0000;
array[26563] <= 16'b0000_0000_0000_0000;
array[26564] <= 16'b0000_0000_0000_0000;
array[26565] <= 16'b0000_0000_0000_0000;
array[26566] <= 16'b0000_0000_0000_0000;
array[26567] <= 16'b0000_0000_0000_0000;
array[26568] <= 16'b0000_0000_0000_0000;
array[26569] <= 16'b0000_0000_0000_0000;
array[26570] <= 16'b0000_0000_0000_0000;
array[26571] <= 16'b0000_0000_0000_0000;
array[26572] <= 16'b0000_0000_0000_0000;
array[26573] <= 16'b0000_0000_0000_0000;
array[26574] <= 16'b0000_0000_0000_0000;
array[26575] <= 16'b0000_0000_0000_0000;
array[26576] <= 16'b0000_0000_0000_0000;
array[26577] <= 16'b0000_0000_0000_0000;
array[26578] <= 16'b0000_0000_0000_0000;
array[26579] <= 16'b0000_0000_0000_0000;
array[26580] <= 16'b0000_0000_0000_0000;
array[26581] <= 16'b0000_0000_0000_0000;
array[26582] <= 16'b0000_0000_0000_0000;
array[26583] <= 16'b0000_0000_0000_0000;
array[26584] <= 16'b0000_0000_0000_0000;
array[26585] <= 16'b0000_0000_0000_0000;
array[26586] <= 16'b0000_0000_0000_0000;
array[26587] <= 16'b0000_0000_0000_0000;
array[26588] <= 16'b0000_0000_0000_0000;
array[26589] <= 16'b0000_0000_0000_0000;
array[26590] <= 16'b0000_0000_0000_0000;
array[26591] <= 16'b0000_0000_0000_0000;
array[26592] <= 16'b0000_0000_0000_0000;
array[26593] <= 16'b0000_0000_0000_0000;
array[26594] <= 16'b0000_0000_0000_0000;
array[26595] <= 16'b0000_0000_0000_0000;
array[26596] <= 16'b0000_0000_0000_0000;
array[26597] <= 16'b0000_0000_0000_0000;
array[26598] <= 16'b0000_0000_0000_0000;
array[26599] <= 16'b0000_0000_0000_0000;
array[26600] <= 16'b0000_0000_0000_0000;
array[26601] <= 16'b0000_0000_0000_0000;
array[26602] <= 16'b0000_0000_0000_0000;
array[26603] <= 16'b0000_0000_0000_0000;
array[26604] <= 16'b0000_0000_0000_0000;
array[26605] <= 16'b0000_0000_0000_0000;
array[26606] <= 16'b0000_0000_0000_0000;
array[26607] <= 16'b0000_0000_0000_0000;
array[26608] <= 16'b0000_0000_0000_0000;
array[26609] <= 16'b0000_0000_0000_0000;
array[26610] <= 16'b0000_0000_0000_0000;
array[26611] <= 16'b0000_0000_0000_0000;
array[26612] <= 16'b0000_0000_0000_0000;
array[26613] <= 16'b0000_0000_0000_0000;
array[26614] <= 16'b0000_0000_0000_0000;
array[26615] <= 16'b0000_0000_0000_0000;
array[26616] <= 16'b0000_0000_0000_0000;
array[26617] <= 16'b0000_0000_0000_0000;
array[26618] <= 16'b0000_0000_0000_0000;
array[26619] <= 16'b0000_0000_0000_0000;
array[26620] <= 16'b0000_0000_0000_0000;
array[26621] <= 16'b0000_0000_0000_0000;
array[26622] <= 16'b0000_0000_0000_0000;
array[26623] <= 16'b0000_0000_0000_0000;
array[26624] <= 16'b0000_0000_0000_0000;
array[26625] <= 16'b0000_0000_0000_0000;
array[26626] <= 16'b0000_0000_0000_0000;
array[26627] <= 16'b0000_0000_0000_0000;
array[26628] <= 16'b0000_0000_0000_0000;
array[26629] <= 16'b0000_0000_0000_0000;
array[26630] <= 16'b0000_0000_0000_0000;
array[26631] <= 16'b0000_0000_0000_0000;
array[26632] <= 16'b0000_0000_0000_0000;
array[26633] <= 16'b0000_0000_0000_0000;
array[26634] <= 16'b0000_0000_0000_0000;
array[26635] <= 16'b0000_0000_0000_0000;
array[26636] <= 16'b0000_0000_0000_0000;
array[26637] <= 16'b0000_0000_0000_0000;
array[26638] <= 16'b0000_0000_0000_0000;
array[26639] <= 16'b0000_0000_0000_0000;
array[26640] <= 16'b0000_0000_0000_0000;
array[26641] <= 16'b0000_0000_0000_0000;
array[26642] <= 16'b0000_0000_0000_0000;
array[26643] <= 16'b0000_0000_0000_0000;
array[26644] <= 16'b0000_0000_0000_0000;
array[26645] <= 16'b0000_0000_0000_0000;
array[26646] <= 16'b0000_0000_0000_0000;
array[26647] <= 16'b0000_0000_0000_0000;
array[26648] <= 16'b0000_0000_0000_0000;
array[26649] <= 16'b0000_0000_0000_0000;
array[26650] <= 16'b0000_0000_0000_0000;
array[26651] <= 16'b0000_0000_0000_0000;
array[26652] <= 16'b0000_0000_0000_0000;
array[26653] <= 16'b0000_0000_0000_0000;
array[26654] <= 16'b0000_0000_0000_0000;
array[26655] <= 16'b0000_0000_0000_0000;
array[26656] <= 16'b0000_0000_0000_0000;
array[26657] <= 16'b0000_0000_0000_0000;
array[26658] <= 16'b0000_0000_0000_0000;
array[26659] <= 16'b0000_0000_0000_0000;
array[26660] <= 16'b0000_0000_0000_0000;
array[26661] <= 16'b0000_0000_0000_0000;
array[26662] <= 16'b0000_0000_0000_0000;
array[26663] <= 16'b0000_0000_0000_0000;
array[26664] <= 16'b0000_0000_0000_0000;
array[26665] <= 16'b0000_0000_0000_0000;
array[26666] <= 16'b0000_0000_0000_0000;
array[26667] <= 16'b0000_0000_0000_0000;
array[26668] <= 16'b0000_0000_0000_0000;
array[26669] <= 16'b0000_0000_0000_0000;
array[26670] <= 16'b0000_0000_0000_0000;
array[26671] <= 16'b0000_0000_0000_0000;
array[26672] <= 16'b0000_0000_0000_0000;
array[26673] <= 16'b0000_0000_0000_0000;
array[26674] <= 16'b0000_0000_0000_0000;
array[26675] <= 16'b0000_0000_0000_0000;
array[26676] <= 16'b0000_0000_0000_0000;
array[26677] <= 16'b0000_0000_0000_0000;
array[26678] <= 16'b0000_0000_0000_0000;
array[26679] <= 16'b0000_0000_0000_0000;
array[26680] <= 16'b0000_0000_0000_0000;
array[26681] <= 16'b0000_0000_0000_0000;
array[26682] <= 16'b0000_0000_0000_0000;
array[26683] <= 16'b0000_0000_0000_0000;
array[26684] <= 16'b0000_0000_0000_0000;
array[26685] <= 16'b0000_0000_0000_0000;
array[26686] <= 16'b0000_0000_0000_0000;
array[26687] <= 16'b0000_0000_0000_0000;
array[26688] <= 16'b0000_0000_0000_0000;
array[26689] <= 16'b0000_0000_0000_0000;
array[26690] <= 16'b0000_0000_0000_0000;
array[26691] <= 16'b0000_0000_0000_0000;
array[26692] <= 16'b0000_0000_0000_0000;
array[26693] <= 16'b0000_0000_0000_0000;
array[26694] <= 16'b0000_0000_0000_0000;
array[26695] <= 16'b0000_0000_0000_0000;
array[26696] <= 16'b0000_0000_0000_0000;
array[26697] <= 16'b0000_0000_0000_0000;
array[26698] <= 16'b0000_0000_0000_0000;
array[26699] <= 16'b0000_0000_0000_0000;
array[26700] <= 16'b0000_0000_0000_0000;
array[26701] <= 16'b0000_0000_0000_0000;
array[26702] <= 16'b0000_0000_0000_0000;
array[26703] <= 16'b0000_0000_0000_0000;
array[26704] <= 16'b0000_0000_0000_0000;
array[26705] <= 16'b0000_0000_0000_0000;
array[26706] <= 16'b0000_0000_0000_0000;
array[26707] <= 16'b0000_0000_0000_0000;
array[26708] <= 16'b0000_0000_0000_0000;
array[26709] <= 16'b0000_0000_0000_0000;
array[26710] <= 16'b0000_0000_0000_0000;
array[26711] <= 16'b0000_0000_0000_0000;
array[26712] <= 16'b0000_0000_0000_0000;
array[26713] <= 16'b0000_0000_0000_0000;
array[26714] <= 16'b0000_0000_0000_0000;
array[26715] <= 16'b0000_0000_0000_0000;
array[26716] <= 16'b0000_0000_0000_0000;
array[26717] <= 16'b0000_0000_0000_0000;
array[26718] <= 16'b0000_0000_0000_0000;
array[26719] <= 16'b0000_0000_0000_0000;
array[26720] <= 16'b0000_0000_0000_0000;
array[26721] <= 16'b0000_0000_0000_0000;
array[26722] <= 16'b0000_0000_0000_0000;
array[26723] <= 16'b0000_0000_0000_0000;
array[26724] <= 16'b0000_0000_0000_0000;
array[26725] <= 16'b0000_0000_0000_0000;
array[26726] <= 16'b0000_0000_0000_0000;
array[26727] <= 16'b0000_0000_0000_0000;
array[26728] <= 16'b0000_0000_0000_0000;
array[26729] <= 16'b0000_0000_0000_0000;
array[26730] <= 16'b0000_0000_0000_0000;
array[26731] <= 16'b0000_0000_0000_0000;
array[26732] <= 16'b0000_0000_0000_0000;
array[26733] <= 16'b0000_0000_0000_0000;
array[26734] <= 16'b0000_0000_0000_0000;
array[26735] <= 16'b0000_0000_0000_0000;
array[26736] <= 16'b0000_0000_0000_0000;
array[26737] <= 16'b0000_0000_0000_0000;
array[26738] <= 16'b0000_0000_0000_0000;
array[26739] <= 16'b0000_0000_0000_0000;
array[26740] <= 16'b0000_0000_0000_0000;
array[26741] <= 16'b0000_0000_0000_0000;
array[26742] <= 16'b0000_0000_0000_0000;
array[26743] <= 16'b0000_0000_0000_0000;
array[26744] <= 16'b0000_0000_0000_0000;
array[26745] <= 16'b0000_0000_0000_0000;
array[26746] <= 16'b0000_0000_0000_0000;
array[26747] <= 16'b0000_0000_0000_0000;
array[26748] <= 16'b0000_0000_0000_0000;
array[26749] <= 16'b0000_0000_0000_0000;
array[26750] <= 16'b0000_0000_0000_0000;
array[26751] <= 16'b0000_0000_0000_0000;
array[26752] <= 16'b0000_0000_0000_0000;
array[26753] <= 16'b0000_0000_0000_0000;
array[26754] <= 16'b0000_0000_0000_0000;
array[26755] <= 16'b0000_0000_0000_0000;
array[26756] <= 16'b0000_0000_0000_0000;
array[26757] <= 16'b0000_0000_0000_0000;
array[26758] <= 16'b0000_0000_0000_0000;
array[26759] <= 16'b0000_0000_0000_0000;
array[26760] <= 16'b0000_0000_0000_0000;
array[26761] <= 16'b0000_0000_0000_0000;
array[26762] <= 16'b0000_0000_0000_0000;
array[26763] <= 16'b0000_0000_0000_0000;
array[26764] <= 16'b0000_0000_0000_0000;
array[26765] <= 16'b0000_0000_0000_0000;
array[26766] <= 16'b0000_0000_0000_0000;
array[26767] <= 16'b0000_0000_0000_0000;
array[26768] <= 16'b0000_0000_0000_0000;
array[26769] <= 16'b0000_0000_0000_0000;
array[26770] <= 16'b0000_0000_0000_0000;
array[26771] <= 16'b0000_0000_0000_0000;
array[26772] <= 16'b0000_0000_0000_0000;
array[26773] <= 16'b0000_0000_0000_0000;
array[26774] <= 16'b0000_0000_0000_0000;
array[26775] <= 16'b0000_0000_0000_0000;
array[26776] <= 16'b0000_0000_0000_0000;
array[26777] <= 16'b0000_0000_0000_0000;
array[26778] <= 16'b0000_0000_0000_0000;
array[26779] <= 16'b0000_0000_0000_0000;
array[26780] <= 16'b0000_0000_0000_0000;
array[26781] <= 16'b0000_0000_0000_0000;
array[26782] <= 16'b0000_0000_0000_0000;
array[26783] <= 16'b0000_0000_0000_0000;
array[26784] <= 16'b0000_0000_0000_0000;
array[26785] <= 16'b0000_0000_0000_0000;
array[26786] <= 16'b0000_0000_0000_0000;
array[26787] <= 16'b0000_0000_0000_0000;
array[26788] <= 16'b0000_0000_0000_0000;
array[26789] <= 16'b0000_0000_0000_0000;
array[26790] <= 16'b0000_0000_0000_0000;
array[26791] <= 16'b0000_0000_0000_0000;
array[26792] <= 16'b0000_0000_0000_0000;
array[26793] <= 16'b0000_0000_0000_0000;
array[26794] <= 16'b0000_0000_0000_0000;
array[26795] <= 16'b0000_0000_0000_0000;
array[26796] <= 16'b0000_0000_0000_0000;
array[26797] <= 16'b0000_0000_0000_0000;
array[26798] <= 16'b0000_0000_0000_0000;
array[26799] <= 16'b0000_0000_0000_0000;
array[26800] <= 16'b0000_0000_0000_0000;
array[26801] <= 16'b0000_0000_0000_0000;
array[26802] <= 16'b0000_0000_0000_0000;
array[26803] <= 16'b0000_0000_0000_0000;
array[26804] <= 16'b0000_0000_0000_0000;
array[26805] <= 16'b0000_0000_0000_0000;
array[26806] <= 16'b0000_0000_0000_0000;
array[26807] <= 16'b0000_0000_0000_0000;
array[26808] <= 16'b0000_0000_0000_0000;
array[26809] <= 16'b0000_0000_0000_0000;
array[26810] <= 16'b0000_0000_0000_0000;
array[26811] <= 16'b0000_0000_0000_0000;
array[26812] <= 16'b0000_0000_0000_0000;
array[26813] <= 16'b0000_0000_0000_0000;
array[26814] <= 16'b0000_0000_0000_0000;
array[26815] <= 16'b0000_0000_0000_0000;
array[26816] <= 16'b0000_0000_0000_0000;
array[26817] <= 16'b0000_0000_0000_0000;
array[26818] <= 16'b0000_0000_0000_0000;
array[26819] <= 16'b0000_0000_0000_0000;
array[26820] <= 16'b0000_0000_0000_0000;
array[26821] <= 16'b0000_0000_0000_0000;
array[26822] <= 16'b0000_0000_0000_0000;
array[26823] <= 16'b0000_0000_0000_0000;
array[26824] <= 16'b0000_0000_0000_0000;
array[26825] <= 16'b0000_0000_0000_0000;
array[26826] <= 16'b0000_0000_0000_0000;
array[26827] <= 16'b0000_0000_0000_0000;
array[26828] <= 16'b0000_0000_0000_0000;
array[26829] <= 16'b0000_0000_0000_0000;
array[26830] <= 16'b0000_0000_0000_0000;
array[26831] <= 16'b0000_0000_0000_0000;
array[26832] <= 16'b0000_0000_0000_0000;
array[26833] <= 16'b0000_0000_0000_0000;
array[26834] <= 16'b0000_0000_0000_0000;
array[26835] <= 16'b0000_0000_0000_0000;
array[26836] <= 16'b0000_0000_0000_0000;
array[26837] <= 16'b0000_0000_0000_0000;
array[26838] <= 16'b0000_0000_0000_0000;
array[26839] <= 16'b0000_0000_0000_0000;
array[26840] <= 16'b0000_0000_0000_0000;
array[26841] <= 16'b0000_0000_0000_0000;
array[26842] <= 16'b0000_0000_0000_0000;
array[26843] <= 16'b0000_0000_0000_0000;
array[26844] <= 16'b0000_0000_0000_0000;
array[26845] <= 16'b0000_0000_0000_0000;
array[26846] <= 16'b0000_0000_0000_0000;
array[26847] <= 16'b0000_0000_0000_0000;
array[26848] <= 16'b0000_0000_0000_0000;
array[26849] <= 16'b0000_0000_0000_0000;
array[26850] <= 16'b0000_0000_0000_0000;
array[26851] <= 16'b0000_0000_0000_0000;
array[26852] <= 16'b0000_0000_0000_0000;
array[26853] <= 16'b0000_0000_0000_0000;
array[26854] <= 16'b0000_0000_0000_0000;
array[26855] <= 16'b0000_0000_0000_0000;
array[26856] <= 16'b0000_0000_0000_0000;
array[26857] <= 16'b0000_0000_0000_0000;
array[26858] <= 16'b0000_0000_0000_0000;
array[26859] <= 16'b0000_0000_0000_0000;
array[26860] <= 16'b0000_0000_0000_0000;
array[26861] <= 16'b0000_0000_0000_0000;
array[26862] <= 16'b0000_0000_0000_0000;
array[26863] <= 16'b0000_0000_0000_0000;
array[26864] <= 16'b0000_0000_0000_0000;
array[26865] <= 16'b0000_0000_0000_0000;
array[26866] <= 16'b0000_0000_0000_0000;
array[26867] <= 16'b0000_0000_0000_0000;
array[26868] <= 16'b0000_0000_0000_0000;
array[26869] <= 16'b0000_0000_0000_0000;
array[26870] <= 16'b0000_0000_0000_0000;
array[26871] <= 16'b0000_0000_0000_0000;
array[26872] <= 16'b0000_0000_0000_0000;
array[26873] <= 16'b0000_0000_0000_0000;
array[26874] <= 16'b0000_0000_0000_0000;
array[26875] <= 16'b0000_0000_0000_0000;
array[26876] <= 16'b0000_0000_0000_0000;
array[26877] <= 16'b0000_0000_0000_0000;
array[26878] <= 16'b0000_0000_0000_0000;
array[26879] <= 16'b0000_0000_0000_0000;
array[26880] <= 16'b0000_0000_0000_0000;
array[26881] <= 16'b0000_0000_0000_0000;
array[26882] <= 16'b0000_0000_0000_0000;
array[26883] <= 16'b0000_0000_0000_0000;
array[26884] <= 16'b0000_0000_0000_0000;
array[26885] <= 16'b0000_0000_0000_0000;
array[26886] <= 16'b0000_0000_0000_0000;
array[26887] <= 16'b0000_0000_0000_0000;
array[26888] <= 16'b0000_0000_0000_0000;
array[26889] <= 16'b0000_0000_0000_0000;
array[26890] <= 16'b0000_0000_0000_0000;
array[26891] <= 16'b0000_0000_0000_0000;
array[26892] <= 16'b0000_0000_0000_0000;
array[26893] <= 16'b0000_0000_0000_0000;
array[26894] <= 16'b0000_0000_0000_0000;
array[26895] <= 16'b0000_0000_0000_0000;
array[26896] <= 16'b0000_0000_0000_0000;
array[26897] <= 16'b0000_0000_0000_0000;
array[26898] <= 16'b0000_0000_0000_0000;
array[26899] <= 16'b0000_0000_0000_0000;
array[26900] <= 16'b0000_0000_0000_0000;
array[26901] <= 16'b0000_0000_0000_0000;
array[26902] <= 16'b0000_0000_0000_0000;
array[26903] <= 16'b0000_0000_0000_0000;
array[26904] <= 16'b0000_0000_0000_0000;
array[26905] <= 16'b0000_0000_0000_0000;
array[26906] <= 16'b0000_0000_0000_0000;
array[26907] <= 16'b0000_0000_0000_0000;
array[26908] <= 16'b0000_0000_0000_0000;
array[26909] <= 16'b0000_0000_0000_0000;
array[26910] <= 16'b0000_0000_0000_0000;
array[26911] <= 16'b0000_0000_0000_0000;
array[26912] <= 16'b0000_0000_0000_0000;
array[26913] <= 16'b0000_0000_0000_0000;
array[26914] <= 16'b0000_0000_0000_0000;
array[26915] <= 16'b0000_0000_0000_0000;
array[26916] <= 16'b0000_0000_0000_0000;
array[26917] <= 16'b0000_0000_0000_0000;
array[26918] <= 16'b0000_0000_0000_0000;
array[26919] <= 16'b0000_0000_0000_0000;
array[26920] <= 16'b0000_0000_0000_0000;
array[26921] <= 16'b0000_0000_0000_0000;
array[26922] <= 16'b0000_0000_0000_0000;
array[26923] <= 16'b0000_0000_0000_0000;
array[26924] <= 16'b0000_0000_0000_0000;
array[26925] <= 16'b0000_0000_0000_0000;
array[26926] <= 16'b0000_0000_0000_0000;
array[26927] <= 16'b0000_0000_0000_0000;
array[26928] <= 16'b0000_0000_0000_0000;
array[26929] <= 16'b0000_0000_0000_0000;
array[26930] <= 16'b0000_0000_0000_0000;
array[26931] <= 16'b0000_0000_0000_0000;
array[26932] <= 16'b0000_0000_0000_0000;
array[26933] <= 16'b0000_0000_0000_0000;
array[26934] <= 16'b0000_0000_0000_0000;
array[26935] <= 16'b0000_0000_0000_0000;
array[26936] <= 16'b0000_0000_0000_0000;
array[26937] <= 16'b0000_0000_0000_0000;
array[26938] <= 16'b0000_0000_0000_0000;
array[26939] <= 16'b0000_0000_0000_0000;
array[26940] <= 16'b0000_0000_0000_0000;
array[26941] <= 16'b0000_0000_0000_0000;
array[26942] <= 16'b0000_0000_0000_0000;
array[26943] <= 16'b0000_0000_0000_0000;
array[26944] <= 16'b0000_0000_0000_0000;
array[26945] <= 16'b0000_0000_0000_0000;
array[26946] <= 16'b0000_0000_0000_0000;
array[26947] <= 16'b0000_0000_0000_0000;
array[26948] <= 16'b0000_0000_0000_0000;
array[26949] <= 16'b0000_0000_0000_0000;
array[26950] <= 16'b0000_0000_0000_0000;
array[26951] <= 16'b0000_0000_0000_0000;
array[26952] <= 16'b0000_0000_0000_0000;
array[26953] <= 16'b0000_0000_0000_0000;
array[26954] <= 16'b0000_0000_0000_0000;
array[26955] <= 16'b0000_0000_0000_0000;
array[26956] <= 16'b0000_0000_0000_0000;
array[26957] <= 16'b0000_0000_0000_0000;
array[26958] <= 16'b0000_0000_0000_0000;
array[26959] <= 16'b0000_0000_0000_0000;
array[26960] <= 16'b0000_0000_0000_0000;
array[26961] <= 16'b0000_0000_0000_0000;
array[26962] <= 16'b0000_0000_0000_0000;
array[26963] <= 16'b0000_0000_0000_0000;
array[26964] <= 16'b0000_0000_0000_0000;
array[26965] <= 16'b0000_0000_0000_0000;
array[26966] <= 16'b0000_0000_0000_0000;
array[26967] <= 16'b0000_0000_0000_0000;
array[26968] <= 16'b0000_0000_0000_0000;
array[26969] <= 16'b0000_0000_0000_0000;
array[26970] <= 16'b0000_0000_0000_0000;
array[26971] <= 16'b0000_0000_0000_0000;
array[26972] <= 16'b0000_0000_0000_0000;
array[26973] <= 16'b0000_0000_0000_0000;
array[26974] <= 16'b0000_0000_0000_0000;
array[26975] <= 16'b0000_0000_0000_0000;
array[26976] <= 16'b0000_0000_0000_0000;
array[26977] <= 16'b0000_0000_0000_0000;
array[26978] <= 16'b0000_0000_0000_0000;
array[26979] <= 16'b0000_0000_0000_0000;
array[26980] <= 16'b0000_0000_0000_0000;
array[26981] <= 16'b0000_0000_0000_0000;
array[26982] <= 16'b0000_0000_0000_0000;
array[26983] <= 16'b0000_0000_0000_0000;
array[26984] <= 16'b0000_0000_0000_0000;
array[26985] <= 16'b0000_0000_0000_0000;
array[26986] <= 16'b0000_0000_0000_0000;
array[26987] <= 16'b0000_0000_0000_0000;
array[26988] <= 16'b0000_0000_0000_0000;
array[26989] <= 16'b0000_0000_0000_0000;
array[26990] <= 16'b0000_0000_0000_0000;
array[26991] <= 16'b0000_0000_0000_0000;
array[26992] <= 16'b0000_0000_0000_0000;
array[26993] <= 16'b0000_0000_0000_0000;
array[26994] <= 16'b0000_0000_0000_0000;
array[26995] <= 16'b0000_0000_0000_0000;
array[26996] <= 16'b0000_0000_0000_0000;
array[26997] <= 16'b0000_0000_0000_0000;
array[26998] <= 16'b0000_0000_0000_0000;
array[26999] <= 16'b0000_0000_0000_0000;
array[27000] <= 16'b0000_0000_0000_0000;
array[27001] <= 16'b0000_0000_0000_0000;
array[27002] <= 16'b0000_0000_0000_0000;
array[27003] <= 16'b0000_0000_0000_0000;
array[27004] <= 16'b0000_0000_0000_0000;
array[27005] <= 16'b0000_0000_0000_0000;
array[27006] <= 16'b0000_0000_0000_0000;
array[27007] <= 16'b0000_0000_0000_0000;
array[27008] <= 16'b0000_0000_0000_0000;
array[27009] <= 16'b0000_0000_0000_0000;
array[27010] <= 16'b0000_0000_0000_0000;
array[27011] <= 16'b0000_0000_0000_0000;
array[27012] <= 16'b0000_0000_0000_0000;
array[27013] <= 16'b0000_0000_0000_0000;
array[27014] <= 16'b0000_0000_0000_0000;
array[27015] <= 16'b0000_0000_0000_0000;
array[27016] <= 16'b0000_0000_0000_0000;
array[27017] <= 16'b0000_0000_0000_0000;
array[27018] <= 16'b0000_0000_0000_0000;
array[27019] <= 16'b0000_0000_0000_0000;
array[27020] <= 16'b0000_0000_0000_0000;
array[27021] <= 16'b0000_0000_0000_0000;
array[27022] <= 16'b0000_0000_0000_0000;
array[27023] <= 16'b0000_0000_0000_0000;
array[27024] <= 16'b0000_0000_0000_0000;
array[27025] <= 16'b0000_0000_0000_0000;
array[27026] <= 16'b0000_0000_0000_0000;
array[27027] <= 16'b0000_0000_0000_0000;
array[27028] <= 16'b0000_0000_0000_0000;
array[27029] <= 16'b0000_0000_0000_0000;
array[27030] <= 16'b0000_0000_0000_0000;
array[27031] <= 16'b0000_0000_0000_0000;
array[27032] <= 16'b0000_0000_0000_0000;
array[27033] <= 16'b0000_0000_0000_0000;
array[27034] <= 16'b0000_0000_0000_0000;
array[27035] <= 16'b0000_0000_0000_0000;
array[27036] <= 16'b0000_0000_0000_0000;
array[27037] <= 16'b0000_0000_0000_0000;
array[27038] <= 16'b0000_0000_0000_0000;
array[27039] <= 16'b0000_0000_0000_0000;
array[27040] <= 16'b0000_0000_0000_0000;
array[27041] <= 16'b0000_0000_0000_0000;
array[27042] <= 16'b0000_0000_0000_0000;
array[27043] <= 16'b0000_0000_0000_0000;
array[27044] <= 16'b0000_0000_0000_0000;
array[27045] <= 16'b0000_0000_0000_0000;
array[27046] <= 16'b0000_0000_0000_0000;
array[27047] <= 16'b0000_0000_0000_0000;
array[27048] <= 16'b0000_0000_0000_0000;
array[27049] <= 16'b0000_0000_0000_0000;
array[27050] <= 16'b0000_0000_0000_0000;
array[27051] <= 16'b0000_0000_0000_0000;
array[27052] <= 16'b0000_0000_0000_0000;
array[27053] <= 16'b0000_0000_0000_0000;
array[27054] <= 16'b0000_0000_0000_0000;
array[27055] <= 16'b0000_0000_0000_0000;
array[27056] <= 16'b0000_0000_0000_0000;
array[27057] <= 16'b0000_0000_0000_0000;
array[27058] <= 16'b0000_0000_0000_0000;
array[27059] <= 16'b0000_0000_0000_0000;
array[27060] <= 16'b0000_0000_0000_0000;
array[27061] <= 16'b0000_0000_0000_0000;
array[27062] <= 16'b0000_0000_0000_0000;
array[27063] <= 16'b0000_0000_0000_0000;
array[27064] <= 16'b0000_0000_0000_0000;
array[27065] <= 16'b0000_0000_0000_0000;
array[27066] <= 16'b0000_0000_0000_0000;
array[27067] <= 16'b0000_0000_0000_0000;
array[27068] <= 16'b0000_0000_0000_0000;
array[27069] <= 16'b0000_0000_0000_0000;
array[27070] <= 16'b0000_0000_0000_0000;
array[27071] <= 16'b0000_0000_0000_0000;
array[27072] <= 16'b0000_0000_0000_0000;
array[27073] <= 16'b0000_0000_0000_0000;
array[27074] <= 16'b0000_0000_0000_0000;
array[27075] <= 16'b0000_0000_0000_0000;
array[27076] <= 16'b0000_0000_0000_0000;
array[27077] <= 16'b0000_0000_0000_0000;
array[27078] <= 16'b0000_0000_0000_0000;
array[27079] <= 16'b0000_0000_0000_0000;
array[27080] <= 16'b0000_0000_0000_0000;
array[27081] <= 16'b0000_0000_0000_0000;
array[27082] <= 16'b0000_0000_0000_0000;
array[27083] <= 16'b0000_0000_0000_0000;
array[27084] <= 16'b0000_0000_0000_0000;
array[27085] <= 16'b0000_0000_0000_0000;
array[27086] <= 16'b0000_0000_0000_0000;
array[27087] <= 16'b0000_0000_0000_0000;
array[27088] <= 16'b0000_0000_0000_0000;
array[27089] <= 16'b0000_0000_0000_0000;
array[27090] <= 16'b0000_0000_0000_0000;
array[27091] <= 16'b0000_0000_0000_0000;
array[27092] <= 16'b0000_0000_0000_0000;
array[27093] <= 16'b0000_0000_0000_0000;
array[27094] <= 16'b0000_0000_0000_0000;
array[27095] <= 16'b0000_0000_0000_0000;
array[27096] <= 16'b0000_0000_0000_0000;
array[27097] <= 16'b0000_0000_0000_0000;
array[27098] <= 16'b0000_0000_0000_0000;
array[27099] <= 16'b0000_0000_0000_0000;
array[27100] <= 16'b0000_0000_0000_0000;
array[27101] <= 16'b0000_0000_0000_0000;
array[27102] <= 16'b0000_0000_0000_0000;
array[27103] <= 16'b0000_0000_0000_0000;
array[27104] <= 16'b0000_0000_0000_0000;
array[27105] <= 16'b0000_0000_0000_0000;
array[27106] <= 16'b0000_0000_0000_0000;
array[27107] <= 16'b0000_0000_0000_0000;
array[27108] <= 16'b0000_0000_0000_0000;
array[27109] <= 16'b0000_0000_0000_0000;
array[27110] <= 16'b0000_0000_0000_0000;
array[27111] <= 16'b0000_0000_0000_0000;
array[27112] <= 16'b0000_0000_0000_0000;
array[27113] <= 16'b0000_0000_0000_0000;
array[27114] <= 16'b0000_0000_0000_0000;
array[27115] <= 16'b0000_0000_0000_0000;
array[27116] <= 16'b0000_0000_0000_0000;
array[27117] <= 16'b0000_0000_0000_0000;
array[27118] <= 16'b0000_0000_0000_0000;
array[27119] <= 16'b0000_0000_0000_0000;
array[27120] <= 16'b0000_0000_0000_0000;
array[27121] <= 16'b0000_0000_0000_0000;
array[27122] <= 16'b0000_0000_0000_0000;
array[27123] <= 16'b0000_0000_0000_0000;
array[27124] <= 16'b0000_0000_0000_0000;
array[27125] <= 16'b0000_0000_0000_0000;
array[27126] <= 16'b0000_0000_0000_0000;
array[27127] <= 16'b0000_0000_0000_0000;
array[27128] <= 16'b0000_0000_0000_0000;
array[27129] <= 16'b0000_0000_0000_0000;
array[27130] <= 16'b0000_0000_0000_0000;
array[27131] <= 16'b0000_0000_0000_0000;
array[27132] <= 16'b0000_0000_0000_0000;
array[27133] <= 16'b0000_0000_0000_0000;
array[27134] <= 16'b0000_0000_0000_0000;
array[27135] <= 16'b0000_0000_0000_0000;
array[27136] <= 16'b0000_0000_0000_0000;
array[27137] <= 16'b0000_0000_0000_0000;
array[27138] <= 16'b0000_0000_0000_0000;
array[27139] <= 16'b0000_0000_0000_0000;
array[27140] <= 16'b0000_0000_0000_0000;
array[27141] <= 16'b0000_0000_0000_0000;
array[27142] <= 16'b0000_0000_0000_0000;
array[27143] <= 16'b0000_0000_0000_0000;
array[27144] <= 16'b0000_0000_0000_0000;
array[27145] <= 16'b0000_0000_0000_0000;
array[27146] <= 16'b0000_0000_0000_0000;
array[27147] <= 16'b0000_0000_0000_0000;
array[27148] <= 16'b0000_0000_0000_0000;
array[27149] <= 16'b0000_0000_0000_0000;
array[27150] <= 16'b0000_0000_0000_0000;
array[27151] <= 16'b0000_0000_0000_0000;
array[27152] <= 16'b0000_0000_0000_0000;
array[27153] <= 16'b0000_0000_0000_0000;
array[27154] <= 16'b0000_0000_0000_0000;
array[27155] <= 16'b0000_0000_0000_0000;
array[27156] <= 16'b0000_0000_0000_0000;
array[27157] <= 16'b0000_0000_0000_0000;
array[27158] <= 16'b0000_0000_0000_0000;
array[27159] <= 16'b0000_0000_0000_0000;
array[27160] <= 16'b0000_0000_0000_0000;
array[27161] <= 16'b0000_0000_0000_0000;
array[27162] <= 16'b0000_0000_0000_0000;
array[27163] <= 16'b0000_0000_0000_0000;
array[27164] <= 16'b0000_0000_0000_0000;
array[27165] <= 16'b0000_0000_0000_0000;
array[27166] <= 16'b0000_0000_0000_0000;
array[27167] <= 16'b0000_0000_0000_0000;
array[27168] <= 16'b0000_0000_0000_0000;
array[27169] <= 16'b0000_0000_0000_0000;
array[27170] <= 16'b0000_0000_0000_0000;
array[27171] <= 16'b0000_0000_0000_0000;
array[27172] <= 16'b0000_0000_0000_0000;
array[27173] <= 16'b0000_0000_0000_0000;
array[27174] <= 16'b0000_0000_0000_0000;
array[27175] <= 16'b0000_0000_0000_0000;
array[27176] <= 16'b0000_0000_0000_0000;
array[27177] <= 16'b0000_0000_0000_0000;
array[27178] <= 16'b0000_0000_0000_0000;
array[27179] <= 16'b0000_0000_0000_0000;
array[27180] <= 16'b0000_0000_0000_0000;
array[27181] <= 16'b0000_0000_0000_0000;
array[27182] <= 16'b0000_0000_0000_0000;
array[27183] <= 16'b0000_0000_0000_0000;
array[27184] <= 16'b0000_0000_0000_0000;
array[27185] <= 16'b0000_0000_0000_0000;
array[27186] <= 16'b0000_0000_0000_0000;
array[27187] <= 16'b0000_0000_0000_0000;
array[27188] <= 16'b0000_0000_0000_0000;
array[27189] <= 16'b0000_0000_0000_0000;
array[27190] <= 16'b0000_0000_0000_0000;
array[27191] <= 16'b0000_0000_0000_0000;
array[27192] <= 16'b0000_0000_0000_0000;
array[27193] <= 16'b0000_0000_0000_0000;
array[27194] <= 16'b0000_0000_0000_0000;
array[27195] <= 16'b0000_0000_0000_0000;
array[27196] <= 16'b0000_0000_0000_0000;
array[27197] <= 16'b0000_0000_0000_0000;
array[27198] <= 16'b0000_0000_0000_0000;
array[27199] <= 16'b0000_0000_0000_0000;
array[27200] <= 16'b0000_0000_0000_0000;
array[27201] <= 16'b0000_0000_0000_0000;
array[27202] <= 16'b0000_0000_0000_0000;
array[27203] <= 16'b0000_0000_0000_0000;
array[27204] <= 16'b0000_0000_0000_0000;
array[27205] <= 16'b0000_0000_0000_0000;
array[27206] <= 16'b0000_0000_0000_0000;
array[27207] <= 16'b0000_0000_0000_0000;
array[27208] <= 16'b0000_0000_0000_0000;
array[27209] <= 16'b0000_0000_0000_0000;
array[27210] <= 16'b0000_0000_0000_0000;
array[27211] <= 16'b0000_0000_0000_0000;
array[27212] <= 16'b0000_0000_0000_0000;
array[27213] <= 16'b0000_0000_0000_0000;
array[27214] <= 16'b0000_0000_0000_0000;
array[27215] <= 16'b0000_0000_0000_0000;
array[27216] <= 16'b0000_0000_0000_0000;
array[27217] <= 16'b0000_0000_0000_0000;
array[27218] <= 16'b0000_0000_0000_0000;
array[27219] <= 16'b0000_0000_0000_0000;
array[27220] <= 16'b0000_0000_0000_0000;
array[27221] <= 16'b0000_0000_0000_0000;
array[27222] <= 16'b0000_0000_0000_0000;
array[27223] <= 16'b0000_0000_0000_0000;
array[27224] <= 16'b0000_0000_0000_0000;
array[27225] <= 16'b0000_0000_0000_0000;
array[27226] <= 16'b0000_0000_0000_0000;
array[27227] <= 16'b0000_0000_0000_0000;
array[27228] <= 16'b0000_0000_0000_0000;
array[27229] <= 16'b0000_0000_0000_0000;
array[27230] <= 16'b0000_0000_0000_0000;
array[27231] <= 16'b0000_0000_0000_0000;
array[27232] <= 16'b0000_0000_0000_0000;
array[27233] <= 16'b0000_0000_0000_0000;
array[27234] <= 16'b0000_0000_0000_0000;
array[27235] <= 16'b0000_0000_0000_0000;
array[27236] <= 16'b0000_0000_0000_0000;
array[27237] <= 16'b0000_0000_0000_0000;
array[27238] <= 16'b0000_0000_0000_0000;
array[27239] <= 16'b0000_0000_0000_0000;
array[27240] <= 16'b0000_0000_0000_0000;
array[27241] <= 16'b0000_0000_0000_0000;
array[27242] <= 16'b0000_0000_0000_0000;
array[27243] <= 16'b0000_0000_0000_0000;
array[27244] <= 16'b0000_0000_0000_0000;
array[27245] <= 16'b0000_0000_0000_0000;
array[27246] <= 16'b0000_0000_0000_0000;
array[27247] <= 16'b0000_0000_0000_0000;
array[27248] <= 16'b0000_0000_0000_0000;
array[27249] <= 16'b0000_0000_0000_0000;
array[27250] <= 16'b0000_0000_0000_0000;
array[27251] <= 16'b0000_0000_0000_0000;
array[27252] <= 16'b0000_0000_0000_0000;
array[27253] <= 16'b0000_0000_0000_0000;
array[27254] <= 16'b0000_0000_0000_0000;
array[27255] <= 16'b0000_0000_0000_0000;
array[27256] <= 16'b0000_0000_0000_0000;
array[27257] <= 16'b0000_0000_0000_0000;
array[27258] <= 16'b0000_0000_0000_0000;
array[27259] <= 16'b0000_0000_0000_0000;
array[27260] <= 16'b0000_0000_0000_0000;
array[27261] <= 16'b0000_0000_0000_0000;
array[27262] <= 16'b0000_0000_0000_0000;
array[27263] <= 16'b0000_0000_0000_0000;
array[27264] <= 16'b0000_0000_0000_0000;
array[27265] <= 16'b0000_0000_0000_0000;
array[27266] <= 16'b0000_0000_0000_0000;
array[27267] <= 16'b0000_0000_0000_0000;
array[27268] <= 16'b0000_0000_0000_0000;
array[27269] <= 16'b0000_0000_0000_0000;
array[27270] <= 16'b0000_0000_0000_0000;
array[27271] <= 16'b0000_0000_0000_0000;
array[27272] <= 16'b0000_0000_0000_0000;
array[27273] <= 16'b0000_0000_0000_0000;
array[27274] <= 16'b0000_0000_0000_0000;
array[27275] <= 16'b0000_0000_0000_0000;
array[27276] <= 16'b0000_0000_0000_0000;
array[27277] <= 16'b0000_0000_0000_0000;
array[27278] <= 16'b0000_0000_0000_0000;
array[27279] <= 16'b0000_0000_0000_0000;
array[27280] <= 16'b0000_0000_0000_0000;
array[27281] <= 16'b0000_0000_0000_0000;
array[27282] <= 16'b0000_0000_0000_0000;
array[27283] <= 16'b0000_0000_0000_0000;
array[27284] <= 16'b0000_0000_0000_0000;
array[27285] <= 16'b0000_0000_0000_0000;
array[27286] <= 16'b0000_0000_0000_0000;
array[27287] <= 16'b0000_0000_0000_0000;
array[27288] <= 16'b0000_0000_0000_0000;
array[27289] <= 16'b0000_0000_0000_0000;
array[27290] <= 16'b0000_0000_0000_0000;
array[27291] <= 16'b0000_0000_0000_0000;
array[27292] <= 16'b0000_0000_0000_0000;
array[27293] <= 16'b0000_0000_0000_0000;
array[27294] <= 16'b0000_0000_0000_0000;
array[27295] <= 16'b0000_0000_0000_0000;
array[27296] <= 16'b0000_0000_0000_0000;
array[27297] <= 16'b0000_0000_0000_0000;
array[27298] <= 16'b0000_0000_0000_0000;
array[27299] <= 16'b0000_0000_0000_0000;
array[27300] <= 16'b0000_0000_0000_0000;
array[27301] <= 16'b0000_0000_0000_0000;
array[27302] <= 16'b0000_0000_0000_0000;
array[27303] <= 16'b0000_0000_0000_0000;
array[27304] <= 16'b0000_0000_0000_0000;
array[27305] <= 16'b0000_0000_0000_0000;
array[27306] <= 16'b0000_0000_0000_0000;
array[27307] <= 16'b0000_0000_0000_0000;
array[27308] <= 16'b0000_0000_0000_0000;
array[27309] <= 16'b0000_0000_0000_0000;
array[27310] <= 16'b0000_0000_0000_0000;
array[27311] <= 16'b0000_0000_0000_0000;
array[27312] <= 16'b0000_0000_0000_0000;
array[27313] <= 16'b0000_0000_0000_0000;
array[27314] <= 16'b0000_0000_0000_0000;
array[27315] <= 16'b0000_0000_0000_0000;
array[27316] <= 16'b0000_0000_0000_0000;
array[27317] <= 16'b0000_0000_0000_0000;
array[27318] <= 16'b0000_0000_0000_0000;
array[27319] <= 16'b0000_0000_0000_0000;
array[27320] <= 16'b0000_0000_0000_0000;
array[27321] <= 16'b0000_0000_0000_0000;
array[27322] <= 16'b0000_0000_0000_0000;
array[27323] <= 16'b0000_0000_0000_0000;
array[27324] <= 16'b0000_0000_0000_0000;
array[27325] <= 16'b0000_0000_0000_0000;
array[27326] <= 16'b0000_0000_0000_0000;
array[27327] <= 16'b0000_0000_0000_0000;
array[27328] <= 16'b0000_0000_0000_0000;
array[27329] <= 16'b0000_0000_0000_0000;
array[27330] <= 16'b0000_0000_0000_0000;
array[27331] <= 16'b0000_0000_0000_0000;
array[27332] <= 16'b0000_0000_0000_0000;
array[27333] <= 16'b0000_0000_0000_0000;
array[27334] <= 16'b0000_0000_0000_0000;
array[27335] <= 16'b0000_0000_0000_0000;
array[27336] <= 16'b0000_0000_0000_0000;
array[27337] <= 16'b0000_0000_0000_0000;
array[27338] <= 16'b0000_0000_0000_0000;
array[27339] <= 16'b0000_0000_0000_0000;
array[27340] <= 16'b0000_0000_0000_0000;
array[27341] <= 16'b0000_0000_0000_0000;
array[27342] <= 16'b0000_0000_0000_0000;
array[27343] <= 16'b0000_0000_0000_0000;
array[27344] <= 16'b0000_0000_0000_0000;
array[27345] <= 16'b0000_0000_0000_0000;
array[27346] <= 16'b0000_0000_0000_0000;
array[27347] <= 16'b0000_0000_0000_0000;
array[27348] <= 16'b0000_0000_0000_0000;
array[27349] <= 16'b0000_0000_0000_0000;
array[27350] <= 16'b0000_0000_0000_0000;
array[27351] <= 16'b0000_0000_0000_0000;
array[27352] <= 16'b0000_0000_0000_0000;
array[27353] <= 16'b0000_0000_0000_0000;
array[27354] <= 16'b0000_0000_0000_0000;
array[27355] <= 16'b0000_0000_0000_0000;
array[27356] <= 16'b0000_0000_0000_0000;
array[27357] <= 16'b0000_0000_0000_0000;
array[27358] <= 16'b0000_0000_0000_0000;
array[27359] <= 16'b0000_0000_0000_0000;
array[27360] <= 16'b0000_0000_0000_0000;
array[27361] <= 16'b0000_0000_0000_0000;
array[27362] <= 16'b0000_0000_0000_0000;
array[27363] <= 16'b0000_0000_0000_0000;
array[27364] <= 16'b0000_0000_0000_0000;
array[27365] <= 16'b0000_0000_0000_0000;
array[27366] <= 16'b0000_0000_0000_0000;
array[27367] <= 16'b0000_0000_0000_0000;
array[27368] <= 16'b0000_0000_0000_0000;
array[27369] <= 16'b0000_0000_0000_0000;
array[27370] <= 16'b0000_0000_0000_0000;
array[27371] <= 16'b0000_0000_0000_0000;
array[27372] <= 16'b0000_0000_0000_0000;
array[27373] <= 16'b0000_0000_0000_0000;
array[27374] <= 16'b0000_0000_0000_0000;
array[27375] <= 16'b0000_0000_0000_0000;
array[27376] <= 16'b0000_0000_0000_0000;
array[27377] <= 16'b0000_0000_0000_0000;
array[27378] <= 16'b0000_0000_0000_0000;
array[27379] <= 16'b0000_0000_0000_0000;
array[27380] <= 16'b0000_0000_0000_0000;
array[27381] <= 16'b0000_0000_0000_0000;
array[27382] <= 16'b0000_0000_0000_0000;
array[27383] <= 16'b0000_0000_0000_0000;
array[27384] <= 16'b0000_0000_0000_0000;
array[27385] <= 16'b0000_0000_0000_0000;
array[27386] <= 16'b0000_0000_0000_0000;
array[27387] <= 16'b0000_0000_0000_0000;
array[27388] <= 16'b0000_0000_0000_0000;
array[27389] <= 16'b0000_0000_0000_0000;
array[27390] <= 16'b0000_0000_0000_0000;
array[27391] <= 16'b0000_0000_0000_0000;
array[27392] <= 16'b0000_0000_0000_0000;
array[27393] <= 16'b0000_0000_0000_0000;
array[27394] <= 16'b0000_0000_0000_0000;
array[27395] <= 16'b0000_0000_0000_0000;
array[27396] <= 16'b0000_0000_0000_0000;
array[27397] <= 16'b0000_0000_0000_0000;
array[27398] <= 16'b0000_0000_0000_0000;
array[27399] <= 16'b0000_0000_0000_0000;
array[27400] <= 16'b0000_0000_0000_0000;
array[27401] <= 16'b0000_0000_0000_0000;
array[27402] <= 16'b0000_0000_0000_0000;
array[27403] <= 16'b0000_0000_0000_0000;
array[27404] <= 16'b0000_0000_0000_0000;
array[27405] <= 16'b0000_0000_0000_0000;
array[27406] <= 16'b0000_0000_0000_0000;
array[27407] <= 16'b0000_0000_0000_0000;
array[27408] <= 16'b0000_0000_0000_0000;
array[27409] <= 16'b0000_0000_0000_0000;
array[27410] <= 16'b0000_0000_0000_0000;
array[27411] <= 16'b0000_0000_0000_0000;
array[27412] <= 16'b0000_0000_0000_0000;
array[27413] <= 16'b0000_0000_0000_0000;
array[27414] <= 16'b0000_0000_0000_0000;
array[27415] <= 16'b0000_0000_0000_0000;
array[27416] <= 16'b0000_0000_0000_0000;
array[27417] <= 16'b0000_0000_0000_0000;
array[27418] <= 16'b0000_0000_0000_0000;
array[27419] <= 16'b0000_0000_0000_0000;
array[27420] <= 16'b0000_0000_0000_0000;
array[27421] <= 16'b0000_0000_0000_0000;
array[27422] <= 16'b0000_0000_0000_0000;
array[27423] <= 16'b0000_0000_0000_0000;
array[27424] <= 16'b0000_0000_0000_0000;
array[27425] <= 16'b0000_0000_0000_0000;
array[27426] <= 16'b0000_0000_0000_0000;
array[27427] <= 16'b0000_0000_0000_0000;
array[27428] <= 16'b0000_0000_0000_0000;
array[27429] <= 16'b0000_0000_0000_0000;
array[27430] <= 16'b0000_0000_0000_0000;
array[27431] <= 16'b0000_0000_0000_0000;
array[27432] <= 16'b0000_0000_0000_0000;
array[27433] <= 16'b0000_0000_0000_0000;
array[27434] <= 16'b0000_0000_0000_0000;
array[27435] <= 16'b0000_0000_0000_0000;
array[27436] <= 16'b0000_0000_0000_0000;
array[27437] <= 16'b0000_0000_0000_0000;
array[27438] <= 16'b0000_0000_0000_0000;
array[27439] <= 16'b0000_0000_0000_0000;
array[27440] <= 16'b0000_0000_0000_0000;
array[27441] <= 16'b0000_0000_0000_0000;
array[27442] <= 16'b0000_0000_0000_0000;
array[27443] <= 16'b0000_0000_0000_0000;
array[27444] <= 16'b0000_0000_0000_0000;
array[27445] <= 16'b0000_0000_0000_0000;
array[27446] <= 16'b0000_0000_0000_0000;
array[27447] <= 16'b0000_0000_0000_0000;
array[27448] <= 16'b0000_0000_0000_0000;
array[27449] <= 16'b0000_0000_0000_0000;
array[27450] <= 16'b0000_0000_0000_0000;
array[27451] <= 16'b0000_0000_0000_0000;
array[27452] <= 16'b0000_0000_0000_0000;
array[27453] <= 16'b0000_0000_0000_0000;
array[27454] <= 16'b0000_0000_0000_0000;
array[27455] <= 16'b0000_0000_0000_0000;
array[27456] <= 16'b0000_0000_0000_0000;
array[27457] <= 16'b0000_0000_0000_0000;
array[27458] <= 16'b0000_0000_0000_0000;
array[27459] <= 16'b0000_0000_0000_0000;
array[27460] <= 16'b0000_0000_0000_0000;
array[27461] <= 16'b0000_0000_0000_0000;
array[27462] <= 16'b0000_0000_0000_0000;
array[27463] <= 16'b0000_0000_0000_0000;
array[27464] <= 16'b0000_0000_0000_0000;
array[27465] <= 16'b0000_0000_0000_0000;
array[27466] <= 16'b0000_0000_0000_0000;
array[27467] <= 16'b0000_0000_0000_0000;
array[27468] <= 16'b0000_0000_0000_0000;
array[27469] <= 16'b0000_0000_0000_0000;
array[27470] <= 16'b0000_0000_0000_0000;
array[27471] <= 16'b0000_0000_0000_0000;
array[27472] <= 16'b0000_0000_0000_0000;
array[27473] <= 16'b0000_0000_0000_0000;
array[27474] <= 16'b0000_0000_0000_0000;
array[27475] <= 16'b0000_0000_0000_0000;
array[27476] <= 16'b0000_0000_0000_0000;
array[27477] <= 16'b0000_0000_0000_0000;
array[27478] <= 16'b0000_0000_0000_0000;
array[27479] <= 16'b0000_0000_0000_0000;
array[27480] <= 16'b0000_0000_0000_0000;
array[27481] <= 16'b0000_0000_0000_0000;
array[27482] <= 16'b0000_0000_0000_0000;
array[27483] <= 16'b0000_0000_0000_0000;
array[27484] <= 16'b0000_0000_0000_0000;
array[27485] <= 16'b0000_0000_0000_0000;
array[27486] <= 16'b0000_0000_0000_0000;
array[27487] <= 16'b0000_0000_0000_0000;
array[27488] <= 16'b0000_0000_0000_0000;
array[27489] <= 16'b0000_0000_0000_0000;
array[27490] <= 16'b0000_0000_0000_0000;
array[27491] <= 16'b0000_0000_0000_0000;
array[27492] <= 16'b0000_0000_0000_0000;
array[27493] <= 16'b0000_0000_0000_0000;
array[27494] <= 16'b0000_0000_0000_0000;
array[27495] <= 16'b0000_0000_0000_0000;
array[27496] <= 16'b0000_0000_0000_0000;
array[27497] <= 16'b0000_0000_0000_0000;
array[27498] <= 16'b0000_0000_0000_0000;
array[27499] <= 16'b0000_0000_0000_0000;
array[27500] <= 16'b0000_0000_0000_0000;
array[27501] <= 16'b0000_0000_0000_0000;
array[27502] <= 16'b0000_0000_0000_0000;
array[27503] <= 16'b0000_0000_0000_0000;
array[27504] <= 16'b0000_0000_0000_0000;
array[27505] <= 16'b0000_0000_0000_0000;
array[27506] <= 16'b0000_0000_0000_0000;
array[27507] <= 16'b0000_0000_0000_0000;
array[27508] <= 16'b0000_0000_0000_0000;
array[27509] <= 16'b0000_0000_0000_0000;
array[27510] <= 16'b0000_0000_0000_0000;
array[27511] <= 16'b0000_0000_0000_0000;
array[27512] <= 16'b0000_0000_0000_0000;
array[27513] <= 16'b0000_0000_0000_0000;
array[27514] <= 16'b0000_0000_0000_0000;
array[27515] <= 16'b0000_0000_0000_0000;
array[27516] <= 16'b0000_0000_0000_0000;
array[27517] <= 16'b0000_0000_0000_0000;
array[27518] <= 16'b0000_0000_0000_0000;
array[27519] <= 16'b0000_0000_0000_0000;
array[27520] <= 16'b0000_0000_0000_0000;
array[27521] <= 16'b0000_0000_0000_0000;
array[27522] <= 16'b0000_0000_0000_0000;
array[27523] <= 16'b0000_0000_0000_0000;
array[27524] <= 16'b0000_0000_0000_0000;
array[27525] <= 16'b0000_0000_0000_0000;
array[27526] <= 16'b0000_0000_0000_0000;
array[27527] <= 16'b0000_0000_0000_0000;
array[27528] <= 16'b0000_0000_0000_0000;
array[27529] <= 16'b0000_0000_0000_0000;
array[27530] <= 16'b0000_0000_0000_0000;
array[27531] <= 16'b0000_0000_0000_0000;
array[27532] <= 16'b0000_0000_0000_0000;
array[27533] <= 16'b0000_0000_0000_0000;
array[27534] <= 16'b0000_0000_0000_0000;
array[27535] <= 16'b0000_0000_0000_0000;
array[27536] <= 16'b0000_0000_0000_0000;
array[27537] <= 16'b0000_0000_0000_0000;
array[27538] <= 16'b0000_0000_0000_0000;
array[27539] <= 16'b0000_0000_0000_0000;
array[27540] <= 16'b0000_0000_0000_0000;
array[27541] <= 16'b0000_0000_0000_0000;
array[27542] <= 16'b0000_0000_0000_0000;
array[27543] <= 16'b0000_0000_0000_0000;
array[27544] <= 16'b0000_0000_0000_0000;
array[27545] <= 16'b0000_0000_0000_0000;
array[27546] <= 16'b0000_0000_0000_0000;
array[27547] <= 16'b0000_0000_0000_0000;
array[27548] <= 16'b0000_0000_0000_0000;
array[27549] <= 16'b0000_0000_0000_0000;
array[27550] <= 16'b0000_0000_0000_0000;
array[27551] <= 16'b0000_0000_0000_0000;
array[27552] <= 16'b0000_0000_0000_0000;
array[27553] <= 16'b0000_0000_0000_0000;
array[27554] <= 16'b0000_0000_0000_0000;
array[27555] <= 16'b0000_0000_0000_0000;
array[27556] <= 16'b0000_0000_0000_0000;
array[27557] <= 16'b0000_0000_0000_0000;
array[27558] <= 16'b0000_0000_0000_0000;
array[27559] <= 16'b0000_0000_0000_0000;
array[27560] <= 16'b0000_0000_0000_0000;
array[27561] <= 16'b0000_0000_0000_0000;
array[27562] <= 16'b0000_0000_0000_0000;
array[27563] <= 16'b0000_0000_0000_0000;
array[27564] <= 16'b0000_0000_0000_0000;
array[27565] <= 16'b0000_0000_0000_0000;
array[27566] <= 16'b0000_0000_0000_0000;
array[27567] <= 16'b0000_0000_0000_0000;
array[27568] <= 16'b0000_0000_0000_0000;
array[27569] <= 16'b0000_0000_0000_0000;
array[27570] <= 16'b0000_0000_0000_0000;
array[27571] <= 16'b0000_0000_0000_0000;
array[27572] <= 16'b0000_0000_0000_0000;
array[27573] <= 16'b0000_0000_0000_0000;
array[27574] <= 16'b0000_0000_0000_0000;
array[27575] <= 16'b0000_0000_0000_0000;
array[27576] <= 16'b0000_0000_0000_0000;
array[27577] <= 16'b0000_0000_0000_0000;
array[27578] <= 16'b0000_0000_0000_0000;
array[27579] <= 16'b0000_0000_0000_0000;
array[27580] <= 16'b0000_0000_0000_0000;
array[27581] <= 16'b0000_0000_0000_0000;
array[27582] <= 16'b0000_0000_0000_0000;
array[27583] <= 16'b0000_0000_0000_0000;
array[27584] <= 16'b0000_0000_0000_0000;
array[27585] <= 16'b0000_0000_0000_0000;
array[27586] <= 16'b0000_0000_0000_0000;
array[27587] <= 16'b0000_0000_0000_0000;
array[27588] <= 16'b0000_0000_0000_0000;
array[27589] <= 16'b0000_0000_0000_0000;
array[27590] <= 16'b0000_0000_0000_0000;
array[27591] <= 16'b0000_0000_0000_0000;
array[27592] <= 16'b0000_0000_0000_0000;
array[27593] <= 16'b0000_0000_0000_0000;
array[27594] <= 16'b0000_0000_0000_0000;
array[27595] <= 16'b0000_0000_0000_0000;
array[27596] <= 16'b0000_0000_0000_0000;
array[27597] <= 16'b0000_0000_0000_0000;
array[27598] <= 16'b0000_0000_0000_0000;
array[27599] <= 16'b0000_0000_0000_0000;
array[27600] <= 16'b0000_0000_0000_0000;
array[27601] <= 16'b0000_0000_0000_0000;
array[27602] <= 16'b0000_0000_0000_0000;
array[27603] <= 16'b0000_0000_0000_0000;
array[27604] <= 16'b0000_0000_0000_0000;
array[27605] <= 16'b0000_0000_0000_0000;
array[27606] <= 16'b0000_0000_0000_0000;
array[27607] <= 16'b0000_0000_0000_0000;
array[27608] <= 16'b0000_0000_0000_0000;
array[27609] <= 16'b0000_0000_0000_0000;
array[27610] <= 16'b0000_0000_0000_0000;
array[27611] <= 16'b0000_0000_0000_0000;
array[27612] <= 16'b0000_0000_0000_0000;
array[27613] <= 16'b0000_0000_0000_0000;
array[27614] <= 16'b0000_0000_0000_0000;
array[27615] <= 16'b0000_0000_0000_0000;
array[27616] <= 16'b0000_0000_0000_0000;
array[27617] <= 16'b0000_0000_0000_0000;
array[27618] <= 16'b0000_0000_0000_0000;
array[27619] <= 16'b0000_0000_0000_0000;
array[27620] <= 16'b0000_0000_0000_0000;
array[27621] <= 16'b0000_0000_0000_0000;
array[27622] <= 16'b0000_0000_0000_0000;
array[27623] <= 16'b0000_0000_0000_0000;
array[27624] <= 16'b0000_0000_0000_0000;
array[27625] <= 16'b0000_0000_0000_0000;
array[27626] <= 16'b0000_0000_0000_0000;
array[27627] <= 16'b0000_0000_0000_0000;
array[27628] <= 16'b0000_0000_0000_0000;
array[27629] <= 16'b0000_0000_0000_0000;
array[27630] <= 16'b0000_0000_0000_0000;
array[27631] <= 16'b0000_0000_0000_0000;
array[27632] <= 16'b0000_0000_0000_0000;
array[27633] <= 16'b0000_0000_0000_0000;
array[27634] <= 16'b0000_0000_0000_0000;
array[27635] <= 16'b0000_0000_0000_0000;
array[27636] <= 16'b0000_0000_0000_0000;
array[27637] <= 16'b0000_0000_0000_0000;
array[27638] <= 16'b0000_0000_0000_0000;
array[27639] <= 16'b0000_0000_0000_0000;
array[27640] <= 16'b0000_0000_0000_0000;
array[27641] <= 16'b0000_0000_0000_0000;
array[27642] <= 16'b0000_0000_0000_0000;
array[27643] <= 16'b0000_0000_0000_0000;
array[27644] <= 16'b0000_0000_0000_0000;
array[27645] <= 16'b0000_0000_0000_0000;
array[27646] <= 16'b0000_0000_0000_0000;
array[27647] <= 16'b0000_0000_0000_0000;
array[27648] <= 16'b0000_0000_0000_0000;
array[27649] <= 16'b0000_0000_0000_0000;
array[27650] <= 16'b0000_0000_0000_0000;
array[27651] <= 16'b0000_0000_0000_0000;
array[27652] <= 16'b0000_0000_0000_0000;
array[27653] <= 16'b0000_0000_0000_0000;
array[27654] <= 16'b0000_0000_0000_0000;
array[27655] <= 16'b0000_0000_0000_0000;
array[27656] <= 16'b0000_0000_0000_0000;
array[27657] <= 16'b0000_0000_0000_0000;
array[27658] <= 16'b0000_0000_0000_0000;
array[27659] <= 16'b0000_0000_0000_0000;
array[27660] <= 16'b0000_0000_0000_0000;
array[27661] <= 16'b0000_0000_0000_0000;
array[27662] <= 16'b0000_0000_0000_0000;
array[27663] <= 16'b0000_0000_0000_0000;
array[27664] <= 16'b0000_0000_0000_0000;
array[27665] <= 16'b0000_0000_0000_0000;
array[27666] <= 16'b0000_0000_0000_0000;
array[27667] <= 16'b0000_0000_0000_0000;
array[27668] <= 16'b0000_0000_0000_0000;
array[27669] <= 16'b0000_0000_0000_0000;
array[27670] <= 16'b0000_0000_0000_0000;
array[27671] <= 16'b0000_0000_0000_0000;
array[27672] <= 16'b0000_0000_0000_0000;
array[27673] <= 16'b0000_0000_0000_0000;
array[27674] <= 16'b0000_0000_0000_0000;
array[27675] <= 16'b0000_0000_0000_0000;
array[27676] <= 16'b0000_0000_0000_0000;
array[27677] <= 16'b0000_0000_0000_0000;
array[27678] <= 16'b0000_0000_0000_0000;
array[27679] <= 16'b0000_0000_0000_0000;
array[27680] <= 16'b0000_0000_0000_0000;
array[27681] <= 16'b0000_0000_0000_0000;
array[27682] <= 16'b0000_0000_0000_0000;
array[27683] <= 16'b0000_0000_0000_0000;
array[27684] <= 16'b0000_0000_0000_0000;
array[27685] <= 16'b0000_0000_0000_0000;
array[27686] <= 16'b0000_0000_0000_0000;
array[27687] <= 16'b0000_0000_0000_0000;
array[27688] <= 16'b0000_0000_0000_0000;
array[27689] <= 16'b0000_0000_0000_0000;
array[27690] <= 16'b0000_0000_0000_0000;
array[27691] <= 16'b0000_0000_0000_0000;
array[27692] <= 16'b0000_0000_0000_0000;
array[27693] <= 16'b0000_0000_0000_0000;
array[27694] <= 16'b0000_0000_0000_0000;
array[27695] <= 16'b0000_0000_0000_0000;
array[27696] <= 16'b0000_0000_0000_0000;
array[27697] <= 16'b0000_0000_0000_0000;
array[27698] <= 16'b0000_0000_0000_0000;
array[27699] <= 16'b0000_0000_0000_0000;
array[27700] <= 16'b0000_0000_0000_0000;
array[27701] <= 16'b0000_0000_0000_0000;
array[27702] <= 16'b0000_0000_0000_0000;
array[27703] <= 16'b0000_0000_0000_0000;
array[27704] <= 16'b0000_0000_0000_0000;
array[27705] <= 16'b0000_0000_0000_0000;
array[27706] <= 16'b0000_0000_0000_0000;
array[27707] <= 16'b0000_0000_0000_0000;
array[27708] <= 16'b0000_0000_0000_0000;
array[27709] <= 16'b0000_0000_0000_0000;
array[27710] <= 16'b0000_0000_0000_0000;
array[27711] <= 16'b0000_0000_0000_0000;
array[27712] <= 16'b0000_0000_0000_0000;
array[27713] <= 16'b0000_0000_0000_0000;
array[27714] <= 16'b0000_0000_0000_0000;
array[27715] <= 16'b0000_0000_0000_0000;
array[27716] <= 16'b0000_0000_0000_0000;
array[27717] <= 16'b0000_0000_0000_0000;
array[27718] <= 16'b0000_0000_0000_0000;
array[27719] <= 16'b0000_0000_0000_0000;
array[27720] <= 16'b0000_0000_0000_0000;
array[27721] <= 16'b0000_0000_0000_0000;
array[27722] <= 16'b0000_0000_0000_0000;
array[27723] <= 16'b0000_0000_0000_0000;
array[27724] <= 16'b0000_0000_0000_0000;
array[27725] <= 16'b0000_0000_0000_0000;
array[27726] <= 16'b0000_0000_0000_0000;
array[27727] <= 16'b0000_0000_0000_0000;
array[27728] <= 16'b0000_0000_0000_0000;
array[27729] <= 16'b0000_0000_0000_0000;
array[27730] <= 16'b0000_0000_0000_0000;
array[27731] <= 16'b0000_0000_0000_0000;
array[27732] <= 16'b0000_0000_0000_0000;
array[27733] <= 16'b0000_0000_0000_0000;
array[27734] <= 16'b0000_0000_0000_0000;
array[27735] <= 16'b0000_0000_0000_0000;
array[27736] <= 16'b0000_0000_0000_0000;
array[27737] <= 16'b0000_0000_0000_0000;
array[27738] <= 16'b0000_0000_0000_0000;
array[27739] <= 16'b0000_0000_0000_0000;
array[27740] <= 16'b0000_0000_0000_0000;
array[27741] <= 16'b0000_0000_0000_0000;
array[27742] <= 16'b0000_0000_0000_0000;
array[27743] <= 16'b0000_0000_0000_0000;
array[27744] <= 16'b0000_0000_0000_0000;
array[27745] <= 16'b0000_0000_0000_0000;
array[27746] <= 16'b0000_0000_0000_0000;
array[27747] <= 16'b0000_0000_0000_0000;
array[27748] <= 16'b0000_0000_0000_0000;
array[27749] <= 16'b0000_0000_0000_0000;
array[27750] <= 16'b0000_0000_0000_0000;
array[27751] <= 16'b0000_0000_0000_0000;
array[27752] <= 16'b0000_0000_0000_0000;
array[27753] <= 16'b0000_0000_0000_0000;
array[27754] <= 16'b0000_0000_0000_0000;
array[27755] <= 16'b0000_0000_0000_0000;
array[27756] <= 16'b0000_0000_0000_0000;
array[27757] <= 16'b0000_0000_0000_0000;
array[27758] <= 16'b0000_0000_0000_0000;
array[27759] <= 16'b0000_0000_0000_0000;
array[27760] <= 16'b0000_0000_0000_0000;
array[27761] <= 16'b0000_0000_0000_0000;
array[27762] <= 16'b0000_0000_0000_0000;
array[27763] <= 16'b0000_0000_0000_0000;
array[27764] <= 16'b0000_0000_0000_0000;
array[27765] <= 16'b0000_0000_0000_0000;
array[27766] <= 16'b0000_0000_0000_0000;
array[27767] <= 16'b0000_0000_0000_0000;
array[27768] <= 16'b0000_0000_0000_0000;
array[27769] <= 16'b0000_0000_0000_0000;
array[27770] <= 16'b0000_0000_0000_0000;
array[27771] <= 16'b0000_0000_0000_0000;
array[27772] <= 16'b0000_0000_0000_0000;
array[27773] <= 16'b0000_0000_0000_0000;
array[27774] <= 16'b0000_0000_0000_0000;
array[27775] <= 16'b0000_0000_0000_0000;
array[27776] <= 16'b0000_0000_0000_0000;
array[27777] <= 16'b0000_0000_0000_0000;
array[27778] <= 16'b0000_0000_0000_0000;
array[27779] <= 16'b0000_0000_0000_0000;
array[27780] <= 16'b0000_0000_0000_0000;
array[27781] <= 16'b0000_0000_0000_0000;
array[27782] <= 16'b0000_0000_0000_0000;
array[27783] <= 16'b0000_0000_0000_0000;
array[27784] <= 16'b0000_0000_0000_0000;
array[27785] <= 16'b0000_0000_0000_0000;
array[27786] <= 16'b0000_0000_0000_0000;
array[27787] <= 16'b0000_0000_0000_0000;
array[27788] <= 16'b0000_0000_0000_0000;
array[27789] <= 16'b0000_0000_0000_0000;
array[27790] <= 16'b0000_0000_0000_0000;
array[27791] <= 16'b0000_0000_0000_0000;
array[27792] <= 16'b0000_0000_0000_0000;
array[27793] <= 16'b0000_0000_0000_0000;
array[27794] <= 16'b0000_0000_0000_0000;
array[27795] <= 16'b0000_0000_0000_0000;
array[27796] <= 16'b0000_0000_0000_0000;
array[27797] <= 16'b0000_0000_0000_0000;
array[27798] <= 16'b0000_0000_0000_0000;
array[27799] <= 16'b0000_0000_0000_0000;
array[27800] <= 16'b0000_0000_0000_0000;
array[27801] <= 16'b0000_0000_0000_0000;
array[27802] <= 16'b0000_0000_0000_0000;
array[27803] <= 16'b0000_0000_0000_0000;
array[27804] <= 16'b0000_0000_0000_0000;
array[27805] <= 16'b0000_0000_0000_0000;
array[27806] <= 16'b0000_0000_0000_0000;
array[27807] <= 16'b0000_0000_0000_0000;
array[27808] <= 16'b0000_0000_0000_0000;
array[27809] <= 16'b0000_0000_0000_0000;
array[27810] <= 16'b0000_0000_0000_0000;
array[27811] <= 16'b0000_0000_0000_0000;
array[27812] <= 16'b0000_0000_0000_0000;
array[27813] <= 16'b0000_0000_0000_0000;
array[27814] <= 16'b0000_0000_0000_0000;
array[27815] <= 16'b0000_0000_0000_0000;
array[27816] <= 16'b0000_0000_0000_0000;
array[27817] <= 16'b0000_0000_0000_0000;
array[27818] <= 16'b0000_0000_0000_0000;
array[27819] <= 16'b0000_0000_0000_0000;
array[27820] <= 16'b0000_0000_0000_0000;
array[27821] <= 16'b0000_0000_0000_0000;
array[27822] <= 16'b0000_0000_0000_0000;
array[27823] <= 16'b0000_0000_0000_0000;
array[27824] <= 16'b0000_0000_0000_0000;
array[27825] <= 16'b0000_0000_0000_0000;
array[27826] <= 16'b0000_0000_0000_0000;
array[27827] <= 16'b0000_0000_0000_0000;
array[27828] <= 16'b0000_0000_0000_0000;
array[27829] <= 16'b0000_0000_0000_0000;
array[27830] <= 16'b0000_0000_0000_0000;
array[27831] <= 16'b0000_0000_0000_0000;
array[27832] <= 16'b0000_0000_0000_0000;
array[27833] <= 16'b0000_0000_0000_0000;
array[27834] <= 16'b0000_0000_0000_0000;
array[27835] <= 16'b0000_0000_0000_0000;
array[27836] <= 16'b0000_0000_0000_0000;
array[27837] <= 16'b0000_0000_0000_0000;
array[27838] <= 16'b0000_0000_0000_0000;
array[27839] <= 16'b0000_0000_0000_0000;
array[27840] <= 16'b0000_0000_0000_0000;
array[27841] <= 16'b0000_0000_0000_0000;
array[27842] <= 16'b0000_0000_0000_0000;
array[27843] <= 16'b0000_0000_0000_0000;
array[27844] <= 16'b0000_0000_0000_0000;
array[27845] <= 16'b0000_0000_0000_0000;
array[27846] <= 16'b0000_0000_0000_0000;
array[27847] <= 16'b0000_0000_0000_0000;
array[27848] <= 16'b0000_0000_0000_0000;
array[27849] <= 16'b0000_0000_0000_0000;
array[27850] <= 16'b0000_0000_0000_0000;
array[27851] <= 16'b0000_0000_0000_0000;
array[27852] <= 16'b0000_0000_0000_0000;
array[27853] <= 16'b0000_0000_0000_0000;
array[27854] <= 16'b0000_0000_0000_0000;
array[27855] <= 16'b0000_0000_0000_0000;
array[27856] <= 16'b0000_0000_0000_0000;
array[27857] <= 16'b0000_0000_0000_0000;
array[27858] <= 16'b0000_0000_0000_0000;
array[27859] <= 16'b0000_0000_0000_0000;
array[27860] <= 16'b0000_0000_0000_0000;
array[27861] <= 16'b0000_0000_0000_0000;
array[27862] <= 16'b0000_0000_0000_0000;
array[27863] <= 16'b0000_0000_0000_0000;
array[27864] <= 16'b0000_0000_0000_0000;
array[27865] <= 16'b0000_0000_0000_0000;
array[27866] <= 16'b0000_0000_0000_0000;
array[27867] <= 16'b0000_0000_0000_0000;
array[27868] <= 16'b0000_0000_0000_0000;
array[27869] <= 16'b0000_0000_0000_0000;
array[27870] <= 16'b0000_0000_0000_0000;
array[27871] <= 16'b0000_0000_0000_0000;
array[27872] <= 16'b0000_0000_0000_0000;
array[27873] <= 16'b0000_0000_0000_0000;
array[27874] <= 16'b0000_0000_0000_0000;
array[27875] <= 16'b0000_0000_0000_0000;
array[27876] <= 16'b0000_0000_0000_0000;
array[27877] <= 16'b0000_0000_0000_0000;
array[27878] <= 16'b0000_0000_0000_0000;
array[27879] <= 16'b0000_0000_0000_0000;
array[27880] <= 16'b0000_0000_0000_0000;
array[27881] <= 16'b0000_0000_0000_0000;
array[27882] <= 16'b0000_0000_0000_0000;
array[27883] <= 16'b0000_0000_0000_0000;
array[27884] <= 16'b0000_0000_0000_0000;
array[27885] <= 16'b0000_0000_0000_0000;
array[27886] <= 16'b0000_0000_0000_0000;
array[27887] <= 16'b0000_0000_0000_0000;
array[27888] <= 16'b0000_0000_0000_0000;
array[27889] <= 16'b0000_0000_0000_0000;
array[27890] <= 16'b0000_0000_0000_0000;
array[27891] <= 16'b0000_0000_0000_0000;
array[27892] <= 16'b0000_0000_0000_0000;
array[27893] <= 16'b0000_0000_0000_0000;
array[27894] <= 16'b0000_0000_0000_0000;
array[27895] <= 16'b0000_0000_0000_0000;
array[27896] <= 16'b0000_0000_0000_0000;
array[27897] <= 16'b0000_0000_0000_0000;
array[27898] <= 16'b0000_0000_0000_0000;
array[27899] <= 16'b0000_0000_0000_0000;
array[27900] <= 16'b0000_0000_0000_0000;
array[27901] <= 16'b0000_0000_0000_0000;
array[27902] <= 16'b0000_0000_0000_0000;
array[27903] <= 16'b0000_0000_0000_0000;
array[27904] <= 16'b0000_0000_0000_0000;
array[27905] <= 16'b0000_0000_0000_0000;
array[27906] <= 16'b0000_0000_0000_0000;
array[27907] <= 16'b0000_0000_0000_0000;
array[27908] <= 16'b0000_0000_0000_0000;
array[27909] <= 16'b0000_0000_0000_0000;
array[27910] <= 16'b0000_0000_0000_0000;
array[27911] <= 16'b0000_0000_0000_0000;
array[27912] <= 16'b0000_0000_0000_0000;
array[27913] <= 16'b0000_0000_0000_0000;
array[27914] <= 16'b0000_0000_0000_0000;
array[27915] <= 16'b0000_0000_0000_0000;
array[27916] <= 16'b0000_0000_0000_0000;
array[27917] <= 16'b0000_0000_0000_0000;
array[27918] <= 16'b0000_0000_0000_0000;
array[27919] <= 16'b0000_0000_0000_0000;
array[27920] <= 16'b0000_0000_0000_0000;
array[27921] <= 16'b0000_0000_0000_0000;
array[27922] <= 16'b0000_0000_0000_0000;
array[27923] <= 16'b0000_0000_0000_0000;
array[27924] <= 16'b0000_0000_0000_0000;
array[27925] <= 16'b0000_0000_0000_0000;
array[27926] <= 16'b0000_0000_0000_0000;
array[27927] <= 16'b0000_0000_0000_0000;
array[27928] <= 16'b0000_0000_0000_0000;
array[27929] <= 16'b0000_0000_0000_0000;
array[27930] <= 16'b0000_0000_0000_0000;
array[27931] <= 16'b0000_0000_0000_0000;
array[27932] <= 16'b0000_0000_0000_0000;
array[27933] <= 16'b0000_0000_0000_0000;
array[27934] <= 16'b0000_0000_0000_0000;
array[27935] <= 16'b0000_0000_0000_0000;
array[27936] <= 16'b0000_0000_0000_0000;
array[27937] <= 16'b0000_0000_0000_0000;
array[27938] <= 16'b0000_0000_0000_0000;
array[27939] <= 16'b0000_0000_0000_0000;
array[27940] <= 16'b0000_0000_0000_0000;
array[27941] <= 16'b0000_0000_0000_0000;
array[27942] <= 16'b0000_0000_0000_0000;
array[27943] <= 16'b0000_0000_0000_0000;
array[27944] <= 16'b0000_0000_0000_0000;
array[27945] <= 16'b0000_0000_0000_0000;
array[27946] <= 16'b0000_0000_0000_0000;
array[27947] <= 16'b0000_0000_0000_0000;
array[27948] <= 16'b0000_0000_0000_0000;
array[27949] <= 16'b0000_0000_0000_0000;
array[27950] <= 16'b0000_0000_0000_0000;
array[27951] <= 16'b0000_0000_0000_0000;
array[27952] <= 16'b0000_0000_0000_0000;
array[27953] <= 16'b0000_0000_0000_0000;
array[27954] <= 16'b0000_0000_0000_0000;
array[27955] <= 16'b0000_0000_0000_0000;
array[27956] <= 16'b0000_0000_0000_0000;
array[27957] <= 16'b0000_0000_0000_0000;
array[27958] <= 16'b0000_0000_0000_0000;
array[27959] <= 16'b0000_0000_0000_0000;
array[27960] <= 16'b0000_0000_0000_0000;
array[27961] <= 16'b0000_0000_0000_0000;
array[27962] <= 16'b0000_0000_0000_0000;
array[27963] <= 16'b0000_0000_0000_0000;
array[27964] <= 16'b0000_0000_0000_0000;
array[27965] <= 16'b0000_0000_0000_0000;
array[27966] <= 16'b0000_0000_0000_0000;
array[27967] <= 16'b0000_0000_0000_0000;
array[27968] <= 16'b0000_0000_0000_0000;
array[27969] <= 16'b0000_0000_0000_0000;
array[27970] <= 16'b0000_0000_0000_0000;
array[27971] <= 16'b0000_0000_0000_0000;
array[27972] <= 16'b0000_0000_0000_0000;
array[27973] <= 16'b0000_0000_0000_0000;
array[27974] <= 16'b0000_0000_0000_0000;
array[27975] <= 16'b0000_0000_0000_0000;
array[27976] <= 16'b0000_0000_0000_0000;
array[27977] <= 16'b0000_0000_0000_0000;
array[27978] <= 16'b0000_0000_0000_0000;
array[27979] <= 16'b0000_0000_0000_0000;
array[27980] <= 16'b0000_0000_0000_0000;
array[27981] <= 16'b0000_0000_0000_0000;
array[27982] <= 16'b0000_0000_0000_0000;
array[27983] <= 16'b0000_0000_0000_0000;
array[27984] <= 16'b0000_0000_0000_0000;
array[27985] <= 16'b0000_0000_0000_0000;
array[27986] <= 16'b0000_0000_0000_0000;
array[27987] <= 16'b0000_0000_0000_0000;
array[27988] <= 16'b0000_0000_0000_0000;
array[27989] <= 16'b0000_0000_0000_0000;
array[27990] <= 16'b0000_0000_0000_0000;
array[27991] <= 16'b0000_0000_0000_0000;
array[27992] <= 16'b0000_0000_0000_0000;
array[27993] <= 16'b0000_0000_0000_0000;
array[27994] <= 16'b0000_0000_0000_0000;
array[27995] <= 16'b0000_0000_0000_0000;
array[27996] <= 16'b0000_0000_0000_0000;
array[27997] <= 16'b0000_0000_0000_0000;
array[27998] <= 16'b0000_0000_0000_0000;
array[27999] <= 16'b0000_0000_0000_0000;
array[28000] <= 16'b0000_0000_0000_0000;
array[28001] <= 16'b0000_0000_0000_0000;
array[28002] <= 16'b0000_0000_0000_0000;
array[28003] <= 16'b0000_0000_0000_0000;
array[28004] <= 16'b0000_0000_0000_0000;
array[28005] <= 16'b0000_0000_0000_0000;
array[28006] <= 16'b0000_0000_0000_0000;
array[28007] <= 16'b0000_0000_0000_0000;
array[28008] <= 16'b0000_0000_0000_0000;
array[28009] <= 16'b0000_0000_0000_0000;
array[28010] <= 16'b0000_0000_0000_0000;
array[28011] <= 16'b0000_0000_0000_0000;
array[28012] <= 16'b0000_0000_0000_0000;
array[28013] <= 16'b0000_0000_0000_0000;
array[28014] <= 16'b0000_0000_0000_0000;
array[28015] <= 16'b0000_0000_0000_0000;
array[28016] <= 16'b0000_0000_0000_0000;
array[28017] <= 16'b0000_0000_0000_0000;
array[28018] <= 16'b0000_0000_0000_0000;
array[28019] <= 16'b0000_0000_0000_0000;
array[28020] <= 16'b0000_0000_0000_0000;
array[28021] <= 16'b0000_0000_0000_0000;
array[28022] <= 16'b0000_0000_0000_0000;
array[28023] <= 16'b0000_0000_0000_0000;
array[28024] <= 16'b0000_0000_0000_0000;
array[28025] <= 16'b0000_0000_0000_0000;
array[28026] <= 16'b0000_0000_0000_0000;
array[28027] <= 16'b0000_0000_0000_0000;
array[28028] <= 16'b0000_0000_0000_0000;
array[28029] <= 16'b0000_0000_0000_0000;
array[28030] <= 16'b0000_0000_0000_0000;
array[28031] <= 16'b0000_0000_0000_0000;
array[28032] <= 16'b0000_0000_0000_0000;
array[28033] <= 16'b0000_0000_0000_0000;
array[28034] <= 16'b0000_0000_0000_0000;
array[28035] <= 16'b0000_0000_0000_0000;
array[28036] <= 16'b0000_0000_0000_0000;
array[28037] <= 16'b0000_0000_0000_0000;
array[28038] <= 16'b0000_0000_0000_0000;
array[28039] <= 16'b0000_0000_0000_0000;
array[28040] <= 16'b0000_0000_0000_0000;
array[28041] <= 16'b0000_0000_0000_0000;
array[28042] <= 16'b0000_0000_0000_0000;
array[28043] <= 16'b0000_0000_0000_0000;
array[28044] <= 16'b0000_0000_0000_0000;
array[28045] <= 16'b0000_0000_0000_0000;
array[28046] <= 16'b0000_0000_0000_0000;
array[28047] <= 16'b0000_0000_0000_0000;
array[28048] <= 16'b0000_0000_0000_0000;
array[28049] <= 16'b0000_0000_0000_0000;
array[28050] <= 16'b0000_0000_0000_0000;
array[28051] <= 16'b0000_0000_0000_0000;
array[28052] <= 16'b0000_0000_0000_0000;
array[28053] <= 16'b0000_0000_0000_0000;
array[28054] <= 16'b0000_0000_0000_0000;
array[28055] <= 16'b0000_0000_0000_0000;
array[28056] <= 16'b0000_0000_0000_0000;
array[28057] <= 16'b0000_0000_0000_0000;
array[28058] <= 16'b0000_0000_0000_0000;
array[28059] <= 16'b0000_0000_0000_0000;
array[28060] <= 16'b0000_0000_0000_0000;
array[28061] <= 16'b0000_0000_0000_0000;
array[28062] <= 16'b0000_0000_0000_0000;
array[28063] <= 16'b0000_0000_0000_0000;
array[28064] <= 16'b0000_0000_0000_0000;
array[28065] <= 16'b0000_0000_0000_0000;
array[28066] <= 16'b0000_0000_0000_0000;
array[28067] <= 16'b0000_0000_0000_0000;
array[28068] <= 16'b0000_0000_0000_0000;
array[28069] <= 16'b0000_0000_0000_0000;
array[28070] <= 16'b0000_0000_0000_0000;
array[28071] <= 16'b0000_0000_0000_0000;
array[28072] <= 16'b0000_0000_0000_0000;
array[28073] <= 16'b0000_0000_0000_0000;
array[28074] <= 16'b0000_0000_0000_0000;
array[28075] <= 16'b0000_0000_0000_0000;
array[28076] <= 16'b0000_0000_0000_0000;
array[28077] <= 16'b0000_0000_0000_0000;
array[28078] <= 16'b0000_0000_0000_0000;
array[28079] <= 16'b0000_0000_0000_0000;
array[28080] <= 16'b0000_0000_0000_0000;
array[28081] <= 16'b0000_0000_0000_0000;
array[28082] <= 16'b0000_0000_0000_0000;
array[28083] <= 16'b0000_0000_0000_0000;
array[28084] <= 16'b0000_0000_0000_0000;
array[28085] <= 16'b0000_0000_0000_0000;
array[28086] <= 16'b0000_0000_0000_0000;
array[28087] <= 16'b0000_0000_0000_0000;
array[28088] <= 16'b0000_0000_0000_0000;
array[28089] <= 16'b0000_0000_0000_0000;
array[28090] <= 16'b0000_0000_0000_0000;
array[28091] <= 16'b0000_0000_0000_0000;
array[28092] <= 16'b0000_0000_0000_0000;
array[28093] <= 16'b0000_0000_0000_0000;
array[28094] <= 16'b0000_0000_0000_0000;
array[28095] <= 16'b0000_0000_0000_0000;
array[28096] <= 16'b0000_0000_0000_0000;
array[28097] <= 16'b0000_0000_0000_0000;
array[28098] <= 16'b0000_0000_0000_0000;
array[28099] <= 16'b0000_0000_0000_0000;
array[28100] <= 16'b0000_0000_0000_0000;
array[28101] <= 16'b0000_0000_0000_0000;
array[28102] <= 16'b0000_0000_0000_0000;
array[28103] <= 16'b0000_0000_0000_0000;
array[28104] <= 16'b0000_0000_0000_0000;
array[28105] <= 16'b0000_0000_0000_0000;
array[28106] <= 16'b0000_0000_0000_0000;
array[28107] <= 16'b0000_0000_0000_0000;
array[28108] <= 16'b0000_0000_0000_0000;
array[28109] <= 16'b0000_0000_0000_0000;
array[28110] <= 16'b0000_0000_0000_0000;
array[28111] <= 16'b0000_0000_0000_0000;
array[28112] <= 16'b0000_0000_0000_0000;
array[28113] <= 16'b0000_0000_0000_0000;
array[28114] <= 16'b0000_0000_0000_0000;
array[28115] <= 16'b0000_0000_0000_0000;
array[28116] <= 16'b0000_0000_0000_0000;
array[28117] <= 16'b0000_0000_0000_0000;
array[28118] <= 16'b0000_0000_0000_0000;
array[28119] <= 16'b0000_0000_0000_0000;
array[28120] <= 16'b0000_0000_0000_0000;
array[28121] <= 16'b0000_0000_0000_0000;
array[28122] <= 16'b0000_0000_0000_0000;
array[28123] <= 16'b0000_0000_0000_0000;
array[28124] <= 16'b0000_0000_0000_0000;
array[28125] <= 16'b0000_0000_0000_0000;
array[28126] <= 16'b0000_0000_0000_0000;
array[28127] <= 16'b0000_0000_0000_0000;
array[28128] <= 16'b0000_0000_0000_0000;
array[28129] <= 16'b0000_0000_0000_0000;
array[28130] <= 16'b0000_0000_0000_0000;
array[28131] <= 16'b0000_0000_0000_0000;
array[28132] <= 16'b0000_0000_0000_0000;
array[28133] <= 16'b0000_0000_0000_0000;
array[28134] <= 16'b0000_0000_0000_0000;
array[28135] <= 16'b0000_0000_0000_0000;
array[28136] <= 16'b0000_0000_0000_0000;
array[28137] <= 16'b0000_0000_0000_0000;
array[28138] <= 16'b0000_0000_0000_0000;
array[28139] <= 16'b0000_0000_0000_0000;
array[28140] <= 16'b0000_0000_0000_0000;
array[28141] <= 16'b0000_0000_0000_0000;
array[28142] <= 16'b0000_0000_0000_0000;
array[28143] <= 16'b0000_0000_0000_0000;
array[28144] <= 16'b0000_0000_0000_0000;
array[28145] <= 16'b0000_0000_0000_0000;
array[28146] <= 16'b0000_0000_0000_0000;
array[28147] <= 16'b0000_0000_0000_0000;
array[28148] <= 16'b0000_0000_0000_0000;
array[28149] <= 16'b0000_0000_0000_0000;
array[28150] <= 16'b0000_0000_0000_0000;
array[28151] <= 16'b0000_0000_0000_0000;
array[28152] <= 16'b0000_0000_0000_0000;
array[28153] <= 16'b0000_0000_0000_0000;
array[28154] <= 16'b0000_0000_0000_0000;
array[28155] <= 16'b0000_0000_0000_0000;
array[28156] <= 16'b0000_0000_0000_0000;
array[28157] <= 16'b0000_0000_0000_0000;
array[28158] <= 16'b0000_0000_0000_0000;
array[28159] <= 16'b0000_0000_0000_0000;
array[28160] <= 16'b0000_0000_0000_0000;
array[28161] <= 16'b0000_0000_0000_0000;
array[28162] <= 16'b0000_0000_0000_0000;
array[28163] <= 16'b0000_0000_0000_0000;
array[28164] <= 16'b0000_0000_0000_0000;
array[28165] <= 16'b0000_0000_0000_0000;
array[28166] <= 16'b0000_0000_0000_0000;
array[28167] <= 16'b0000_0000_0000_0000;
array[28168] <= 16'b0000_0000_0000_0000;
array[28169] <= 16'b0000_0000_0000_0000;
array[28170] <= 16'b0000_0000_0000_0000;
array[28171] <= 16'b0000_0000_0000_0000;
array[28172] <= 16'b0000_0000_0000_0000;
array[28173] <= 16'b0000_0000_0000_0000;
array[28174] <= 16'b0000_0000_0000_0000;
array[28175] <= 16'b0000_0000_0000_0000;
array[28176] <= 16'b0000_0000_0000_0000;
array[28177] <= 16'b0000_0000_0000_0000;
array[28178] <= 16'b0000_0000_0000_0000;
array[28179] <= 16'b0000_0000_0000_0000;
array[28180] <= 16'b0000_0000_0000_0000;
array[28181] <= 16'b0000_0000_0000_0000;
array[28182] <= 16'b0000_0000_0000_0000;
array[28183] <= 16'b0000_0000_0000_0000;
array[28184] <= 16'b0000_0000_0000_0000;
array[28185] <= 16'b0000_0000_0000_0000;
array[28186] <= 16'b0000_0000_0000_0000;
array[28187] <= 16'b0000_0000_0000_0000;
array[28188] <= 16'b0000_0000_0000_0000;
array[28189] <= 16'b0000_0000_0000_0000;
array[28190] <= 16'b0000_0000_0000_0000;
array[28191] <= 16'b0000_0000_0000_0000;
array[28192] <= 16'b0000_0000_0000_0000;
array[28193] <= 16'b0000_0000_0000_0000;
array[28194] <= 16'b0000_0000_0000_0000;
array[28195] <= 16'b0000_0000_0000_0000;
array[28196] <= 16'b0000_0000_0000_0000;
array[28197] <= 16'b0000_0000_0000_0000;
array[28198] <= 16'b0000_0000_0000_0000;
array[28199] <= 16'b0000_0000_0000_0000;
array[28200] <= 16'b0000_0000_0000_0000;
array[28201] <= 16'b0000_0000_0000_0000;
array[28202] <= 16'b0000_0000_0000_0000;
array[28203] <= 16'b0000_0000_0000_0000;
array[28204] <= 16'b0000_0000_0000_0000;
array[28205] <= 16'b0000_0000_0000_0000;
array[28206] <= 16'b0000_0000_0000_0000;
array[28207] <= 16'b0000_0000_0000_0000;
array[28208] <= 16'b0000_0000_0000_0000;
array[28209] <= 16'b0000_0000_0000_0000;
array[28210] <= 16'b0000_0000_0000_0000;
array[28211] <= 16'b0000_0000_0000_0000;
array[28212] <= 16'b0000_0000_0000_0000;
array[28213] <= 16'b0000_0000_0000_0000;
array[28214] <= 16'b0000_0000_0000_0000;
array[28215] <= 16'b0000_0000_0000_0000;
array[28216] <= 16'b0000_0000_0000_0000;
array[28217] <= 16'b0000_0000_0000_0000;
array[28218] <= 16'b0000_0000_0000_0000;
array[28219] <= 16'b0000_0000_0000_0000;
array[28220] <= 16'b0000_0000_0000_0000;
array[28221] <= 16'b0000_0000_0000_0000;
array[28222] <= 16'b0000_0000_0000_0000;
array[28223] <= 16'b0000_0000_0000_0000;
array[28224] <= 16'b0000_0000_0000_0000;
array[28225] <= 16'b0000_0000_0000_0000;
array[28226] <= 16'b0000_0000_0000_0000;
array[28227] <= 16'b0000_0000_0000_0000;
array[28228] <= 16'b0000_0000_0000_0000;
array[28229] <= 16'b0000_0000_0000_0000;
array[28230] <= 16'b0000_0000_0000_0000;
array[28231] <= 16'b0000_0000_0000_0000;
array[28232] <= 16'b0000_0000_0000_0000;
array[28233] <= 16'b0000_0000_0000_0000;
array[28234] <= 16'b0000_0000_0000_0000;
array[28235] <= 16'b0000_0000_0000_0000;
array[28236] <= 16'b0000_0000_0000_0000;
array[28237] <= 16'b0000_0000_0000_0000;
array[28238] <= 16'b0000_0000_0000_0000;
array[28239] <= 16'b0000_0000_0000_0000;
array[28240] <= 16'b0000_0000_0000_0000;
array[28241] <= 16'b0000_0000_0000_0000;
array[28242] <= 16'b0000_0000_0000_0000;
array[28243] <= 16'b0000_0000_0000_0000;
array[28244] <= 16'b0000_0000_0000_0000;
array[28245] <= 16'b0000_0000_0000_0000;
array[28246] <= 16'b0000_0000_0000_0000;
array[28247] <= 16'b0000_0000_0000_0000;
array[28248] <= 16'b0000_0000_0000_0000;
array[28249] <= 16'b0000_0000_0000_0000;
array[28250] <= 16'b0000_0000_0000_0000;
array[28251] <= 16'b0000_0000_0000_0000;
array[28252] <= 16'b0000_0000_0000_0000;
array[28253] <= 16'b0000_0000_0000_0000;
array[28254] <= 16'b0000_0000_0000_0000;
array[28255] <= 16'b0000_0000_0000_0000;
array[28256] <= 16'b0000_0000_0000_0000;
array[28257] <= 16'b0000_0000_0000_0000;
array[28258] <= 16'b0000_0000_0000_0000;
array[28259] <= 16'b0000_0000_0000_0000;
array[28260] <= 16'b0000_0000_0000_0000;
array[28261] <= 16'b0000_0000_0000_0000;
array[28262] <= 16'b0000_0000_0000_0000;
array[28263] <= 16'b0000_0000_0000_0000;
array[28264] <= 16'b0000_0000_0000_0000;
array[28265] <= 16'b0000_0000_0000_0000;
array[28266] <= 16'b0000_0000_0000_0000;
array[28267] <= 16'b0000_0000_0000_0000;
array[28268] <= 16'b0000_0000_0000_0000;
array[28269] <= 16'b0000_0000_0000_0000;
array[28270] <= 16'b0000_0000_0000_0000;
array[28271] <= 16'b0000_0000_0000_0000;
array[28272] <= 16'b0000_0000_0000_0000;
array[28273] <= 16'b0000_0000_0000_0000;
array[28274] <= 16'b0000_0000_0000_0000;
array[28275] <= 16'b0000_0000_0000_0000;
array[28276] <= 16'b0000_0000_0000_0000;
array[28277] <= 16'b0000_0000_0000_0000;
array[28278] <= 16'b0000_0000_0000_0000;
array[28279] <= 16'b0000_0000_0000_0000;
array[28280] <= 16'b0000_0000_0000_0000;
array[28281] <= 16'b0000_0000_0000_0000;
array[28282] <= 16'b0000_0000_0000_0000;
array[28283] <= 16'b0000_0000_0000_0000;
array[28284] <= 16'b0000_0000_0000_0000;
array[28285] <= 16'b0000_0000_0000_0000;
array[28286] <= 16'b0000_0000_0000_0000;
array[28287] <= 16'b0000_0000_0000_0000;
array[28288] <= 16'b0000_0000_0000_0000;
array[28289] <= 16'b0000_0000_0000_0000;
array[28290] <= 16'b0000_0000_0000_0000;
array[28291] <= 16'b0000_0000_0000_0000;
array[28292] <= 16'b0000_0000_0000_0000;
array[28293] <= 16'b0000_0000_0000_0000;
array[28294] <= 16'b0000_0000_0000_0000;
array[28295] <= 16'b0000_0000_0000_0000;
array[28296] <= 16'b0000_0000_0000_0000;
array[28297] <= 16'b0000_0000_0000_0000;
array[28298] <= 16'b0000_0000_0000_0000;
array[28299] <= 16'b0000_0000_0000_0000;
array[28300] <= 16'b0000_0000_0000_0000;
array[28301] <= 16'b0000_0000_0000_0000;
array[28302] <= 16'b0000_0000_0000_0000;
array[28303] <= 16'b0000_0000_0000_0000;
array[28304] <= 16'b0000_0000_0000_0000;
array[28305] <= 16'b0000_0000_0000_0000;
array[28306] <= 16'b0000_0000_0000_0000;
array[28307] <= 16'b0000_0000_0000_0000;
array[28308] <= 16'b0000_0000_0000_0000;
array[28309] <= 16'b0000_0000_0000_0000;
array[28310] <= 16'b0000_0000_0000_0000;
array[28311] <= 16'b0000_0000_0000_0000;
array[28312] <= 16'b0000_0000_0000_0000;
array[28313] <= 16'b0000_0000_0000_0000;
array[28314] <= 16'b0000_0000_0000_0000;
array[28315] <= 16'b0000_0000_0000_0000;
array[28316] <= 16'b0000_0000_0000_0000;
array[28317] <= 16'b0000_0000_0000_0000;
array[28318] <= 16'b0000_0000_0000_0000;
array[28319] <= 16'b0000_0000_0000_0000;
array[28320] <= 16'b0000_0000_0000_0000;
array[28321] <= 16'b0000_0000_0000_0000;
array[28322] <= 16'b0000_0000_0000_0000;
array[28323] <= 16'b0000_0000_0000_0000;
array[28324] <= 16'b0000_0000_0000_0000;
array[28325] <= 16'b0000_0000_0000_0000;
array[28326] <= 16'b0000_0000_0000_0000;
array[28327] <= 16'b0000_0000_0000_0000;
array[28328] <= 16'b0000_0000_0000_0000;
array[28329] <= 16'b0000_0000_0000_0000;
array[28330] <= 16'b0000_0000_0000_0000;
array[28331] <= 16'b0000_0000_0000_0000;
array[28332] <= 16'b0000_0000_0000_0000;
array[28333] <= 16'b0000_0000_0000_0000;
array[28334] <= 16'b0000_0000_0000_0000;
array[28335] <= 16'b0000_0000_0000_0000;
array[28336] <= 16'b0000_0000_0000_0000;
array[28337] <= 16'b0000_0000_0000_0000;
array[28338] <= 16'b0000_0000_0000_0000;
array[28339] <= 16'b0000_0000_0000_0000;
array[28340] <= 16'b0000_0000_0000_0000;
array[28341] <= 16'b0000_0000_0000_0000;
array[28342] <= 16'b0000_0000_0000_0000;
array[28343] <= 16'b0000_0000_0000_0000;
array[28344] <= 16'b0000_0000_0000_0000;
array[28345] <= 16'b0000_0000_0000_0000;
array[28346] <= 16'b0000_0000_0000_0000;
array[28347] <= 16'b0000_0000_0000_0000;
array[28348] <= 16'b0000_0000_0000_0000;
array[28349] <= 16'b0000_0000_0000_0000;
array[28350] <= 16'b0000_0000_0000_0000;
array[28351] <= 16'b0000_0000_0000_0000;
array[28352] <= 16'b0000_0000_0000_0000;
array[28353] <= 16'b0000_0000_0000_0000;
array[28354] <= 16'b0000_0000_0000_0000;
array[28355] <= 16'b0000_0000_0000_0000;
array[28356] <= 16'b0000_0000_0000_0000;
array[28357] <= 16'b0000_0000_0000_0000;
array[28358] <= 16'b0000_0000_0000_0000;
array[28359] <= 16'b0000_0000_0000_0000;
array[28360] <= 16'b0000_0000_0000_0000;
array[28361] <= 16'b0000_0000_0000_0000;
array[28362] <= 16'b0000_0000_0000_0000;
array[28363] <= 16'b0000_0000_0000_0000;
array[28364] <= 16'b0000_0000_0000_0000;
array[28365] <= 16'b0000_0000_0000_0000;
array[28366] <= 16'b0000_0000_0000_0000;
array[28367] <= 16'b0000_0000_0000_0000;
array[28368] <= 16'b0000_0000_0000_0000;
array[28369] <= 16'b0000_0000_0000_0000;
array[28370] <= 16'b0000_0000_0000_0000;
array[28371] <= 16'b0000_0000_0000_0000;
array[28372] <= 16'b0000_0000_0000_0000;
array[28373] <= 16'b0000_0000_0000_0000;
array[28374] <= 16'b0000_0000_0000_0000;
array[28375] <= 16'b0000_0000_0000_0000;
array[28376] <= 16'b0000_0000_0000_0000;
array[28377] <= 16'b0000_0000_0000_0000;
array[28378] <= 16'b0000_0000_0000_0000;
array[28379] <= 16'b0000_0000_0000_0000;
array[28380] <= 16'b0000_0000_0000_0000;
array[28381] <= 16'b0000_0000_0000_0000;
array[28382] <= 16'b0000_0000_0000_0000;
array[28383] <= 16'b0000_0000_0000_0000;
array[28384] <= 16'b0000_0000_0000_0000;
array[28385] <= 16'b0000_0000_0000_0000;
array[28386] <= 16'b0000_0000_0000_0000;
array[28387] <= 16'b0000_0000_0000_0000;
array[28388] <= 16'b0000_0000_0000_0000;
array[28389] <= 16'b0000_0000_0000_0000;
array[28390] <= 16'b0000_0000_0000_0000;
array[28391] <= 16'b0000_0000_0000_0000;
array[28392] <= 16'b0000_0000_0000_0000;
array[28393] <= 16'b0000_0000_0000_0000;
array[28394] <= 16'b0000_0000_0000_0000;
array[28395] <= 16'b0000_0000_0000_0000;
array[28396] <= 16'b0000_0000_0000_0000;
array[28397] <= 16'b0000_0000_0000_0000;
array[28398] <= 16'b0000_0000_0000_0000;
array[28399] <= 16'b0000_0000_0000_0000;
array[28400] <= 16'b0000_0000_0000_0000;
array[28401] <= 16'b0000_0000_0000_0000;
array[28402] <= 16'b0000_0000_0000_0000;
array[28403] <= 16'b0000_0000_0000_0000;
array[28404] <= 16'b0000_0000_0000_0000;
array[28405] <= 16'b0000_0000_0000_0000;
array[28406] <= 16'b0000_0000_0000_0000;
array[28407] <= 16'b0000_0000_0000_0000;
array[28408] <= 16'b0000_0000_0000_0000;
array[28409] <= 16'b0000_0000_0000_0000;
array[28410] <= 16'b0000_0000_0000_0000;
array[28411] <= 16'b0000_0000_0000_0000;
array[28412] <= 16'b0000_0000_0000_0000;
array[28413] <= 16'b0000_0000_0000_0000;
array[28414] <= 16'b0000_0000_0000_0000;
array[28415] <= 16'b0000_0000_0000_0000;
array[28416] <= 16'b0000_0000_0000_0000;
array[28417] <= 16'b0000_0000_0000_0000;
array[28418] <= 16'b0000_0000_0000_0000;
array[28419] <= 16'b0000_0000_0000_0000;
array[28420] <= 16'b0000_0000_0000_0000;
array[28421] <= 16'b0000_0000_0000_0000;
array[28422] <= 16'b0000_0000_0000_0000;
array[28423] <= 16'b0000_0000_0000_0000;
array[28424] <= 16'b0000_0000_0000_0000;
array[28425] <= 16'b0000_0000_0000_0000;
array[28426] <= 16'b0000_0000_0000_0000;
array[28427] <= 16'b0000_0000_0000_0000;
array[28428] <= 16'b0000_0000_0000_0000;
array[28429] <= 16'b0000_0000_0000_0000;
array[28430] <= 16'b0000_0000_0000_0000;
array[28431] <= 16'b0000_0000_0000_0000;
array[28432] <= 16'b0000_0000_0000_0000;
array[28433] <= 16'b0000_0000_0000_0000;
array[28434] <= 16'b0000_0000_0000_0000;
array[28435] <= 16'b0000_0000_0000_0000;
array[28436] <= 16'b0000_0000_0000_0000;
array[28437] <= 16'b0000_0000_0000_0000;
array[28438] <= 16'b0000_0000_0000_0000;
array[28439] <= 16'b0000_0000_0000_0000;
array[28440] <= 16'b0000_0000_0000_0000;
array[28441] <= 16'b0000_0000_0000_0000;
array[28442] <= 16'b0000_0000_0000_0000;
array[28443] <= 16'b0000_0000_0000_0000;
array[28444] <= 16'b0000_0000_0000_0000;
array[28445] <= 16'b0000_0000_0000_0000;
array[28446] <= 16'b0000_0000_0000_0000;
array[28447] <= 16'b0000_0000_0000_0000;
array[28448] <= 16'b0000_0000_0000_0000;
array[28449] <= 16'b0000_0000_0000_0000;
array[28450] <= 16'b0000_0000_0000_0000;
array[28451] <= 16'b0000_0000_0000_0000;
array[28452] <= 16'b0000_0000_0000_0000;
array[28453] <= 16'b0000_0000_0000_0000;
array[28454] <= 16'b0000_0000_0000_0000;
array[28455] <= 16'b0000_0000_0000_0000;
array[28456] <= 16'b0000_0000_0000_0000;
array[28457] <= 16'b0000_0000_0000_0000;
array[28458] <= 16'b0000_0000_0000_0000;
array[28459] <= 16'b0000_0000_0000_0000;
array[28460] <= 16'b0000_0000_0000_0000;
array[28461] <= 16'b0000_0000_0000_0000;
array[28462] <= 16'b0000_0000_0000_0000;
array[28463] <= 16'b0000_0000_0000_0000;
array[28464] <= 16'b0000_0000_0000_0000;
array[28465] <= 16'b0000_0000_0000_0000;
array[28466] <= 16'b0000_0000_0000_0000;
array[28467] <= 16'b0000_0000_0000_0000;
array[28468] <= 16'b0000_0000_0000_0000;
array[28469] <= 16'b0000_0000_0000_0000;
array[28470] <= 16'b0000_0000_0000_0000;
array[28471] <= 16'b0000_0000_0000_0000;
array[28472] <= 16'b0000_0000_0000_0000;
array[28473] <= 16'b0000_0000_0000_0000;
array[28474] <= 16'b0000_0000_0000_0000;
array[28475] <= 16'b0000_0000_0000_0000;
array[28476] <= 16'b0000_0000_0000_0000;
array[28477] <= 16'b0000_0000_0000_0000;
array[28478] <= 16'b0000_0000_0000_0000;
array[28479] <= 16'b0000_0000_0000_0000;
array[28480] <= 16'b0000_0000_0000_0000;
array[28481] <= 16'b0000_0000_0000_0000;
array[28482] <= 16'b0000_0000_0000_0000;
array[28483] <= 16'b0000_0000_0000_0000;
array[28484] <= 16'b0000_0000_0000_0000;
array[28485] <= 16'b0000_0000_0000_0000;
array[28486] <= 16'b0000_0000_0000_0000;
array[28487] <= 16'b0000_0000_0000_0000;
array[28488] <= 16'b0000_0000_0000_0000;
array[28489] <= 16'b0000_0000_0000_0000;
array[28490] <= 16'b0000_0000_0000_0000;
array[28491] <= 16'b0000_0000_0000_0000;
array[28492] <= 16'b0000_0000_0000_0000;
array[28493] <= 16'b0000_0000_0000_0000;
array[28494] <= 16'b0000_0000_0000_0000;
array[28495] <= 16'b0000_0000_0000_0000;
array[28496] <= 16'b0000_0000_0000_0000;
array[28497] <= 16'b0000_0000_0000_0000;
array[28498] <= 16'b0000_0000_0000_0000;
array[28499] <= 16'b0000_0000_0000_0000;
array[28500] <= 16'b0000_0000_0000_0000;
array[28501] <= 16'b0000_0000_0000_0000;
array[28502] <= 16'b0000_0000_0000_0000;
array[28503] <= 16'b0000_0000_0000_0000;
array[28504] <= 16'b0000_0000_0000_0000;
array[28505] <= 16'b0000_0000_0000_0000;
array[28506] <= 16'b0000_0000_0000_0000;
array[28507] <= 16'b0000_0000_0000_0000;
array[28508] <= 16'b0000_0000_0000_0000;
array[28509] <= 16'b0000_0000_0000_0000;
array[28510] <= 16'b0000_0000_0000_0000;
array[28511] <= 16'b0000_0000_0000_0000;
array[28512] <= 16'b0000_0000_0000_0000;
array[28513] <= 16'b0000_0000_0000_0000;
array[28514] <= 16'b0000_0000_0000_0000;
array[28515] <= 16'b0000_0000_0000_0000;
array[28516] <= 16'b0000_0000_0000_0000;
array[28517] <= 16'b0000_0000_0000_0000;
array[28518] <= 16'b0000_0000_0000_0000;
array[28519] <= 16'b0000_0000_0000_0000;
array[28520] <= 16'b0000_0000_0000_0000;
array[28521] <= 16'b0000_0000_0000_0000;
array[28522] <= 16'b0000_0000_0000_0000;
array[28523] <= 16'b0000_0000_0000_0000;
array[28524] <= 16'b0000_0000_0000_0000;
array[28525] <= 16'b0000_0000_0000_0000;
array[28526] <= 16'b0000_0000_0000_0000;
array[28527] <= 16'b0000_0000_0000_0000;
array[28528] <= 16'b0000_0000_0000_0000;
array[28529] <= 16'b0000_0000_0000_0000;
array[28530] <= 16'b0000_0000_0000_0000;
array[28531] <= 16'b0000_0000_0000_0000;
array[28532] <= 16'b0000_0000_0000_0000;
array[28533] <= 16'b0000_0000_0000_0000;
array[28534] <= 16'b0000_0000_0000_0000;
array[28535] <= 16'b0000_0000_0000_0000;
array[28536] <= 16'b0000_0000_0000_0000;
array[28537] <= 16'b0000_0000_0000_0000;
array[28538] <= 16'b0000_0000_0000_0000;
array[28539] <= 16'b0000_0000_0000_0000;
array[28540] <= 16'b0000_0000_0000_0000;
array[28541] <= 16'b0000_0000_0000_0000;
array[28542] <= 16'b0000_0000_0000_0000;
array[28543] <= 16'b0000_0000_0000_0000;
array[28544] <= 16'b0000_0000_0000_0000;
array[28545] <= 16'b0000_0000_0000_0000;
array[28546] <= 16'b0000_0000_0000_0000;
array[28547] <= 16'b0000_0000_0000_0000;
array[28548] <= 16'b0000_0000_0000_0000;
array[28549] <= 16'b0000_0000_0000_0000;
array[28550] <= 16'b0000_0000_0000_0000;
array[28551] <= 16'b0000_0000_0000_0000;
array[28552] <= 16'b0000_0000_0000_0000;
array[28553] <= 16'b0000_0000_0000_0000;
array[28554] <= 16'b0000_0000_0000_0000;
array[28555] <= 16'b0000_0000_0000_0000;
array[28556] <= 16'b0000_0000_0000_0000;
array[28557] <= 16'b0000_0000_0000_0000;
array[28558] <= 16'b0000_0000_0000_0000;
array[28559] <= 16'b0000_0000_0000_0000;
array[28560] <= 16'b0000_0000_0000_0000;
array[28561] <= 16'b0000_0000_0000_0000;
array[28562] <= 16'b0000_0000_0000_0000;
array[28563] <= 16'b0000_0000_0000_0000;
array[28564] <= 16'b0000_0000_0000_0000;
array[28565] <= 16'b0000_0000_0000_0000;
array[28566] <= 16'b0000_0000_0000_0000;
array[28567] <= 16'b0000_0000_0000_0000;
array[28568] <= 16'b0000_0000_0000_0000;
array[28569] <= 16'b0000_0000_0000_0000;
array[28570] <= 16'b0000_0000_0000_0000;
array[28571] <= 16'b0000_0000_0000_0000;
array[28572] <= 16'b0000_0000_0000_0000;
array[28573] <= 16'b0000_0000_0000_0000;
array[28574] <= 16'b0000_0000_0000_0000;
array[28575] <= 16'b0000_0000_0000_0000;
array[28576] <= 16'b0000_0000_0000_0000;
array[28577] <= 16'b0000_0000_0000_0000;
array[28578] <= 16'b0000_0000_0000_0000;
array[28579] <= 16'b0000_0000_0000_0000;
array[28580] <= 16'b0000_0000_0000_0000;
array[28581] <= 16'b0000_0000_0000_0000;
array[28582] <= 16'b0000_0000_0000_0000;
array[28583] <= 16'b0000_0000_0000_0000;
array[28584] <= 16'b0000_0000_0000_0000;
array[28585] <= 16'b0000_0000_0000_0000;
array[28586] <= 16'b0000_0000_0000_0000;
array[28587] <= 16'b0000_0000_0000_0000;
array[28588] <= 16'b0000_0000_0000_0000;
array[28589] <= 16'b0000_0000_0000_0000;
array[28590] <= 16'b0000_0000_0000_0000;
array[28591] <= 16'b0000_0000_0000_0000;
array[28592] <= 16'b0000_0000_0000_0000;
array[28593] <= 16'b0000_0000_0000_0000;
array[28594] <= 16'b0000_0000_0000_0000;
array[28595] <= 16'b0000_0000_0000_0000;
array[28596] <= 16'b0000_0000_0000_0000;
array[28597] <= 16'b0000_0000_0000_0000;
array[28598] <= 16'b0000_0000_0000_0000;
array[28599] <= 16'b0000_0000_0000_0000;
array[28600] <= 16'b0000_0000_0000_0000;
array[28601] <= 16'b0000_0000_0000_0000;
array[28602] <= 16'b0000_0000_0000_0000;
array[28603] <= 16'b0000_0000_0000_0000;
array[28604] <= 16'b0000_0000_0000_0000;
array[28605] <= 16'b0000_0000_0000_0000;
array[28606] <= 16'b0000_0000_0000_0000;
array[28607] <= 16'b0000_0000_0000_0000;
array[28608] <= 16'b0000_0000_0000_0000;
array[28609] <= 16'b0000_0000_0000_0000;
array[28610] <= 16'b0000_0000_0000_0000;
array[28611] <= 16'b0000_0000_0000_0000;
array[28612] <= 16'b0000_0000_0000_0000;
array[28613] <= 16'b0000_0000_0000_0000;
array[28614] <= 16'b0000_0000_0000_0000;
array[28615] <= 16'b0000_0000_0000_0000;
array[28616] <= 16'b0000_0000_0000_0000;
array[28617] <= 16'b0000_0000_0000_0000;
array[28618] <= 16'b0000_0000_0000_0000;
array[28619] <= 16'b0000_0000_0000_0000;
array[28620] <= 16'b0000_0000_0000_0000;
array[28621] <= 16'b0000_0000_0000_0000;
array[28622] <= 16'b0000_0000_0000_0000;
array[28623] <= 16'b0000_0000_0000_0000;
array[28624] <= 16'b0000_0000_0000_0000;
array[28625] <= 16'b0000_0000_0000_0000;
array[28626] <= 16'b0000_0000_0000_0000;
array[28627] <= 16'b0000_0000_0000_0000;
array[28628] <= 16'b0000_0000_0000_0000;
array[28629] <= 16'b0000_0000_0000_0000;
array[28630] <= 16'b0000_0000_0000_0000;
array[28631] <= 16'b0000_0000_0000_0000;
array[28632] <= 16'b0000_0000_0000_0000;
array[28633] <= 16'b0000_0000_0000_0000;
array[28634] <= 16'b0000_0000_0000_0000;
array[28635] <= 16'b0000_0000_0000_0000;
array[28636] <= 16'b0000_0000_0000_0000;
array[28637] <= 16'b0000_0000_0000_0000;
array[28638] <= 16'b0000_0000_0000_0000;
array[28639] <= 16'b0000_0000_0000_0000;
array[28640] <= 16'b0000_0000_0000_0000;
array[28641] <= 16'b0000_0000_0000_0000;
array[28642] <= 16'b0000_0000_0000_0000;
array[28643] <= 16'b0000_0000_0000_0000;
array[28644] <= 16'b0000_0000_0000_0000;
array[28645] <= 16'b0000_0000_0000_0000;
array[28646] <= 16'b0000_0000_0000_0000;
array[28647] <= 16'b0000_0000_0000_0000;
array[28648] <= 16'b0000_0000_0000_0000;
array[28649] <= 16'b0000_0000_0000_0000;
array[28650] <= 16'b0000_0000_0000_0000;
array[28651] <= 16'b0000_0000_0000_0000;
array[28652] <= 16'b0000_0000_0000_0000;
array[28653] <= 16'b0000_0000_0000_0000;
array[28654] <= 16'b0000_0000_0000_0000;
array[28655] <= 16'b0000_0000_0000_0000;
array[28656] <= 16'b0000_0000_0000_0000;
array[28657] <= 16'b0000_0000_0000_0000;
array[28658] <= 16'b0000_0000_0000_0000;
array[28659] <= 16'b0000_0000_0000_0000;
array[28660] <= 16'b0000_0000_0000_0000;
array[28661] <= 16'b0000_0000_0000_0000;
array[28662] <= 16'b0000_0000_0000_0000;
array[28663] <= 16'b0000_0000_0000_0000;
array[28664] <= 16'b0000_0000_0000_0000;
array[28665] <= 16'b0000_0000_0000_0000;
array[28666] <= 16'b0000_0000_0000_0000;
array[28667] <= 16'b0000_0000_0000_0000;
array[28668] <= 16'b0000_0000_0000_0000;
array[28669] <= 16'b0000_0000_0000_0000;
array[28670] <= 16'b0000_0000_0000_0000;
array[28671] <= 16'b0000_0000_0000_0000;
array[28672] <= 16'b0000_0000_0000_0000;
array[28673] <= 16'b0000_0000_0000_0000;
array[28674] <= 16'b0000_0000_0000_0000;
array[28675] <= 16'b0000_0000_0000_0000;
array[28676] <= 16'b0000_0000_0000_0000;
array[28677] <= 16'b0000_0000_0000_0000;
array[28678] <= 16'b0000_0000_0000_0000;
array[28679] <= 16'b0000_0000_0000_0000;
array[28680] <= 16'b0000_0000_0000_0000;
array[28681] <= 16'b0000_0000_0000_0000;
array[28682] <= 16'b0000_0000_0000_0000;
array[28683] <= 16'b0000_0000_0000_0000;
array[28684] <= 16'b0000_0000_0000_0000;
array[28685] <= 16'b0000_0000_0000_0000;
array[28686] <= 16'b0000_0000_0000_0000;
array[28687] <= 16'b0000_0000_0000_0000;
array[28688] <= 16'b0000_0000_0000_0000;
array[28689] <= 16'b0000_0000_0000_0000;
array[28690] <= 16'b0000_0000_0000_0000;
array[28691] <= 16'b0000_0000_0000_0000;
array[28692] <= 16'b0000_0000_0000_0000;
array[28693] <= 16'b0000_0000_0000_0000;
array[28694] <= 16'b0000_0000_0000_0000;
array[28695] <= 16'b0000_0000_0000_0000;
array[28696] <= 16'b0000_0000_0000_0000;
array[28697] <= 16'b0000_0000_0000_0000;
array[28698] <= 16'b0000_0000_0000_0000;
array[28699] <= 16'b0000_0000_0000_0000;
array[28700] <= 16'b0000_0000_0000_0000;
array[28701] <= 16'b0000_0000_0000_0000;
array[28702] <= 16'b0000_0000_0000_0000;
array[28703] <= 16'b0000_0000_0000_0000;
array[28704] <= 16'b0000_0000_0000_0000;
array[28705] <= 16'b0000_0000_0000_0000;
array[28706] <= 16'b0000_0000_0000_0000;
array[28707] <= 16'b0000_0000_0000_0000;
array[28708] <= 16'b0000_0000_0000_0000;
array[28709] <= 16'b0000_0000_0000_0000;
array[28710] <= 16'b0000_0000_0000_0000;
array[28711] <= 16'b0000_0000_0000_0000;
array[28712] <= 16'b0000_0000_0000_0000;
array[28713] <= 16'b0000_0000_0000_0000;
array[28714] <= 16'b0000_0000_0000_0000;
array[28715] <= 16'b0000_0000_0000_0000;
array[28716] <= 16'b0000_0000_0000_0000;
array[28717] <= 16'b0000_0000_0000_0000;
array[28718] <= 16'b0000_0000_0000_0000;
array[28719] <= 16'b0000_0000_0000_0000;
array[28720] <= 16'b0000_0000_0000_0000;
array[28721] <= 16'b0000_0000_0000_0000;
array[28722] <= 16'b0000_0000_0000_0000;
array[28723] <= 16'b0000_0000_0000_0000;
array[28724] <= 16'b0000_0000_0000_0000;
array[28725] <= 16'b0000_0000_0000_0000;
array[28726] <= 16'b0000_0000_0000_0000;
array[28727] <= 16'b0000_0000_0000_0000;
array[28728] <= 16'b0000_0000_0000_0000;
array[28729] <= 16'b0000_0000_0000_0000;
array[28730] <= 16'b0000_0000_0000_0000;
array[28731] <= 16'b0000_0000_0000_0000;
array[28732] <= 16'b0000_0000_0000_0000;
array[28733] <= 16'b0000_0000_0000_0000;
array[28734] <= 16'b0000_0000_0000_0000;
array[28735] <= 16'b0000_0000_0000_0000;
array[28736] <= 16'b0000_0000_0000_0000;
array[28737] <= 16'b0000_0000_0000_0000;
array[28738] <= 16'b0000_0000_0000_0000;
array[28739] <= 16'b0000_0000_0000_0000;
array[28740] <= 16'b0000_0000_0000_0000;
array[28741] <= 16'b0000_0000_0000_0000;
array[28742] <= 16'b0000_0000_0000_0000;
array[28743] <= 16'b0000_0000_0000_0000;
array[28744] <= 16'b0000_0000_0000_0000;
array[28745] <= 16'b0000_0000_0000_0000;
array[28746] <= 16'b0000_0000_0000_0000;
array[28747] <= 16'b0000_0000_0000_0000;
array[28748] <= 16'b0000_0000_0000_0000;
array[28749] <= 16'b0000_0000_0000_0000;
array[28750] <= 16'b0000_0000_0000_0000;
array[28751] <= 16'b0000_0000_0000_0000;
array[28752] <= 16'b0000_0000_0000_0000;
array[28753] <= 16'b0000_0000_0000_0000;
array[28754] <= 16'b0000_0000_0000_0000;
array[28755] <= 16'b0000_0000_0000_0000;
array[28756] <= 16'b0000_0000_0000_0000;
array[28757] <= 16'b0000_0000_0000_0000;
array[28758] <= 16'b0000_0000_0000_0000;
array[28759] <= 16'b0000_0000_0000_0000;
array[28760] <= 16'b0000_0000_0000_0000;
array[28761] <= 16'b0000_0000_0000_0000;
array[28762] <= 16'b0000_0000_0000_0000;
array[28763] <= 16'b0000_0000_0000_0000;
array[28764] <= 16'b0000_0000_0000_0000;
array[28765] <= 16'b0000_0000_0000_0000;
array[28766] <= 16'b0000_0000_0000_0000;
array[28767] <= 16'b0000_0000_0000_0000;
array[28768] <= 16'b0000_0000_0000_0000;
array[28769] <= 16'b0000_0000_0000_0000;
array[28770] <= 16'b0000_0000_0000_0000;
array[28771] <= 16'b0000_0000_0000_0000;
array[28772] <= 16'b0000_0000_0000_0000;
array[28773] <= 16'b0000_0000_0000_0000;
array[28774] <= 16'b0000_0000_0000_0000;
array[28775] <= 16'b0000_0000_0000_0000;
array[28776] <= 16'b0000_0000_0000_0000;
array[28777] <= 16'b0000_0000_0000_0000;
array[28778] <= 16'b0000_0000_0000_0000;
array[28779] <= 16'b0000_0000_0000_0000;
array[28780] <= 16'b0000_0000_0000_0000;
array[28781] <= 16'b0000_0000_0000_0000;
array[28782] <= 16'b0000_0000_0000_0000;
array[28783] <= 16'b0000_0000_0000_0000;
array[28784] <= 16'b0000_0000_0000_0000;
array[28785] <= 16'b0000_0000_0000_0000;
array[28786] <= 16'b0000_0000_0000_0000;
array[28787] <= 16'b0000_0000_0000_0000;
array[28788] <= 16'b0000_0000_0000_0000;
array[28789] <= 16'b0000_0000_0000_0000;
array[28790] <= 16'b0000_0000_0000_0000;
array[28791] <= 16'b0000_0000_0000_0000;
array[28792] <= 16'b0000_0000_0000_0000;
array[28793] <= 16'b0000_0000_0000_0000;
array[28794] <= 16'b0000_0000_0000_0000;
array[28795] <= 16'b0000_0000_0000_0000;
array[28796] <= 16'b0000_0000_0000_0000;
array[28797] <= 16'b0000_0000_0000_0000;
array[28798] <= 16'b0000_0000_0000_0000;
array[28799] <= 16'b0000_0000_0000_0000;
array[28800] <= 16'b0000_0000_0000_0000;
array[28801] <= 16'b0000_0000_0000_0000;
array[28802] <= 16'b0000_0000_0000_0000;
array[28803] <= 16'b0000_0000_0000_0000;
array[28804] <= 16'b0000_0000_0000_0000;
array[28805] <= 16'b0000_0000_0000_0000;
array[28806] <= 16'b0000_0000_0000_0000;
array[28807] <= 16'b0000_0000_0000_0000;
array[28808] <= 16'b0000_0000_0000_0000;
array[28809] <= 16'b0000_0000_0000_0000;
array[28810] <= 16'b0000_0000_0000_0000;
array[28811] <= 16'b0000_0000_0000_0000;
array[28812] <= 16'b0000_0000_0000_0000;
array[28813] <= 16'b0000_0000_0000_0000;
array[28814] <= 16'b0000_0000_0000_0000;
array[28815] <= 16'b0000_0000_0000_0000;
array[28816] <= 16'b0000_0000_0000_0000;
array[28817] <= 16'b0000_0000_0000_0000;
array[28818] <= 16'b0000_0000_0000_0000;
array[28819] <= 16'b0000_0000_0000_0000;
array[28820] <= 16'b0000_0000_0000_0000;
array[28821] <= 16'b0000_0000_0000_0000;
array[28822] <= 16'b0000_0000_0000_0000;
array[28823] <= 16'b0000_0000_0000_0000;
array[28824] <= 16'b0000_0000_0000_0000;
array[28825] <= 16'b0000_0000_0000_0000;
array[28826] <= 16'b0000_0000_0000_0000;
array[28827] <= 16'b0000_0000_0000_0000;
array[28828] <= 16'b0000_0000_0000_0000;
array[28829] <= 16'b0000_0000_0000_0000;
array[28830] <= 16'b0000_0000_0000_0000;
array[28831] <= 16'b0000_0000_0000_0000;
array[28832] <= 16'b0000_0000_0000_0000;
array[28833] <= 16'b0000_0000_0000_0000;
array[28834] <= 16'b0000_0000_0000_0000;
array[28835] <= 16'b0000_0000_0000_0000;
array[28836] <= 16'b0000_0000_0000_0000;
array[28837] <= 16'b0000_0000_0000_0000;
array[28838] <= 16'b0000_0000_0000_0000;
array[28839] <= 16'b0000_0000_0000_0000;
array[28840] <= 16'b0000_0000_0000_0000;
array[28841] <= 16'b0000_0000_0000_0000;
array[28842] <= 16'b0000_0000_0000_0000;
array[28843] <= 16'b0000_0000_0000_0000;
array[28844] <= 16'b0000_0000_0000_0000;
array[28845] <= 16'b0000_0000_0000_0000;
array[28846] <= 16'b0000_0000_0000_0000;
array[28847] <= 16'b0000_0000_0000_0000;
array[28848] <= 16'b0000_0000_0000_0000;
array[28849] <= 16'b0000_0000_0000_0000;
array[28850] <= 16'b0000_0000_0000_0000;
array[28851] <= 16'b0000_0000_0000_0000;
array[28852] <= 16'b0000_0000_0000_0000;
array[28853] <= 16'b0000_0000_0000_0000;
array[28854] <= 16'b0000_0000_0000_0000;
array[28855] <= 16'b0000_0000_0000_0000;
array[28856] <= 16'b0000_0000_0000_0000;
array[28857] <= 16'b0000_0000_0000_0000;
array[28858] <= 16'b0000_0000_0000_0000;
array[28859] <= 16'b0000_0000_0000_0000;
array[28860] <= 16'b0000_0000_0000_0000;
array[28861] <= 16'b0000_0000_0000_0000;
array[28862] <= 16'b0000_0000_0000_0000;
array[28863] <= 16'b0000_0000_0000_0000;
array[28864] <= 16'b0000_0000_0000_0000;
array[28865] <= 16'b0000_0000_0000_0000;
array[28866] <= 16'b0000_0000_0000_0000;
array[28867] <= 16'b0000_0000_0000_0000;
array[28868] <= 16'b0000_0000_0000_0000;
array[28869] <= 16'b0000_0000_0000_0000;
array[28870] <= 16'b0000_0000_0000_0000;
array[28871] <= 16'b0000_0000_0000_0000;
array[28872] <= 16'b0000_0000_0000_0000;
array[28873] <= 16'b0000_0000_0000_0000;
array[28874] <= 16'b0000_0000_0000_0000;
array[28875] <= 16'b0000_0000_0000_0000;
array[28876] <= 16'b0000_0000_0000_0000;
array[28877] <= 16'b0000_0000_0000_0000;
array[28878] <= 16'b0000_0000_0000_0000;
array[28879] <= 16'b0000_0000_0000_0000;
array[28880] <= 16'b0000_0000_0000_0000;
array[28881] <= 16'b0000_0000_0000_0000;
array[28882] <= 16'b0000_0000_0000_0000;
array[28883] <= 16'b0000_0000_0000_0000;
array[28884] <= 16'b0000_0000_0000_0000;
array[28885] <= 16'b0000_0000_0000_0000;
array[28886] <= 16'b0000_0000_0000_0000;
array[28887] <= 16'b0000_0000_0000_0000;
array[28888] <= 16'b0000_0000_0000_0000;
array[28889] <= 16'b0000_0000_0000_0000;
array[28890] <= 16'b0000_0000_0000_0000;
array[28891] <= 16'b0000_0000_0000_0000;
array[28892] <= 16'b0000_0000_0000_0000;
array[28893] <= 16'b0000_0000_0000_0000;
array[28894] <= 16'b0000_0000_0000_0000;
array[28895] <= 16'b0000_0000_0000_0000;
array[28896] <= 16'b0000_0000_0000_0000;
array[28897] <= 16'b0000_0000_0000_0000;
array[28898] <= 16'b0000_0000_0000_0000;
array[28899] <= 16'b0000_0000_0000_0000;
array[28900] <= 16'b0000_0000_0000_0000;
array[28901] <= 16'b0000_0000_0000_0000;
array[28902] <= 16'b0000_0000_0000_0000;
array[28903] <= 16'b0000_0000_0000_0000;
array[28904] <= 16'b0000_0000_0000_0000;
array[28905] <= 16'b0000_0000_0000_0000;
array[28906] <= 16'b0000_0000_0000_0000;
array[28907] <= 16'b0000_0000_0000_0000;
array[28908] <= 16'b0000_0000_0000_0000;
array[28909] <= 16'b0000_0000_0000_0000;
array[28910] <= 16'b0000_0000_0000_0000;
array[28911] <= 16'b0000_0000_0000_0000;
array[28912] <= 16'b0000_0000_0000_0000;
array[28913] <= 16'b0000_0000_0000_0000;
array[28914] <= 16'b0000_0000_0000_0000;
array[28915] <= 16'b0000_0000_0000_0000;
array[28916] <= 16'b0000_0000_0000_0000;
array[28917] <= 16'b0000_0000_0000_0000;
array[28918] <= 16'b0000_0000_0000_0000;
array[28919] <= 16'b0000_0000_0000_0000;
array[28920] <= 16'b0000_0000_0000_0000;
array[28921] <= 16'b0000_0000_0000_0000;
array[28922] <= 16'b0000_0000_0000_0000;
array[28923] <= 16'b0000_0000_0000_0000;
array[28924] <= 16'b0000_0000_0000_0000;
array[28925] <= 16'b0000_0000_0000_0000;
array[28926] <= 16'b0000_0000_0000_0000;
array[28927] <= 16'b0000_0000_0000_0000;
array[28928] <= 16'b0000_0000_0000_0000;
array[28929] <= 16'b0000_0000_0000_0000;
array[28930] <= 16'b0000_0000_0000_0000;
array[28931] <= 16'b0000_0000_0000_0000;
array[28932] <= 16'b0000_0000_0000_0000;
array[28933] <= 16'b0000_0000_0000_0000;
array[28934] <= 16'b0000_0000_0000_0000;
array[28935] <= 16'b0000_0000_0000_0000;
array[28936] <= 16'b0000_0000_0000_0000;
array[28937] <= 16'b0000_0000_0000_0000;
array[28938] <= 16'b0000_0000_0000_0000;
array[28939] <= 16'b0000_0000_0000_0000;
array[28940] <= 16'b0000_0000_0000_0000;
array[28941] <= 16'b0000_0000_0000_0000;
array[28942] <= 16'b0000_0000_0000_0000;
array[28943] <= 16'b0000_0000_0000_0000;
array[28944] <= 16'b0000_0000_0000_0000;
array[28945] <= 16'b0000_0000_0000_0000;
array[28946] <= 16'b0000_0000_0000_0000;
array[28947] <= 16'b0000_0000_0000_0000;
array[28948] <= 16'b0000_0000_0000_0000;
array[28949] <= 16'b0000_0000_0000_0000;
array[28950] <= 16'b0000_0000_0000_0000;
array[28951] <= 16'b0000_0000_0000_0000;
array[28952] <= 16'b0000_0000_0000_0000;
array[28953] <= 16'b0000_0000_0000_0000;
array[28954] <= 16'b0000_0000_0000_0000;
array[28955] <= 16'b0000_0000_0000_0000;
array[28956] <= 16'b0000_0000_0000_0000;
array[28957] <= 16'b0000_0000_0000_0000;
array[28958] <= 16'b0000_0000_0000_0000;
array[28959] <= 16'b0000_0000_0000_0000;
array[28960] <= 16'b0000_0000_0000_0000;
array[28961] <= 16'b0000_0000_0000_0000;
array[28962] <= 16'b0000_0000_0000_0000;
array[28963] <= 16'b0000_0000_0000_0000;
array[28964] <= 16'b0000_0000_0000_0000;
array[28965] <= 16'b0000_0000_0000_0000;
array[28966] <= 16'b0000_0000_0000_0000;
array[28967] <= 16'b0000_0000_0000_0000;
array[28968] <= 16'b0000_0000_0000_0000;
array[28969] <= 16'b0000_0000_0000_0000;
array[28970] <= 16'b0000_0000_0000_0000;
array[28971] <= 16'b0000_0000_0000_0000;
array[28972] <= 16'b0000_0000_0000_0000;
array[28973] <= 16'b0000_0000_0000_0000;
array[28974] <= 16'b0000_0000_0000_0000;
array[28975] <= 16'b0000_0000_0000_0000;
array[28976] <= 16'b0000_0000_0000_0000;
array[28977] <= 16'b0000_0000_0000_0000;
array[28978] <= 16'b0000_0000_0000_0000;
array[28979] <= 16'b0000_0000_0000_0000;
array[28980] <= 16'b0000_0000_0000_0000;
array[28981] <= 16'b0000_0000_0000_0000;
array[28982] <= 16'b0000_0000_0000_0000;
array[28983] <= 16'b0000_0000_0000_0000;
array[28984] <= 16'b0000_0000_0000_0000;
array[28985] <= 16'b0000_0000_0000_0000;
array[28986] <= 16'b0000_0000_0000_0000;
array[28987] <= 16'b0000_0000_0000_0000;
array[28988] <= 16'b0000_0000_0000_0000;
array[28989] <= 16'b0000_0000_0000_0000;
array[28990] <= 16'b0000_0000_0000_0000;
array[28991] <= 16'b0000_0000_0000_0000;
array[28992] <= 16'b0000_0000_0000_0000;
array[28993] <= 16'b0000_0000_0000_0000;
array[28994] <= 16'b0000_0000_0000_0000;
array[28995] <= 16'b0000_0000_0000_0000;
array[28996] <= 16'b0000_0000_0000_0000;
array[28997] <= 16'b0000_0000_0000_0000;
array[28998] <= 16'b0000_0000_0000_0000;
array[28999] <= 16'b0000_0000_0000_0000;
array[29000] <= 16'b0000_0000_0000_0000;
array[29001] <= 16'b0000_0000_0000_0000;
array[29002] <= 16'b0000_0000_0000_0000;
array[29003] <= 16'b0000_0000_0000_0000;
array[29004] <= 16'b0000_0000_0000_0000;
array[29005] <= 16'b0000_0000_0000_0000;
array[29006] <= 16'b0000_0000_0000_0000;
array[29007] <= 16'b0000_0000_0000_0000;
array[29008] <= 16'b0000_0000_0000_0000;
array[29009] <= 16'b0000_0000_0000_0000;
array[29010] <= 16'b0000_0000_0000_0000;
array[29011] <= 16'b0000_0000_0000_0000;
array[29012] <= 16'b0000_0000_0000_0000;
array[29013] <= 16'b0000_0000_0000_0000;
array[29014] <= 16'b0000_0000_0000_0000;
array[29015] <= 16'b0000_0000_0000_0000;
array[29016] <= 16'b0000_0000_0000_0000;
array[29017] <= 16'b0000_0000_0000_0000;
array[29018] <= 16'b0000_0000_0000_0000;
array[29019] <= 16'b0000_0000_0000_0000;
array[29020] <= 16'b0000_0000_0000_0000;
array[29021] <= 16'b0000_0000_0000_0000;
array[29022] <= 16'b0000_0000_0000_0000;
array[29023] <= 16'b0000_0000_0000_0000;
array[29024] <= 16'b0000_0000_0000_0000;
array[29025] <= 16'b0000_0000_0000_0000;
array[29026] <= 16'b0000_0000_0000_0000;
array[29027] <= 16'b0000_0000_0000_0000;
array[29028] <= 16'b0000_0000_0000_0000;
array[29029] <= 16'b0000_0000_0000_0000;
array[29030] <= 16'b0000_0000_0000_0000;
array[29031] <= 16'b0000_0000_0000_0000;
array[29032] <= 16'b0000_0000_0000_0000;
array[29033] <= 16'b0000_0000_0000_0000;
array[29034] <= 16'b0000_0000_0000_0000;
array[29035] <= 16'b0000_0000_0000_0000;
array[29036] <= 16'b0000_0000_0000_0000;
array[29037] <= 16'b0000_0000_0000_0000;
array[29038] <= 16'b0000_0000_0000_0000;
array[29039] <= 16'b0000_0000_0000_0000;
array[29040] <= 16'b0000_0000_0000_0000;
array[29041] <= 16'b0000_0000_0000_0000;
array[29042] <= 16'b0000_0000_0000_0000;
array[29043] <= 16'b0000_0000_0000_0000;
array[29044] <= 16'b0000_0000_0000_0000;
array[29045] <= 16'b0000_0000_0000_0000;
array[29046] <= 16'b0000_0000_0000_0000;
array[29047] <= 16'b0000_0000_0000_0000;
array[29048] <= 16'b0000_0000_0000_0000;
array[29049] <= 16'b0000_0000_0000_0000;
array[29050] <= 16'b0000_0000_0000_0000;
array[29051] <= 16'b0000_0000_0000_0000;
array[29052] <= 16'b0000_0000_0000_0000;
array[29053] <= 16'b0000_0000_0000_0000;
array[29054] <= 16'b0000_0000_0000_0000;
array[29055] <= 16'b0000_0000_0000_0000;
array[29056] <= 16'b0000_0000_0000_0000;
array[29057] <= 16'b0000_0000_0000_0000;
array[29058] <= 16'b0000_0000_0000_0000;
array[29059] <= 16'b0000_0000_0000_0000;
array[29060] <= 16'b0000_0000_0000_0000;
array[29061] <= 16'b0000_0000_0000_0000;
array[29062] <= 16'b0000_0000_0000_0000;
array[29063] <= 16'b0000_0000_0000_0000;
array[29064] <= 16'b0000_0000_0000_0000;
array[29065] <= 16'b0000_0000_0000_0000;
array[29066] <= 16'b0000_0000_0000_0000;
array[29067] <= 16'b0000_0000_0000_0000;
array[29068] <= 16'b0000_0000_0000_0000;
array[29069] <= 16'b0000_0000_0000_0000;
array[29070] <= 16'b0000_0000_0000_0000;
array[29071] <= 16'b0000_0000_0000_0000;
array[29072] <= 16'b0000_0000_0000_0000;
array[29073] <= 16'b0000_0000_0000_0000;
array[29074] <= 16'b0000_0000_0000_0000;
array[29075] <= 16'b0000_0000_0000_0000;
array[29076] <= 16'b0000_0000_0000_0000;
array[29077] <= 16'b0000_0000_0000_0000;
array[29078] <= 16'b0000_0000_0000_0000;
array[29079] <= 16'b0000_0000_0000_0000;
array[29080] <= 16'b0000_0000_0000_0000;
array[29081] <= 16'b0000_0000_0000_0000;
array[29082] <= 16'b0000_0000_0000_0000;
array[29083] <= 16'b0000_0000_0000_0000;
array[29084] <= 16'b0000_0000_0000_0000;
array[29085] <= 16'b0000_0000_0000_0000;
array[29086] <= 16'b0000_0000_0000_0000;
array[29087] <= 16'b0000_0000_0000_0000;
array[29088] <= 16'b0000_0000_0000_0000;
array[29089] <= 16'b0000_0000_0000_0000;
array[29090] <= 16'b0000_0000_0000_0000;
array[29091] <= 16'b0000_0000_0000_0000;
array[29092] <= 16'b0000_0000_0000_0000;
array[29093] <= 16'b0000_0000_0000_0000;
array[29094] <= 16'b0000_0000_0000_0000;
array[29095] <= 16'b0000_0000_0000_0000;
array[29096] <= 16'b0000_0000_0000_0000;
array[29097] <= 16'b0000_0000_0000_0000;
array[29098] <= 16'b0000_0000_0000_0000;
array[29099] <= 16'b0000_0000_0000_0000;
array[29100] <= 16'b0000_0000_0000_0000;
array[29101] <= 16'b0000_0000_0000_0000;
array[29102] <= 16'b0000_0000_0000_0000;
array[29103] <= 16'b0000_0000_0000_0000;
array[29104] <= 16'b0000_0000_0000_0000;
array[29105] <= 16'b0000_0000_0000_0000;
array[29106] <= 16'b0000_0000_0000_0000;
array[29107] <= 16'b0000_0000_0000_0000;
array[29108] <= 16'b0000_0000_0000_0000;
array[29109] <= 16'b0000_0000_0000_0000;
array[29110] <= 16'b0000_0000_0000_0000;
array[29111] <= 16'b0000_0000_0000_0000;
array[29112] <= 16'b0000_0000_0000_0000;
array[29113] <= 16'b0000_0000_0000_0000;
array[29114] <= 16'b0000_0000_0000_0000;
array[29115] <= 16'b0000_0000_0000_0000;
array[29116] <= 16'b0000_0000_0000_0000;
array[29117] <= 16'b0000_0000_0000_0000;
array[29118] <= 16'b0000_0000_0000_0000;
array[29119] <= 16'b0000_0000_0000_0000;
array[29120] <= 16'b0000_0000_0000_0000;
array[29121] <= 16'b0000_0000_0000_0000;
array[29122] <= 16'b0000_0000_0000_0000;
array[29123] <= 16'b0000_0000_0000_0000;
array[29124] <= 16'b0000_0000_0000_0000;
array[29125] <= 16'b0000_0000_0000_0000;
array[29126] <= 16'b0000_0000_0000_0000;
array[29127] <= 16'b0000_0000_0000_0000;
array[29128] <= 16'b0000_0000_0000_0000;
array[29129] <= 16'b0000_0000_0000_0000;
array[29130] <= 16'b0000_0000_0000_0000;
array[29131] <= 16'b0000_0000_0000_0000;
array[29132] <= 16'b0000_0000_0000_0000;
array[29133] <= 16'b0000_0000_0000_0000;
array[29134] <= 16'b0000_0000_0000_0000;
array[29135] <= 16'b0000_0000_0000_0000;
array[29136] <= 16'b0000_0000_0000_0000;
array[29137] <= 16'b0000_0000_0000_0000;
array[29138] <= 16'b0000_0000_0000_0000;
array[29139] <= 16'b0000_0000_0000_0000;
array[29140] <= 16'b0000_0000_0000_0000;
array[29141] <= 16'b0000_0000_0000_0000;
array[29142] <= 16'b0000_0000_0000_0000;
array[29143] <= 16'b0000_0000_0000_0000;
array[29144] <= 16'b0000_0000_0000_0000;
array[29145] <= 16'b0000_0000_0000_0000;
array[29146] <= 16'b0000_0000_0000_0000;
array[29147] <= 16'b0000_0000_0000_0000;
array[29148] <= 16'b0000_0000_0000_0000;
array[29149] <= 16'b0000_0000_0000_0000;
array[29150] <= 16'b0000_0000_0000_0000;
array[29151] <= 16'b0000_0000_0000_0000;
array[29152] <= 16'b0000_0000_0000_0000;
array[29153] <= 16'b0000_0000_0000_0000;
array[29154] <= 16'b0000_0000_0000_0000;
array[29155] <= 16'b0000_0000_0000_0000;
array[29156] <= 16'b0000_0000_0000_0000;
array[29157] <= 16'b0000_0000_0000_0000;
array[29158] <= 16'b0000_0000_0000_0000;
array[29159] <= 16'b0000_0000_0000_0000;
array[29160] <= 16'b0000_0000_0000_0000;
array[29161] <= 16'b0000_0000_0000_0000;
array[29162] <= 16'b0000_0000_0000_0000;
array[29163] <= 16'b0000_0000_0000_0000;
array[29164] <= 16'b0000_0000_0000_0000;
array[29165] <= 16'b0000_0000_0000_0000;
array[29166] <= 16'b0000_0000_0000_0000;
array[29167] <= 16'b0000_0000_0000_0000;
array[29168] <= 16'b0000_0000_0000_0000;
array[29169] <= 16'b0000_0000_0000_0000;
array[29170] <= 16'b0000_0000_0000_0000;
array[29171] <= 16'b0000_0000_0000_0000;
array[29172] <= 16'b0000_0000_0000_0000;
array[29173] <= 16'b0000_0000_0000_0000;
array[29174] <= 16'b0000_0000_0000_0000;
array[29175] <= 16'b0000_0000_0000_0000;
array[29176] <= 16'b0000_0000_0000_0000;
array[29177] <= 16'b0000_0000_0000_0000;
array[29178] <= 16'b0000_0000_0000_0000;
array[29179] <= 16'b0000_0000_0000_0000;
array[29180] <= 16'b0000_0000_0000_0000;
array[29181] <= 16'b0000_0000_0000_0000;
array[29182] <= 16'b0000_0000_0000_0000;
array[29183] <= 16'b0000_0000_0000_0000;
array[29184] <= 16'b0000_0000_0000_0000;
array[29185] <= 16'b0000_0000_0000_0000;
array[29186] <= 16'b0000_0000_0000_0000;
array[29187] <= 16'b0000_0000_0000_0000;
array[29188] <= 16'b0000_0000_0000_0000;
array[29189] <= 16'b0000_0000_0000_0000;
array[29190] <= 16'b0000_0000_0000_0000;
array[29191] <= 16'b0000_0000_0000_0000;
array[29192] <= 16'b0000_0000_0000_0000;
array[29193] <= 16'b0000_0000_0000_0000;
array[29194] <= 16'b0000_0000_0000_0000;
array[29195] <= 16'b0000_0000_0000_0000;
array[29196] <= 16'b0000_0000_0000_0000;
array[29197] <= 16'b0000_0000_0000_0000;
array[29198] <= 16'b0000_0000_0000_0000;
array[29199] <= 16'b0000_0000_0000_0000;
array[29200] <= 16'b0000_0000_0000_0000;
array[29201] <= 16'b0000_0000_0000_0000;
array[29202] <= 16'b0000_0000_0000_0000;
array[29203] <= 16'b0000_0000_0000_0000;
array[29204] <= 16'b0000_0000_0000_0000;
array[29205] <= 16'b0000_0000_0000_0000;
array[29206] <= 16'b0000_0000_0000_0000;
array[29207] <= 16'b0000_0000_0000_0000;
array[29208] <= 16'b0000_0000_0000_0000;
array[29209] <= 16'b0000_0000_0000_0000;
array[29210] <= 16'b0000_0000_0000_0000;
array[29211] <= 16'b0000_0000_0000_0000;
array[29212] <= 16'b0000_0000_0000_0000;
array[29213] <= 16'b0000_0000_0000_0000;
array[29214] <= 16'b0000_0000_0000_0000;
array[29215] <= 16'b0000_0000_0000_0000;
array[29216] <= 16'b0000_0000_0000_0000;
array[29217] <= 16'b0000_0000_0000_0000;
array[29218] <= 16'b0000_0000_0000_0000;
array[29219] <= 16'b0000_0000_0000_0000;
array[29220] <= 16'b0000_0000_0000_0000;
array[29221] <= 16'b0000_0000_0000_0000;
array[29222] <= 16'b0000_0000_0000_0000;
array[29223] <= 16'b0000_0000_0000_0000;
array[29224] <= 16'b0000_0000_0000_0000;
array[29225] <= 16'b0000_0000_0000_0000;
array[29226] <= 16'b0000_0000_0000_0000;
array[29227] <= 16'b0000_0000_0000_0000;
array[29228] <= 16'b0000_0000_0000_0000;
array[29229] <= 16'b0000_0000_0000_0000;
array[29230] <= 16'b0000_0000_0000_0000;
array[29231] <= 16'b0000_0000_0000_0000;
array[29232] <= 16'b0000_0000_0000_0000;
array[29233] <= 16'b0000_0000_0000_0000;
array[29234] <= 16'b0000_0000_0000_0000;
array[29235] <= 16'b0000_0000_0000_0000;
array[29236] <= 16'b0000_0000_0000_0000;
array[29237] <= 16'b0000_0000_0000_0000;
array[29238] <= 16'b0000_0000_0000_0000;
array[29239] <= 16'b0000_0000_0000_0000;
array[29240] <= 16'b0000_0000_0000_0000;
array[29241] <= 16'b0000_0000_0000_0000;
array[29242] <= 16'b0000_0000_0000_0000;
array[29243] <= 16'b0000_0000_0000_0000;
array[29244] <= 16'b0000_0000_0000_0000;
array[29245] <= 16'b0000_0000_0000_0000;
array[29246] <= 16'b0000_0000_0000_0000;
array[29247] <= 16'b0000_0000_0000_0000;
array[29248] <= 16'b0000_0000_0000_0000;
array[29249] <= 16'b0000_0000_0000_0000;
array[29250] <= 16'b0000_0000_0000_0000;
array[29251] <= 16'b0000_0000_0000_0000;
array[29252] <= 16'b0000_0000_0000_0000;
array[29253] <= 16'b0000_0000_0000_0000;
array[29254] <= 16'b0000_0000_0000_0000;
array[29255] <= 16'b0000_0000_0000_0000;
array[29256] <= 16'b0000_0000_0000_0000;
array[29257] <= 16'b0000_0000_0000_0000;
array[29258] <= 16'b0000_0000_0000_0000;
array[29259] <= 16'b0000_0000_0000_0000;
array[29260] <= 16'b0000_0000_0000_0000;
array[29261] <= 16'b0000_0000_0000_0000;
array[29262] <= 16'b0000_0000_0000_0000;
array[29263] <= 16'b0000_0000_0000_0000;
array[29264] <= 16'b0000_0000_0000_0000;
array[29265] <= 16'b0000_0000_0000_0000;
array[29266] <= 16'b0000_0000_0000_0000;
array[29267] <= 16'b0000_0000_0000_0000;
array[29268] <= 16'b0000_0000_0000_0000;
array[29269] <= 16'b0000_0000_0000_0000;
array[29270] <= 16'b0000_0000_0000_0000;
array[29271] <= 16'b0000_0000_0000_0000;
array[29272] <= 16'b0000_0000_0000_0000;
array[29273] <= 16'b0000_0000_0000_0000;
array[29274] <= 16'b0000_0000_0000_0000;
array[29275] <= 16'b0000_0000_0000_0000;
array[29276] <= 16'b0000_0000_0000_0000;
array[29277] <= 16'b0000_0000_0000_0000;
array[29278] <= 16'b0000_0000_0000_0000;
array[29279] <= 16'b0000_0000_0000_0000;
array[29280] <= 16'b0000_0000_0000_0000;
array[29281] <= 16'b0000_0000_0000_0000;
array[29282] <= 16'b0000_0000_0000_0000;
array[29283] <= 16'b0000_0000_0000_0000;
array[29284] <= 16'b0000_0000_0000_0000;
array[29285] <= 16'b0000_0000_0000_0000;
array[29286] <= 16'b0000_0000_0000_0000;
array[29287] <= 16'b0000_0000_0000_0000;
array[29288] <= 16'b0000_0000_0000_0000;
array[29289] <= 16'b0000_0000_0000_0000;
array[29290] <= 16'b0000_0000_0000_0000;
array[29291] <= 16'b0000_0000_0000_0000;
array[29292] <= 16'b0000_0000_0000_0000;
array[29293] <= 16'b0000_0000_0000_0000;
array[29294] <= 16'b0000_0000_0000_0000;
array[29295] <= 16'b0000_0000_0000_0000;
array[29296] <= 16'b0000_0000_0000_0000;
array[29297] <= 16'b0000_0000_0000_0000;
array[29298] <= 16'b0000_0000_0000_0000;
array[29299] <= 16'b0000_0000_0000_0000;
array[29300] <= 16'b0000_0000_0000_0000;
array[29301] <= 16'b0000_0000_0000_0000;
array[29302] <= 16'b0000_0000_0000_0000;
array[29303] <= 16'b0000_0000_0000_0000;
array[29304] <= 16'b0000_0000_0000_0000;
array[29305] <= 16'b0000_0000_0000_0000;
array[29306] <= 16'b0000_0000_0000_0000;
array[29307] <= 16'b0000_0000_0000_0000;
array[29308] <= 16'b0000_0000_0000_0000;
array[29309] <= 16'b0000_0000_0000_0000;
array[29310] <= 16'b0000_0000_0000_0000;
array[29311] <= 16'b0000_0000_0000_0000;
array[29312] <= 16'b0000_0000_0000_0000;
array[29313] <= 16'b0000_0000_0000_0000;
array[29314] <= 16'b0000_0000_0000_0000;
array[29315] <= 16'b0000_0000_0000_0000;
array[29316] <= 16'b0000_0000_0000_0000;
array[29317] <= 16'b0000_0000_0000_0000;
array[29318] <= 16'b0000_0000_0000_0000;
array[29319] <= 16'b0000_0000_0000_0000;
array[29320] <= 16'b0000_0000_0000_0000;
array[29321] <= 16'b0000_0000_0000_0000;
array[29322] <= 16'b0000_0000_0000_0000;
array[29323] <= 16'b0000_0000_0000_0000;
array[29324] <= 16'b0000_0000_0000_0000;
array[29325] <= 16'b0000_0000_0000_0000;
array[29326] <= 16'b0000_0000_0000_0000;
array[29327] <= 16'b0000_0000_0000_0000;
array[29328] <= 16'b0000_0000_0000_0000;
array[29329] <= 16'b0000_0000_0000_0000;
array[29330] <= 16'b0000_0000_0000_0000;
array[29331] <= 16'b0000_0000_0000_0000;
array[29332] <= 16'b0000_0000_0000_0000;
array[29333] <= 16'b0000_0000_0000_0000;
array[29334] <= 16'b0000_0000_0000_0000;
array[29335] <= 16'b0000_0000_0000_0000;
array[29336] <= 16'b0000_0000_0000_0000;
array[29337] <= 16'b0000_0000_0000_0000;
array[29338] <= 16'b0000_0000_0000_0000;
array[29339] <= 16'b0000_0000_0000_0000;
array[29340] <= 16'b0000_0000_0000_0000;
array[29341] <= 16'b0000_0000_0000_0000;
array[29342] <= 16'b0000_0000_0000_0000;
array[29343] <= 16'b0000_0000_0000_0000;
array[29344] <= 16'b0000_0000_0000_0000;
array[29345] <= 16'b0000_0000_0000_0000;
array[29346] <= 16'b0000_0000_0000_0000;
array[29347] <= 16'b0000_0000_0000_0000;
array[29348] <= 16'b0000_0000_0000_0000;
array[29349] <= 16'b0000_0000_0000_0000;
array[29350] <= 16'b0000_0000_0000_0000;
array[29351] <= 16'b0000_0000_0000_0000;
array[29352] <= 16'b0000_0000_0000_0000;
array[29353] <= 16'b0000_0000_0000_0000;
array[29354] <= 16'b0000_0000_0000_0000;
array[29355] <= 16'b0000_0000_0000_0000;
array[29356] <= 16'b0000_0000_0000_0000;
array[29357] <= 16'b0000_0000_0000_0000;
array[29358] <= 16'b0000_0000_0000_0000;
array[29359] <= 16'b0000_0000_0000_0000;
array[29360] <= 16'b0000_0000_0000_0000;
array[29361] <= 16'b0000_0000_0000_0000;
array[29362] <= 16'b0000_0000_0000_0000;
array[29363] <= 16'b0000_0000_0000_0000;
array[29364] <= 16'b0000_0000_0000_0000;
array[29365] <= 16'b0000_0000_0000_0000;
array[29366] <= 16'b0000_0000_0000_0000;
array[29367] <= 16'b0000_0000_0000_0000;
array[29368] <= 16'b0000_0000_0000_0000;
array[29369] <= 16'b0000_0000_0000_0000;
array[29370] <= 16'b0000_0000_0000_0000;
array[29371] <= 16'b0000_0000_0000_0000;
array[29372] <= 16'b0000_0000_0000_0000;
array[29373] <= 16'b0000_0000_0000_0000;
array[29374] <= 16'b0000_0000_0000_0000;
array[29375] <= 16'b0000_0000_0000_0000;
array[29376] <= 16'b0000_0000_0000_0000;
array[29377] <= 16'b0000_0000_0000_0000;
array[29378] <= 16'b0000_0000_0000_0000;
array[29379] <= 16'b0000_0000_0000_0000;
array[29380] <= 16'b0000_0000_0000_0000;
array[29381] <= 16'b0000_0000_0000_0000;
array[29382] <= 16'b0000_0000_0000_0000;
array[29383] <= 16'b0000_0000_0000_0000;
array[29384] <= 16'b0000_0000_0000_0000;
array[29385] <= 16'b0000_0000_0000_0000;
array[29386] <= 16'b0000_0000_0000_0000;
array[29387] <= 16'b0000_0000_0000_0000;
array[29388] <= 16'b0000_0000_0000_0000;
array[29389] <= 16'b0000_0000_0000_0000;
array[29390] <= 16'b0000_0000_0000_0000;
array[29391] <= 16'b0000_0000_0000_0000;
array[29392] <= 16'b0000_0000_0000_0000;
array[29393] <= 16'b0000_0000_0000_0000;
array[29394] <= 16'b0000_0000_0000_0000;
array[29395] <= 16'b0000_0000_0000_0000;
array[29396] <= 16'b0000_0000_0000_0000;
array[29397] <= 16'b0000_0000_0000_0000;
array[29398] <= 16'b0000_0000_0000_0000;
array[29399] <= 16'b0000_0000_0000_0000;
array[29400] <= 16'b0000_0000_0000_0000;
array[29401] <= 16'b0000_0000_0000_0000;
array[29402] <= 16'b0000_0000_0000_0000;
array[29403] <= 16'b0000_0000_0000_0000;
array[29404] <= 16'b0000_0000_0000_0000;
array[29405] <= 16'b0000_0000_0000_0000;
array[29406] <= 16'b0000_0000_0000_0000;
array[29407] <= 16'b0000_0000_0000_0000;
array[29408] <= 16'b0000_0000_0000_0000;
array[29409] <= 16'b0000_0000_0000_0000;
array[29410] <= 16'b0000_0000_0000_0000;
array[29411] <= 16'b0000_0000_0000_0000;
array[29412] <= 16'b0000_0000_0000_0000;
array[29413] <= 16'b0000_0000_0000_0000;
array[29414] <= 16'b0000_0000_0000_0000;
array[29415] <= 16'b0000_0000_0000_0000;
array[29416] <= 16'b0000_0000_0000_0000;
array[29417] <= 16'b0000_0000_0000_0000;
array[29418] <= 16'b0000_0000_0000_0000;
array[29419] <= 16'b0000_0000_0000_0000;
array[29420] <= 16'b0000_0000_0000_0000;
array[29421] <= 16'b0000_0000_0000_0000;
array[29422] <= 16'b0000_0000_0000_0000;
array[29423] <= 16'b0000_0000_0000_0000;
array[29424] <= 16'b0000_0000_0000_0000;
array[29425] <= 16'b0000_0000_0000_0000;
array[29426] <= 16'b0000_0000_0000_0000;
array[29427] <= 16'b0000_0000_0000_0000;
array[29428] <= 16'b0000_0000_0000_0000;
array[29429] <= 16'b0000_0000_0000_0000;
array[29430] <= 16'b0000_0000_0000_0000;
array[29431] <= 16'b0000_0000_0000_0000;
array[29432] <= 16'b0000_0000_0000_0000;
array[29433] <= 16'b0000_0000_0000_0000;
array[29434] <= 16'b0000_0000_0000_0000;
array[29435] <= 16'b0000_0000_0000_0000;
array[29436] <= 16'b0000_0000_0000_0000;
array[29437] <= 16'b0000_0000_0000_0000;
array[29438] <= 16'b0000_0000_0000_0000;
array[29439] <= 16'b0000_0000_0000_0000;
array[29440] <= 16'b0000_0000_0000_0000;
array[29441] <= 16'b0000_0000_0000_0000;
array[29442] <= 16'b0000_0000_0000_0000;
array[29443] <= 16'b0000_0000_0000_0000;
array[29444] <= 16'b0000_0000_0000_0000;
array[29445] <= 16'b0000_0000_0000_0000;
array[29446] <= 16'b0000_0000_0000_0000;
array[29447] <= 16'b0000_0000_0000_0000;
array[29448] <= 16'b0000_0000_0000_0000;
array[29449] <= 16'b0000_0000_0000_0000;
array[29450] <= 16'b0000_0000_0000_0000;
array[29451] <= 16'b0000_0000_0000_0000;
array[29452] <= 16'b0000_0000_0000_0000;
array[29453] <= 16'b0000_0000_0000_0000;
array[29454] <= 16'b0000_0000_0000_0000;
array[29455] <= 16'b0000_0000_0000_0000;
array[29456] <= 16'b0000_0000_0000_0000;
array[29457] <= 16'b0000_0000_0000_0000;
array[29458] <= 16'b0000_0000_0000_0000;
array[29459] <= 16'b0000_0000_0000_0000;
array[29460] <= 16'b0000_0000_0000_0000;
array[29461] <= 16'b0000_0000_0000_0000;
array[29462] <= 16'b0000_0000_0000_0000;
array[29463] <= 16'b0000_0000_0000_0000;
array[29464] <= 16'b0000_0000_0000_0000;
array[29465] <= 16'b0000_0000_0000_0000;
array[29466] <= 16'b0000_0000_0000_0000;
array[29467] <= 16'b0000_0000_0000_0000;
array[29468] <= 16'b0000_0000_0000_0000;
array[29469] <= 16'b0000_0000_0000_0000;
array[29470] <= 16'b0000_0000_0000_0000;
array[29471] <= 16'b0000_0000_0000_0000;
array[29472] <= 16'b0000_0000_0000_0000;
array[29473] <= 16'b0000_0000_0000_0000;
array[29474] <= 16'b0000_0000_0000_0000;
array[29475] <= 16'b0000_0000_0000_0000;
array[29476] <= 16'b0000_0000_0000_0000;
array[29477] <= 16'b0000_0000_0000_0000;
array[29478] <= 16'b0000_0000_0000_0000;
array[29479] <= 16'b0000_0000_0000_0000;
array[29480] <= 16'b0000_0000_0000_0000;
array[29481] <= 16'b0000_0000_0000_0000;
array[29482] <= 16'b0000_0000_0000_0000;
array[29483] <= 16'b0000_0000_0000_0000;
array[29484] <= 16'b0000_0000_0000_0000;
array[29485] <= 16'b0000_0000_0000_0000;
array[29486] <= 16'b0000_0000_0000_0000;
array[29487] <= 16'b0000_0000_0000_0000;
array[29488] <= 16'b0000_0000_0000_0000;
array[29489] <= 16'b0000_0000_0000_0000;
array[29490] <= 16'b0000_0000_0000_0000;
array[29491] <= 16'b0000_0000_0000_0000;
array[29492] <= 16'b0000_0000_0000_0000;
array[29493] <= 16'b0000_0000_0000_0000;
array[29494] <= 16'b0000_0000_0000_0000;
array[29495] <= 16'b0000_0000_0000_0000;
array[29496] <= 16'b0000_0000_0000_0000;
array[29497] <= 16'b0000_0000_0000_0000;
array[29498] <= 16'b0000_0000_0000_0000;
array[29499] <= 16'b0000_0000_0000_0000;
array[29500] <= 16'b0000_0000_0000_0000;
array[29501] <= 16'b0000_0000_0000_0000;
array[29502] <= 16'b0000_0000_0000_0000;
array[29503] <= 16'b0000_0000_0000_0000;
array[29504] <= 16'b0000_0000_0000_0000;
array[29505] <= 16'b0000_0000_0000_0000;
array[29506] <= 16'b0000_0000_0000_0000;
array[29507] <= 16'b0000_0000_0000_0000;
array[29508] <= 16'b0000_0000_0000_0000;
array[29509] <= 16'b0000_0000_0000_0000;
array[29510] <= 16'b0000_0000_0000_0000;
array[29511] <= 16'b0000_0000_0000_0000;
array[29512] <= 16'b0000_0000_0000_0000;
array[29513] <= 16'b0000_0000_0000_0000;
array[29514] <= 16'b0000_0000_0000_0000;
array[29515] <= 16'b0000_0000_0000_0000;
array[29516] <= 16'b0000_0000_0000_0000;
array[29517] <= 16'b0000_0000_0000_0000;
array[29518] <= 16'b0000_0000_0000_0000;
array[29519] <= 16'b0000_0000_0000_0000;
array[29520] <= 16'b0000_0000_0000_0000;
array[29521] <= 16'b0000_0000_0000_0000;
array[29522] <= 16'b0000_0000_0000_0000;
array[29523] <= 16'b0000_0000_0000_0000;
array[29524] <= 16'b0000_0000_0000_0000;
array[29525] <= 16'b0000_0000_0000_0000;
array[29526] <= 16'b0000_0000_0000_0000;
array[29527] <= 16'b0000_0000_0000_0000;
array[29528] <= 16'b0000_0000_0000_0000;
array[29529] <= 16'b0000_0000_0000_0000;
array[29530] <= 16'b0000_0000_0000_0000;
array[29531] <= 16'b0000_0000_0000_0000;
array[29532] <= 16'b0000_0000_0000_0000;
array[29533] <= 16'b0000_0000_0000_0000;
array[29534] <= 16'b0000_0000_0000_0000;
array[29535] <= 16'b0000_0000_0000_0000;
array[29536] <= 16'b0000_0000_0000_0000;
array[29537] <= 16'b0000_0000_0000_0000;
array[29538] <= 16'b0000_0000_0000_0000;
array[29539] <= 16'b0000_0000_0000_0000;
array[29540] <= 16'b0000_0000_0000_0000;
array[29541] <= 16'b0000_0000_0000_0000;
array[29542] <= 16'b0000_0000_0000_0000;
array[29543] <= 16'b0000_0000_0000_0000;
array[29544] <= 16'b0000_0000_0000_0000;
array[29545] <= 16'b0000_0000_0000_0000;
array[29546] <= 16'b0000_0000_0000_0000;
array[29547] <= 16'b0000_0000_0000_0000;
array[29548] <= 16'b0000_0000_0000_0000;
array[29549] <= 16'b0000_0000_0000_0000;
array[29550] <= 16'b0000_0000_0000_0000;
array[29551] <= 16'b0000_0000_0000_0000;
array[29552] <= 16'b0000_0000_0000_0000;
array[29553] <= 16'b0000_0000_0000_0000;
array[29554] <= 16'b0000_0000_0000_0000;
array[29555] <= 16'b0000_0000_0000_0000;
array[29556] <= 16'b0000_0000_0000_0000;
array[29557] <= 16'b0000_0000_0000_0000;
array[29558] <= 16'b0000_0000_0000_0000;
array[29559] <= 16'b0000_0000_0000_0000;
array[29560] <= 16'b0000_0000_0000_0000;
array[29561] <= 16'b0000_0000_0000_0000;
array[29562] <= 16'b0000_0000_0000_0000;
array[29563] <= 16'b0000_0000_0000_0000;
array[29564] <= 16'b0000_0000_0000_0000;
array[29565] <= 16'b0000_0000_0000_0000;
array[29566] <= 16'b0000_0000_0000_0000;
array[29567] <= 16'b0000_0000_0000_0000;
array[29568] <= 16'b0000_0000_0000_0000;
array[29569] <= 16'b0000_0000_0000_0000;
array[29570] <= 16'b0000_0000_0000_0000;
array[29571] <= 16'b0000_0000_0000_0000;
array[29572] <= 16'b0000_0000_0000_0000;
array[29573] <= 16'b0000_0000_0000_0000;
array[29574] <= 16'b0000_0000_0000_0000;
array[29575] <= 16'b0000_0000_0000_0000;
array[29576] <= 16'b0000_0000_0000_0000;
array[29577] <= 16'b0000_0000_0000_0000;
array[29578] <= 16'b0000_0000_0000_0000;
array[29579] <= 16'b0000_0000_0000_0000;
array[29580] <= 16'b0000_0000_0000_0000;
array[29581] <= 16'b0000_0000_0000_0000;
array[29582] <= 16'b0000_0000_0000_0000;
array[29583] <= 16'b0000_0000_0000_0000;
array[29584] <= 16'b0000_0000_0000_0000;
array[29585] <= 16'b0000_0000_0000_0000;
array[29586] <= 16'b0000_0000_0000_0000;
array[29587] <= 16'b0000_0000_0000_0000;
array[29588] <= 16'b0000_0000_0000_0000;
array[29589] <= 16'b0000_0000_0000_0000;
array[29590] <= 16'b0000_0000_0000_0000;
array[29591] <= 16'b0000_0000_0000_0000;
array[29592] <= 16'b0000_0000_0000_0000;
array[29593] <= 16'b0000_0000_0000_0000;
array[29594] <= 16'b0000_0000_0000_0000;
array[29595] <= 16'b0000_0000_0000_0000;
array[29596] <= 16'b0000_0000_0000_0000;
array[29597] <= 16'b0000_0000_0000_0000;
array[29598] <= 16'b0000_0000_0000_0000;
array[29599] <= 16'b0000_0000_0000_0000;
array[29600] <= 16'b0000_0000_0000_0000;
array[29601] <= 16'b0000_0000_0000_0000;
array[29602] <= 16'b0000_0000_0000_0000;
array[29603] <= 16'b0000_0000_0000_0000;
array[29604] <= 16'b0000_0000_0000_0000;
array[29605] <= 16'b0000_0000_0000_0000;
array[29606] <= 16'b0000_0000_0000_0000;
array[29607] <= 16'b0000_0000_0000_0000;
array[29608] <= 16'b0000_0000_0000_0000;
array[29609] <= 16'b0000_0000_0000_0000;
array[29610] <= 16'b0000_0000_0000_0000;
array[29611] <= 16'b0000_0000_0000_0000;
array[29612] <= 16'b0000_0000_0000_0000;
array[29613] <= 16'b0000_0000_0000_0000;
array[29614] <= 16'b0000_0000_0000_0000;
array[29615] <= 16'b0000_0000_0000_0000;
array[29616] <= 16'b0000_0000_0000_0000;
array[29617] <= 16'b0000_0000_0000_0000;
array[29618] <= 16'b0000_0000_0000_0000;
array[29619] <= 16'b0000_0000_0000_0000;
array[29620] <= 16'b0000_0000_0000_0000;
array[29621] <= 16'b0000_0000_0000_0000;
array[29622] <= 16'b0000_0000_0000_0000;
array[29623] <= 16'b0000_0000_0000_0000;
array[29624] <= 16'b0000_0000_0000_0000;
array[29625] <= 16'b0000_0000_0000_0000;
array[29626] <= 16'b0000_0000_0000_0000;
array[29627] <= 16'b0000_0000_0000_0000;
array[29628] <= 16'b0000_0000_0000_0000;
array[29629] <= 16'b0000_0000_0000_0000;
array[29630] <= 16'b0000_0000_0000_0000;
array[29631] <= 16'b0000_0000_0000_0000;
array[29632] <= 16'b0000_0000_0000_0000;
array[29633] <= 16'b0000_0000_0000_0000;
array[29634] <= 16'b0000_0000_0000_0000;
array[29635] <= 16'b0000_0000_0000_0000;
array[29636] <= 16'b0000_0000_0000_0000;
array[29637] <= 16'b0000_0000_0000_0000;
array[29638] <= 16'b0000_0000_0000_0000;
array[29639] <= 16'b0000_0000_0000_0000;
array[29640] <= 16'b0000_0000_0000_0000;
array[29641] <= 16'b0000_0000_0000_0000;
array[29642] <= 16'b0000_0000_0000_0000;
array[29643] <= 16'b0000_0000_0000_0000;
array[29644] <= 16'b0000_0000_0000_0000;
array[29645] <= 16'b0000_0000_0000_0000;
array[29646] <= 16'b0000_0000_0000_0000;
array[29647] <= 16'b0000_0000_0000_0000;
array[29648] <= 16'b0000_0000_0000_0000;
array[29649] <= 16'b0000_0000_0000_0000;
array[29650] <= 16'b0000_0000_0000_0000;
array[29651] <= 16'b0000_0000_0000_0000;
array[29652] <= 16'b0000_0000_0000_0000;
array[29653] <= 16'b0000_0000_0000_0000;
array[29654] <= 16'b0000_0000_0000_0000;
array[29655] <= 16'b0000_0000_0000_0000;
array[29656] <= 16'b0000_0000_0000_0000;
array[29657] <= 16'b0000_0000_0000_0000;
array[29658] <= 16'b0000_0000_0000_0000;
array[29659] <= 16'b0000_0000_0000_0000;
array[29660] <= 16'b0000_0000_0000_0000;
array[29661] <= 16'b0000_0000_0000_0000;
array[29662] <= 16'b0000_0000_0000_0000;
array[29663] <= 16'b0000_0000_0000_0000;
array[29664] <= 16'b0000_0000_0000_0000;
array[29665] <= 16'b0000_0000_0000_0000;
array[29666] <= 16'b0000_0000_0000_0000;
array[29667] <= 16'b0000_0000_0000_0000;
array[29668] <= 16'b0000_0000_0000_0000;
array[29669] <= 16'b0000_0000_0000_0000;
array[29670] <= 16'b0000_0000_0000_0000;
array[29671] <= 16'b0000_0000_0000_0000;
array[29672] <= 16'b0000_0000_0000_0000;
array[29673] <= 16'b0000_0000_0000_0000;
array[29674] <= 16'b0000_0000_0000_0000;
array[29675] <= 16'b0000_0000_0000_0000;
array[29676] <= 16'b0000_0000_0000_0000;
array[29677] <= 16'b0000_0000_0000_0000;
array[29678] <= 16'b0000_0000_0000_0000;
array[29679] <= 16'b0000_0000_0000_0000;
array[29680] <= 16'b0000_0000_0000_0000;
array[29681] <= 16'b0000_0000_0000_0000;
array[29682] <= 16'b0000_0000_0000_0000;
array[29683] <= 16'b0000_0000_0000_0000;
array[29684] <= 16'b0000_0000_0000_0000;
array[29685] <= 16'b0000_0000_0000_0000;
array[29686] <= 16'b0000_0000_0000_0000;
array[29687] <= 16'b0000_0000_0000_0000;
array[29688] <= 16'b0000_0000_0000_0000;
array[29689] <= 16'b0000_0000_0000_0000;
array[29690] <= 16'b0000_0000_0000_0000;
array[29691] <= 16'b0000_0000_0000_0000;
array[29692] <= 16'b0000_0000_0000_0000;
array[29693] <= 16'b0000_0000_0000_0000;
array[29694] <= 16'b0000_0000_0000_0000;
array[29695] <= 16'b0000_0000_0000_0000;
array[29696] <= 16'b0000_0000_0000_0000;
array[29697] <= 16'b0000_0000_0000_0000;
array[29698] <= 16'b0000_0000_0000_0000;
array[29699] <= 16'b0000_0000_0000_0000;
array[29700] <= 16'b0000_0000_0000_0000;
array[29701] <= 16'b0000_0000_0000_0000;
array[29702] <= 16'b0000_0000_0000_0000;
array[29703] <= 16'b0000_0000_0000_0000;
array[29704] <= 16'b0000_0000_0000_0000;
array[29705] <= 16'b0000_0000_0000_0000;
array[29706] <= 16'b0000_0000_0000_0000;
array[29707] <= 16'b0000_0000_0000_0000;
array[29708] <= 16'b0000_0000_0000_0000;
array[29709] <= 16'b0000_0000_0000_0000;
array[29710] <= 16'b0000_0000_0000_0000;
array[29711] <= 16'b0000_0000_0000_0000;
array[29712] <= 16'b0000_0000_0000_0000;
array[29713] <= 16'b0000_0000_0000_0000;
array[29714] <= 16'b0000_0000_0000_0000;
array[29715] <= 16'b0000_0000_0000_0000;
array[29716] <= 16'b0000_0000_0000_0000;
array[29717] <= 16'b0000_0000_0000_0000;
array[29718] <= 16'b0000_0000_0000_0000;
array[29719] <= 16'b0000_0000_0000_0000;
array[29720] <= 16'b0000_0000_0000_0000;
array[29721] <= 16'b0000_0000_0000_0000;
array[29722] <= 16'b0000_0000_0000_0000;
array[29723] <= 16'b0000_0000_0000_0000;
array[29724] <= 16'b0000_0000_0000_0000;
array[29725] <= 16'b0000_0000_0000_0000;
array[29726] <= 16'b0000_0000_0000_0000;
array[29727] <= 16'b0000_0000_0000_0000;
array[29728] <= 16'b0000_0000_0000_0000;
array[29729] <= 16'b0000_0000_0000_0000;
array[29730] <= 16'b0000_0000_0000_0000;
array[29731] <= 16'b0000_0000_0000_0000;
array[29732] <= 16'b0000_0000_0000_0000;
array[29733] <= 16'b0000_0000_0000_0000;
array[29734] <= 16'b0000_0000_0000_0000;
array[29735] <= 16'b0000_0000_0000_0000;
array[29736] <= 16'b0000_0000_0000_0000;
array[29737] <= 16'b0000_0000_0000_0000;
array[29738] <= 16'b0000_0000_0000_0000;
array[29739] <= 16'b0000_0000_0000_0000;
array[29740] <= 16'b0000_0000_0000_0000;
array[29741] <= 16'b0000_0000_0000_0000;
array[29742] <= 16'b0000_0000_0000_0000;
array[29743] <= 16'b0000_0000_0000_0000;
array[29744] <= 16'b0000_0000_0000_0000;
array[29745] <= 16'b0000_0000_0000_0000;
array[29746] <= 16'b0000_0000_0000_0000;
array[29747] <= 16'b0000_0000_0000_0000;
array[29748] <= 16'b0000_0000_0000_0000;
array[29749] <= 16'b0000_0000_0000_0000;
array[29750] <= 16'b0000_0000_0000_0000;
array[29751] <= 16'b0000_0000_0000_0000;
array[29752] <= 16'b0000_0000_0000_0000;
array[29753] <= 16'b0000_0000_0000_0000;
array[29754] <= 16'b0000_0000_0000_0000;
array[29755] <= 16'b0000_0000_0000_0000;
array[29756] <= 16'b0000_0000_0000_0000;
array[29757] <= 16'b0000_0000_0000_0000;
array[29758] <= 16'b0000_0000_0000_0000;
array[29759] <= 16'b0000_0000_0000_0000;
array[29760] <= 16'b0000_0000_0000_0000;
array[29761] <= 16'b0000_0000_0000_0000;
array[29762] <= 16'b0000_0000_0000_0000;
array[29763] <= 16'b0000_0000_0000_0000;
array[29764] <= 16'b0000_0000_0000_0000;
array[29765] <= 16'b0000_0000_0000_0000;
array[29766] <= 16'b0000_0000_0000_0000;
array[29767] <= 16'b0000_0000_0000_0000;
array[29768] <= 16'b0000_0000_0000_0000;
array[29769] <= 16'b0000_0000_0000_0000;
array[29770] <= 16'b0000_0000_0000_0000;
array[29771] <= 16'b0000_0000_0000_0000;
array[29772] <= 16'b0000_0000_0000_0000;
array[29773] <= 16'b0000_0000_0000_0000;
array[29774] <= 16'b0000_0000_0000_0000;
array[29775] <= 16'b0000_0000_0000_0000;
array[29776] <= 16'b0000_0000_0000_0000;
array[29777] <= 16'b0000_0000_0000_0000;
array[29778] <= 16'b0000_0000_0000_0000;
array[29779] <= 16'b0000_0000_0000_0000;
array[29780] <= 16'b0000_0000_0000_0000;
array[29781] <= 16'b0000_0000_0000_0000;
array[29782] <= 16'b0000_0000_0000_0000;
array[29783] <= 16'b0000_0000_0000_0000;
array[29784] <= 16'b0000_0000_0000_0000;
array[29785] <= 16'b0000_0000_0000_0000;
array[29786] <= 16'b0000_0000_0000_0000;
array[29787] <= 16'b0000_0000_0000_0000;
array[29788] <= 16'b0000_0000_0000_0000;
array[29789] <= 16'b0000_0000_0000_0000;
array[29790] <= 16'b0000_0000_0000_0000;
array[29791] <= 16'b0000_0000_0000_0000;
array[29792] <= 16'b0000_0000_0000_0000;
array[29793] <= 16'b0000_0000_0000_0000;
array[29794] <= 16'b0000_0000_0000_0000;
array[29795] <= 16'b0000_0000_0000_0000;
array[29796] <= 16'b0000_0000_0000_0000;
array[29797] <= 16'b0000_0000_0000_0000;
array[29798] <= 16'b0000_0000_0000_0000;
array[29799] <= 16'b0000_0000_0000_0000;
array[29800] <= 16'b0000_0000_0000_0000;
array[29801] <= 16'b0000_0000_0000_0000;
array[29802] <= 16'b0000_0000_0000_0000;
array[29803] <= 16'b0000_0000_0000_0000;
array[29804] <= 16'b0000_0000_0000_0000;
array[29805] <= 16'b0000_0000_0000_0000;
array[29806] <= 16'b0000_0000_0000_0000;
array[29807] <= 16'b0000_0000_0000_0000;
array[29808] <= 16'b0000_0000_0000_0000;
array[29809] <= 16'b0000_0000_0000_0000;
array[29810] <= 16'b0000_0000_0000_0000;
array[29811] <= 16'b0000_0000_0000_0000;
array[29812] <= 16'b0000_0000_0000_0000;
array[29813] <= 16'b0000_0000_0000_0000;
array[29814] <= 16'b0000_0000_0000_0000;
array[29815] <= 16'b0000_0000_0000_0000;
array[29816] <= 16'b0000_0000_0000_0000;
array[29817] <= 16'b0000_0000_0000_0000;
array[29818] <= 16'b0000_0000_0000_0000;
array[29819] <= 16'b0000_0000_0000_0000;
array[29820] <= 16'b0000_0000_0000_0000;
array[29821] <= 16'b0000_0000_0000_0000;
array[29822] <= 16'b0000_0000_0000_0000;
array[29823] <= 16'b0000_0000_0000_0000;
array[29824] <= 16'b0000_0000_0000_0000;
array[29825] <= 16'b0000_0000_0000_0000;
array[29826] <= 16'b0000_0000_0000_0000;
array[29827] <= 16'b0000_0000_0000_0000;
array[29828] <= 16'b0000_0000_0000_0000;
array[29829] <= 16'b0000_0000_0000_0000;
array[29830] <= 16'b0000_0000_0000_0000;
array[29831] <= 16'b0000_0000_0000_0000;
array[29832] <= 16'b0000_0000_0000_0000;
array[29833] <= 16'b0000_0000_0000_0000;
array[29834] <= 16'b0000_0000_0000_0000;
array[29835] <= 16'b0000_0000_0000_0000;
array[29836] <= 16'b0000_0000_0000_0000;
array[29837] <= 16'b0000_0000_0000_0000;
array[29838] <= 16'b0000_0000_0000_0000;
array[29839] <= 16'b0000_0000_0000_0000;
array[29840] <= 16'b0000_0000_0000_0000;
array[29841] <= 16'b0000_0000_0000_0000;
array[29842] <= 16'b0000_0000_0000_0000;
array[29843] <= 16'b0000_0000_0000_0000;
array[29844] <= 16'b0000_0000_0000_0000;
array[29845] <= 16'b0000_0000_0000_0000;
array[29846] <= 16'b0000_0000_0000_0000;
array[29847] <= 16'b0000_0000_0000_0000;
array[29848] <= 16'b0000_0000_0000_0000;
array[29849] <= 16'b0000_0000_0000_0000;
array[29850] <= 16'b0000_0000_0000_0000;
array[29851] <= 16'b0000_0000_0000_0000;
array[29852] <= 16'b0000_0000_0000_0000;
array[29853] <= 16'b0000_0000_0000_0000;
array[29854] <= 16'b0000_0000_0000_0000;
array[29855] <= 16'b0000_0000_0000_0000;
array[29856] <= 16'b0000_0000_0000_0000;
array[29857] <= 16'b0000_0000_0000_0000;
array[29858] <= 16'b0000_0000_0000_0000;
array[29859] <= 16'b0000_0000_0000_0000;
array[29860] <= 16'b0000_0000_0000_0000;
array[29861] <= 16'b0000_0000_0000_0000;
array[29862] <= 16'b0000_0000_0000_0000;
array[29863] <= 16'b0000_0000_0000_0000;
array[29864] <= 16'b0000_0000_0000_0000;
array[29865] <= 16'b0000_0000_0000_0000;
array[29866] <= 16'b0000_0000_0000_0000;
array[29867] <= 16'b0000_0000_0000_0000;
array[29868] <= 16'b0000_0000_0000_0000;
array[29869] <= 16'b0000_0000_0000_0000;
array[29870] <= 16'b0000_0000_0000_0000;
array[29871] <= 16'b0000_0000_0000_0000;
array[29872] <= 16'b0000_0000_0000_0000;
array[29873] <= 16'b0000_0000_0000_0000;
array[29874] <= 16'b0000_0000_0000_0000;
array[29875] <= 16'b0000_0000_0000_0000;
array[29876] <= 16'b0000_0000_0000_0000;
array[29877] <= 16'b0000_0000_0000_0000;
array[29878] <= 16'b0000_0000_0000_0000;
array[29879] <= 16'b0000_0000_0000_0000;
array[29880] <= 16'b0000_0000_0000_0000;
array[29881] <= 16'b0000_0000_0000_0000;
array[29882] <= 16'b0000_0000_0000_0000;
array[29883] <= 16'b0000_0000_0000_0000;
array[29884] <= 16'b0000_0000_0000_0000;
array[29885] <= 16'b0000_0000_0000_0000;
array[29886] <= 16'b0000_0000_0000_0000;
array[29887] <= 16'b0000_0000_0000_0000;
array[29888] <= 16'b0000_0000_0000_0000;
array[29889] <= 16'b0000_0000_0000_0000;
array[29890] <= 16'b0000_0000_0000_0000;
array[29891] <= 16'b0000_0000_0000_0000;
array[29892] <= 16'b0000_0000_0000_0000;
array[29893] <= 16'b0000_0000_0000_0000;
array[29894] <= 16'b0000_0000_0000_0000;
array[29895] <= 16'b0000_0000_0000_0000;
array[29896] <= 16'b0000_0000_0000_0000;
array[29897] <= 16'b0000_0000_0000_0000;
array[29898] <= 16'b0000_0000_0000_0000;
array[29899] <= 16'b0000_0000_0000_0000;
array[29900] <= 16'b0000_0000_0000_0000;
array[29901] <= 16'b0000_0000_0000_0000;
array[29902] <= 16'b0000_0000_0000_0000;
array[29903] <= 16'b0000_0000_0000_0000;
array[29904] <= 16'b0000_0000_0000_0000;
array[29905] <= 16'b0000_0000_0000_0000;
array[29906] <= 16'b0000_0000_0000_0000;
array[29907] <= 16'b0000_0000_0000_0000;
array[29908] <= 16'b0000_0000_0000_0000;
array[29909] <= 16'b0000_0000_0000_0000;
array[29910] <= 16'b0000_0000_0000_0000;
array[29911] <= 16'b0000_0000_0000_0000;
array[29912] <= 16'b0000_0000_0000_0000;
array[29913] <= 16'b0000_0000_0000_0000;
array[29914] <= 16'b0000_0000_0000_0000;
array[29915] <= 16'b0000_0000_0000_0000;
array[29916] <= 16'b0000_0000_0000_0000;
array[29917] <= 16'b0000_0000_0000_0000;
array[29918] <= 16'b0000_0000_0000_0000;
array[29919] <= 16'b0000_0000_0000_0000;
array[29920] <= 16'b0000_0000_0000_0000;
array[29921] <= 16'b0000_0000_0000_0000;
array[29922] <= 16'b0000_0000_0000_0000;
array[29923] <= 16'b0000_0000_0000_0000;
array[29924] <= 16'b0000_0000_0000_0000;
array[29925] <= 16'b0000_0000_0000_0000;
array[29926] <= 16'b0000_0000_0000_0000;
array[29927] <= 16'b0000_0000_0000_0000;
array[29928] <= 16'b0000_0000_0000_0000;
array[29929] <= 16'b0000_0000_0000_0000;
array[29930] <= 16'b0000_0000_0000_0000;
array[29931] <= 16'b0000_0000_0000_0000;
array[29932] <= 16'b0000_0000_0000_0000;
array[29933] <= 16'b0000_0000_0000_0000;
array[29934] <= 16'b0000_0000_0000_0000;
array[29935] <= 16'b0000_0000_0000_0000;
array[29936] <= 16'b0000_0000_0000_0000;
array[29937] <= 16'b0000_0000_0000_0000;
array[29938] <= 16'b0000_0000_0000_0000;
array[29939] <= 16'b0000_0000_0000_0000;
array[29940] <= 16'b0000_0000_0000_0000;
array[29941] <= 16'b0000_0000_0000_0000;
array[29942] <= 16'b0000_0000_0000_0000;
array[29943] <= 16'b0000_0000_0000_0000;
array[29944] <= 16'b0000_0000_0000_0000;
array[29945] <= 16'b0000_0000_0000_0000;
array[29946] <= 16'b0000_0000_0000_0000;
array[29947] <= 16'b0000_0000_0000_0000;
array[29948] <= 16'b0000_0000_0000_0000;
array[29949] <= 16'b0000_0000_0000_0000;
array[29950] <= 16'b0000_0000_0000_0000;
array[29951] <= 16'b0000_0000_0000_0000;
array[29952] <= 16'b0000_0000_0000_0000;
array[29953] <= 16'b0000_0000_0000_0000;
array[29954] <= 16'b0000_0000_0000_0000;
array[29955] <= 16'b0000_0000_0000_0000;
array[29956] <= 16'b0000_0000_0000_0000;
array[29957] <= 16'b0000_0000_0000_0000;
array[29958] <= 16'b0000_0000_0000_0000;
array[29959] <= 16'b0000_0000_0000_0000;
array[29960] <= 16'b0000_0000_0000_0000;
array[29961] <= 16'b0000_0000_0000_0000;
array[29962] <= 16'b0000_0000_0000_0000;
array[29963] <= 16'b0000_0000_0000_0000;
array[29964] <= 16'b0000_0000_0000_0000;
array[29965] <= 16'b0000_0000_0000_0000;
array[29966] <= 16'b0000_0000_0000_0000;
array[29967] <= 16'b0000_0000_0000_0000;
array[29968] <= 16'b0000_0000_0000_0000;
array[29969] <= 16'b0000_0000_0000_0000;
array[29970] <= 16'b0000_0000_0000_0000;
array[29971] <= 16'b0000_0000_0000_0000;
array[29972] <= 16'b0000_0000_0000_0000;
array[29973] <= 16'b0000_0000_0000_0000;
array[29974] <= 16'b0000_0000_0000_0000;
array[29975] <= 16'b0000_0000_0000_0000;
array[29976] <= 16'b0000_0000_0000_0000;
array[29977] <= 16'b0000_0000_0000_0000;
array[29978] <= 16'b0000_0000_0000_0000;
array[29979] <= 16'b0000_0000_0000_0000;
array[29980] <= 16'b0000_0000_0000_0000;
array[29981] <= 16'b0000_0000_0000_0000;
array[29982] <= 16'b0000_0000_0000_0000;
array[29983] <= 16'b0000_0000_0000_0000;
array[29984] <= 16'b0000_0000_0000_0000;
array[29985] <= 16'b0000_0000_0000_0000;
array[29986] <= 16'b0000_0000_0000_0000;
array[29987] <= 16'b0000_0000_0000_0000;
array[29988] <= 16'b0000_0000_0000_0000;
array[29989] <= 16'b0000_0000_0000_0000;
array[29990] <= 16'b0000_0000_0000_0000;
array[29991] <= 16'b0000_0000_0000_0000;
array[29992] <= 16'b0000_0000_0000_0000;
array[29993] <= 16'b0000_0000_0000_0000;
array[29994] <= 16'b0000_0000_0000_0000;
array[29995] <= 16'b0000_0000_0000_0000;
array[29996] <= 16'b0000_0000_0000_0000;
array[29997] <= 16'b0000_0000_0000_0000;
array[29998] <= 16'b0000_0000_0000_0000;
array[29999] <= 16'b0000_0000_0000_0000;
array[30000] <= 16'b0000_0000_0000_0000;
array[30001] <= 16'b0000_0000_0000_0000;
array[30002] <= 16'b0000_0000_0000_0000;
array[30003] <= 16'b0000_0000_0000_0000;
array[30004] <= 16'b0000_0000_0000_0000;
array[30005] <= 16'b0000_0000_0000_0000;
array[30006] <= 16'b0000_0000_0000_0000;
array[30007] <= 16'b0000_0000_0000_0000;
array[30008] <= 16'b0000_0000_0000_0000;
array[30009] <= 16'b0000_0000_0000_0000;
array[30010] <= 16'b0000_0000_0000_0000;
array[30011] <= 16'b0000_0000_0000_0000;
array[30012] <= 16'b0000_0000_0000_0000;
array[30013] <= 16'b0000_0000_0000_0000;
array[30014] <= 16'b0000_0000_0000_0000;
array[30015] <= 16'b0000_0000_0000_0000;
array[30016] <= 16'b0000_0000_0000_0000;
array[30017] <= 16'b0000_0000_0000_0000;
array[30018] <= 16'b0000_0000_0000_0000;
array[30019] <= 16'b0000_0000_0000_0000;
array[30020] <= 16'b0000_0000_0000_0000;
array[30021] <= 16'b0000_0000_0000_0000;
array[30022] <= 16'b0000_0000_0000_0000;
array[30023] <= 16'b0000_0000_0000_0000;
array[30024] <= 16'b0000_0000_0000_0000;
array[30025] <= 16'b0000_0000_0000_0000;
array[30026] <= 16'b0000_0000_0000_0000;
array[30027] <= 16'b0000_0000_0000_0000;
array[30028] <= 16'b0000_0000_0000_0000;
array[30029] <= 16'b0000_0000_0000_0000;
array[30030] <= 16'b0000_0000_0000_0000;
array[30031] <= 16'b0000_0000_0000_0000;
array[30032] <= 16'b0000_0000_0000_0000;
array[30033] <= 16'b0000_0000_0000_0000;
array[30034] <= 16'b0000_0000_0000_0000;
array[30035] <= 16'b0000_0000_0000_0000;
array[30036] <= 16'b0000_0000_0000_0000;
array[30037] <= 16'b0000_0000_0000_0000;
array[30038] <= 16'b0000_0000_0000_0000;
array[30039] <= 16'b0000_0000_0000_0000;
array[30040] <= 16'b0000_0000_0000_0000;
array[30041] <= 16'b0000_0000_0000_0000;
array[30042] <= 16'b0000_0000_0000_0000;
array[30043] <= 16'b0000_0000_0000_0000;
array[30044] <= 16'b0000_0000_0000_0000;
array[30045] <= 16'b0000_0000_0000_0000;
array[30046] <= 16'b0000_0000_0000_0000;
array[30047] <= 16'b0000_0000_0000_0000;
array[30048] <= 16'b0000_0000_0000_0000;
array[30049] <= 16'b0000_0000_0000_0000;
array[30050] <= 16'b0000_0000_0000_0000;
array[30051] <= 16'b0000_0000_0000_0000;
array[30052] <= 16'b0000_0000_0000_0000;
array[30053] <= 16'b0000_0000_0000_0000;
array[30054] <= 16'b0000_0000_0000_0000;
array[30055] <= 16'b0000_0000_0000_0000;
array[30056] <= 16'b0000_0000_0000_0000;
array[30057] <= 16'b0000_0000_0000_0000;
array[30058] <= 16'b0000_0000_0000_0000;
array[30059] <= 16'b0000_0000_0000_0000;
array[30060] <= 16'b0000_0000_0000_0000;
array[30061] <= 16'b0000_0000_0000_0000;
array[30062] <= 16'b0000_0000_0000_0000;
array[30063] <= 16'b0000_0000_0000_0000;
array[30064] <= 16'b0000_0000_0000_0000;
array[30065] <= 16'b0000_0000_0000_0000;
array[30066] <= 16'b0000_0000_0000_0000;
array[30067] <= 16'b0000_0000_0000_0000;
array[30068] <= 16'b0000_0000_0000_0000;
array[30069] <= 16'b0000_0000_0000_0000;
array[30070] <= 16'b0000_0000_0000_0000;
array[30071] <= 16'b0000_0000_0000_0000;
array[30072] <= 16'b0000_0000_0000_0000;
array[30073] <= 16'b0000_0000_0000_0000;
array[30074] <= 16'b0000_0000_0000_0000;
array[30075] <= 16'b0000_0000_0000_0000;
array[30076] <= 16'b0000_0000_0000_0000;
array[30077] <= 16'b0000_0000_0000_0000;
array[30078] <= 16'b0000_0000_0000_0000;
array[30079] <= 16'b0000_0000_0000_0000;
array[30080] <= 16'b0000_0000_0000_0000;
array[30081] <= 16'b0000_0000_0000_0000;
array[30082] <= 16'b0000_0000_0000_0000;
array[30083] <= 16'b0000_0000_0000_0000;
array[30084] <= 16'b0000_0000_0000_0000;
array[30085] <= 16'b0000_0000_0000_0000;
array[30086] <= 16'b0000_0000_0000_0000;
array[30087] <= 16'b0000_0000_0000_0000;
array[30088] <= 16'b0000_0000_0000_0000;
array[30089] <= 16'b0000_0000_0000_0000;
array[30090] <= 16'b0000_0000_0000_0000;
array[30091] <= 16'b0000_0000_0000_0000;
array[30092] <= 16'b0000_0000_0000_0000;
array[30093] <= 16'b0000_0000_0000_0000;
array[30094] <= 16'b0000_0000_0000_0000;
array[30095] <= 16'b0000_0000_0000_0000;
array[30096] <= 16'b0000_0000_0000_0000;
array[30097] <= 16'b0000_0000_0000_0000;
array[30098] <= 16'b0000_0000_0000_0000;
array[30099] <= 16'b0000_0000_0000_0000;
array[30100] <= 16'b0000_0000_0000_0000;
array[30101] <= 16'b0000_0000_0000_0000;
array[30102] <= 16'b0000_0000_0000_0000;
array[30103] <= 16'b0000_0000_0000_0000;
array[30104] <= 16'b0000_0000_0000_0000;
array[30105] <= 16'b0000_0000_0000_0000;
array[30106] <= 16'b0000_0000_0000_0000;
array[30107] <= 16'b0000_0000_0000_0000;
array[30108] <= 16'b0000_0000_0000_0000;
array[30109] <= 16'b0000_0000_0000_0000;
array[30110] <= 16'b0000_0000_0000_0000;
array[30111] <= 16'b0000_0000_0000_0000;
array[30112] <= 16'b0000_0000_0000_0000;
array[30113] <= 16'b0000_0000_0000_0000;
array[30114] <= 16'b0000_0000_0000_0000;
array[30115] <= 16'b0000_0000_0000_0000;
array[30116] <= 16'b0000_0000_0000_0000;
array[30117] <= 16'b0000_0000_0000_0000;
array[30118] <= 16'b0000_0000_0000_0000;
array[30119] <= 16'b0000_0000_0000_0000;
array[30120] <= 16'b0000_0000_0000_0000;
array[30121] <= 16'b0000_0000_0000_0000;
array[30122] <= 16'b0000_0000_0000_0000;
array[30123] <= 16'b0000_0000_0000_0000;
array[30124] <= 16'b0000_0000_0000_0000;
array[30125] <= 16'b0000_0000_0000_0000;
array[30126] <= 16'b0000_0000_0000_0000;
array[30127] <= 16'b0000_0000_0000_0000;
array[30128] <= 16'b0000_0000_0000_0000;
array[30129] <= 16'b0000_0000_0000_0000;
array[30130] <= 16'b0000_0000_0000_0000;
array[30131] <= 16'b0000_0000_0000_0000;
array[30132] <= 16'b0000_0000_0000_0000;
array[30133] <= 16'b0000_0000_0000_0000;
array[30134] <= 16'b0000_0000_0000_0000;
array[30135] <= 16'b0000_0000_0000_0000;
array[30136] <= 16'b0000_0000_0000_0000;
array[30137] <= 16'b0000_0000_0000_0000;
array[30138] <= 16'b0000_0000_0000_0000;
array[30139] <= 16'b0000_0000_0000_0000;
array[30140] <= 16'b0000_0000_0000_0000;
array[30141] <= 16'b0000_0000_0000_0000;
array[30142] <= 16'b0000_0000_0000_0000;
array[30143] <= 16'b0000_0000_0000_0000;
array[30144] <= 16'b0000_0000_0000_0000;
array[30145] <= 16'b0000_0000_0000_0000;
array[30146] <= 16'b0000_0000_0000_0000;
array[30147] <= 16'b0000_0000_0000_0000;
array[30148] <= 16'b0000_0000_0000_0000;
array[30149] <= 16'b0000_0000_0000_0000;
array[30150] <= 16'b0000_0000_0000_0000;
array[30151] <= 16'b0000_0000_0000_0000;
array[30152] <= 16'b0000_0000_0000_0000;
array[30153] <= 16'b0000_0000_0000_0000;
array[30154] <= 16'b0000_0000_0000_0000;
array[30155] <= 16'b0000_0000_0000_0000;
array[30156] <= 16'b0000_0000_0000_0000;
array[30157] <= 16'b0000_0000_0000_0000;
array[30158] <= 16'b0000_0000_0000_0000;
array[30159] <= 16'b0000_0000_0000_0000;
array[30160] <= 16'b0000_0000_0000_0000;
array[30161] <= 16'b0000_0000_0000_0000;
array[30162] <= 16'b0000_0000_0000_0000;
array[30163] <= 16'b0000_0000_0000_0000;
array[30164] <= 16'b0000_0000_0000_0000;
array[30165] <= 16'b0000_0000_0000_0000;
array[30166] <= 16'b0000_0000_0000_0000;
array[30167] <= 16'b0000_0000_0000_0000;
array[30168] <= 16'b0000_0000_0000_0000;
array[30169] <= 16'b0000_0000_0000_0000;
array[30170] <= 16'b0000_0000_0000_0000;
array[30171] <= 16'b0000_0000_0000_0000;
array[30172] <= 16'b0000_0000_0000_0000;
array[30173] <= 16'b0000_0000_0000_0000;
array[30174] <= 16'b0000_0000_0000_0000;
array[30175] <= 16'b0000_0000_0000_0000;
array[30176] <= 16'b0000_0000_0000_0000;
array[30177] <= 16'b0000_0000_0000_0000;
array[30178] <= 16'b0000_0000_0000_0000;
array[30179] <= 16'b0000_0000_0000_0000;
array[30180] <= 16'b0000_0000_0000_0000;
array[30181] <= 16'b0000_0000_0000_0000;
array[30182] <= 16'b0000_0000_0000_0000;
array[30183] <= 16'b0000_0000_0000_0000;
array[30184] <= 16'b0000_0000_0000_0000;
array[30185] <= 16'b0000_0000_0000_0000;
array[30186] <= 16'b0000_0000_0000_0000;
array[30187] <= 16'b0000_0000_0000_0000;
array[30188] <= 16'b0000_0000_0000_0000;
array[30189] <= 16'b0000_0000_0000_0000;
array[30190] <= 16'b0000_0000_0000_0000;
array[30191] <= 16'b0000_0000_0000_0000;
array[30192] <= 16'b0000_0000_0000_0000;
array[30193] <= 16'b0000_0000_0000_0000;
array[30194] <= 16'b0000_0000_0000_0000;
array[30195] <= 16'b0000_0000_0000_0000;
array[30196] <= 16'b0000_0000_0000_0000;
array[30197] <= 16'b0000_0000_0000_0000;
array[30198] <= 16'b0000_0000_0000_0000;
array[30199] <= 16'b0000_0000_0000_0000;
array[30200] <= 16'b0000_0000_0000_0000;
array[30201] <= 16'b0000_0000_0000_0000;
array[30202] <= 16'b0000_0000_0000_0000;
array[30203] <= 16'b0000_0000_0000_0000;
array[30204] <= 16'b0000_0000_0000_0000;
array[30205] <= 16'b0000_0000_0000_0000;
array[30206] <= 16'b0000_0000_0000_0000;
array[30207] <= 16'b0000_0000_0000_0000;
array[30208] <= 16'b0000_0000_0000_0000;
array[30209] <= 16'b0000_0000_0000_0000;
array[30210] <= 16'b0000_0000_0000_0000;
array[30211] <= 16'b0000_0000_0000_0000;
array[30212] <= 16'b0000_0000_0000_0000;
array[30213] <= 16'b0000_0000_0000_0000;
array[30214] <= 16'b0000_0000_0000_0000;
array[30215] <= 16'b0000_0000_0000_0000;
array[30216] <= 16'b0000_0000_0000_0000;
array[30217] <= 16'b0000_0000_0000_0000;
array[30218] <= 16'b0000_0000_0000_0000;
array[30219] <= 16'b0000_0000_0000_0000;
array[30220] <= 16'b0000_0000_0000_0000;
array[30221] <= 16'b0000_0000_0000_0000;
array[30222] <= 16'b0000_0000_0000_0000;
array[30223] <= 16'b0000_0000_0000_0000;
array[30224] <= 16'b0000_0000_0000_0000;
array[30225] <= 16'b0000_0000_0000_0000;
array[30226] <= 16'b0000_0000_0000_0000;
array[30227] <= 16'b0000_0000_0000_0000;
array[30228] <= 16'b0000_0000_0000_0000;
array[30229] <= 16'b0000_0000_0000_0000;
array[30230] <= 16'b0000_0000_0000_0000;
array[30231] <= 16'b0000_0000_0000_0000;
array[30232] <= 16'b0000_0000_0000_0000;
array[30233] <= 16'b0000_0000_0000_0000;
array[30234] <= 16'b0000_0000_0000_0000;
array[30235] <= 16'b0000_0000_0000_0000;
array[30236] <= 16'b0000_0000_0000_0000;
array[30237] <= 16'b0000_0000_0000_0000;
array[30238] <= 16'b0000_0000_0000_0000;
array[30239] <= 16'b0000_0000_0000_0000;
array[30240] <= 16'b0000_0000_0000_0000;
array[30241] <= 16'b0000_0000_0000_0000;
array[30242] <= 16'b0000_0000_0000_0000;
array[30243] <= 16'b0000_0000_0000_0000;
array[30244] <= 16'b0000_0000_0000_0000;
array[30245] <= 16'b0000_0000_0000_0000;
array[30246] <= 16'b0000_0000_0000_0000;
array[30247] <= 16'b0000_0000_0000_0000;
array[30248] <= 16'b0000_0000_0000_0000;
array[30249] <= 16'b0000_0000_0000_0000;
array[30250] <= 16'b0000_0000_0000_0000;
array[30251] <= 16'b0000_0000_0000_0000;
array[30252] <= 16'b0000_0000_0000_0000;
array[30253] <= 16'b0000_0000_0000_0000;
array[30254] <= 16'b0000_0000_0000_0000;
array[30255] <= 16'b0000_0000_0000_0000;
array[30256] <= 16'b0000_0000_0000_0000;
array[30257] <= 16'b0000_0000_0000_0000;
array[30258] <= 16'b0000_0000_0000_0000;
array[30259] <= 16'b0000_0000_0000_0000;
array[30260] <= 16'b0000_0000_0000_0000;
array[30261] <= 16'b0000_0000_0000_0000;
array[30262] <= 16'b0000_0000_0000_0000;
array[30263] <= 16'b0000_0000_0000_0000;
array[30264] <= 16'b0000_0000_0000_0000;
array[30265] <= 16'b0000_0000_0000_0000;
array[30266] <= 16'b0000_0000_0000_0000;
array[30267] <= 16'b0000_0000_0000_0000;
array[30268] <= 16'b0000_0000_0000_0000;
array[30269] <= 16'b0000_0000_0000_0000;
array[30270] <= 16'b0000_0000_0000_0000;
array[30271] <= 16'b0000_0000_0000_0000;
array[30272] <= 16'b0000_0000_0000_0000;
array[30273] <= 16'b0000_0000_0000_0000;
array[30274] <= 16'b0000_0000_0000_0000;
array[30275] <= 16'b0000_0000_0000_0000;
array[30276] <= 16'b0000_0000_0000_0000;
array[30277] <= 16'b0000_0000_0000_0000;
array[30278] <= 16'b0000_0000_0000_0000;
array[30279] <= 16'b0000_0000_0000_0000;
array[30280] <= 16'b0000_0000_0000_0000;
array[30281] <= 16'b0000_0000_0000_0000;
array[30282] <= 16'b0000_0000_0000_0000;
array[30283] <= 16'b0000_0000_0000_0000;
array[30284] <= 16'b0000_0000_0000_0000;
array[30285] <= 16'b0000_0000_0000_0000;
array[30286] <= 16'b0000_0000_0000_0000;
array[30287] <= 16'b0000_0000_0000_0000;
array[30288] <= 16'b0000_0000_0000_0000;
array[30289] <= 16'b0000_0000_0000_0000;
array[30290] <= 16'b0000_0000_0000_0000;
array[30291] <= 16'b0000_0000_0000_0000;
array[30292] <= 16'b0000_0000_0000_0000;
array[30293] <= 16'b0000_0000_0000_0000;
array[30294] <= 16'b0000_0000_0000_0000;
array[30295] <= 16'b0000_0000_0000_0000;
array[30296] <= 16'b0000_0000_0000_0000;
array[30297] <= 16'b0000_0000_0000_0000;
array[30298] <= 16'b0000_0000_0000_0000;
array[30299] <= 16'b0000_0000_0000_0000;
array[30300] <= 16'b0000_0000_0000_0000;
array[30301] <= 16'b0000_0000_0000_0000;
array[30302] <= 16'b0000_0000_0000_0000;
array[30303] <= 16'b0000_0000_0000_0000;
array[30304] <= 16'b0000_0000_0000_0000;
array[30305] <= 16'b0000_0000_0000_0000;
array[30306] <= 16'b0000_0000_0000_0000;
array[30307] <= 16'b0000_0000_0000_0000;
array[30308] <= 16'b0000_0000_0000_0000;
array[30309] <= 16'b0000_0000_0000_0000;
array[30310] <= 16'b0000_0000_0000_0000;
array[30311] <= 16'b0000_0000_0000_0000;
array[30312] <= 16'b0000_0000_0000_0000;
array[30313] <= 16'b0000_0000_0000_0000;
array[30314] <= 16'b0000_0000_0000_0000;
array[30315] <= 16'b0000_0000_0000_0000;
array[30316] <= 16'b0000_0000_0000_0000;
array[30317] <= 16'b0000_0000_0000_0000;
array[30318] <= 16'b0000_0000_0000_0000;
array[30319] <= 16'b0000_0000_0000_0000;
array[30320] <= 16'b0000_0000_0000_0000;
array[30321] <= 16'b0000_0000_0000_0000;
array[30322] <= 16'b0000_0000_0000_0000;
array[30323] <= 16'b0000_0000_0000_0000;
array[30324] <= 16'b0000_0000_0000_0000;
array[30325] <= 16'b0000_0000_0000_0000;
array[30326] <= 16'b0000_0000_0000_0000;
array[30327] <= 16'b0000_0000_0000_0000;
array[30328] <= 16'b0000_0000_0000_0000;
array[30329] <= 16'b0000_0000_0000_0000;
array[30330] <= 16'b0000_0000_0000_0000;
array[30331] <= 16'b0000_0000_0000_0000;
array[30332] <= 16'b0000_0000_0000_0000;
array[30333] <= 16'b0000_0000_0000_0000;
array[30334] <= 16'b0000_0000_0000_0000;
array[30335] <= 16'b0000_0000_0000_0000;
array[30336] <= 16'b0000_0000_0000_0000;
array[30337] <= 16'b0000_0000_0000_0000;
array[30338] <= 16'b0000_0000_0000_0000;
array[30339] <= 16'b0000_0000_0000_0000;
array[30340] <= 16'b0000_0000_0000_0000;
array[30341] <= 16'b0000_0000_0000_0000;
array[30342] <= 16'b0000_0000_0000_0000;
array[30343] <= 16'b0000_0000_0000_0000;
array[30344] <= 16'b0000_0000_0000_0000;
array[30345] <= 16'b0000_0000_0000_0000;
array[30346] <= 16'b0000_0000_0000_0000;
array[30347] <= 16'b0000_0000_0000_0000;
array[30348] <= 16'b0000_0000_0000_0000;
array[30349] <= 16'b0000_0000_0000_0000;
array[30350] <= 16'b0000_0000_0000_0000;
array[30351] <= 16'b0000_0000_0000_0000;
array[30352] <= 16'b0000_0000_0000_0000;
array[30353] <= 16'b0000_0000_0000_0000;
array[30354] <= 16'b0000_0000_0000_0000;
array[30355] <= 16'b0000_0000_0000_0000;
array[30356] <= 16'b0000_0000_0000_0000;
array[30357] <= 16'b0000_0000_0000_0000;
array[30358] <= 16'b0000_0000_0000_0000;
array[30359] <= 16'b0000_0000_0000_0000;
array[30360] <= 16'b0000_0000_0000_0000;
array[30361] <= 16'b0000_0000_0000_0000;
array[30362] <= 16'b0000_0000_0000_0000;
array[30363] <= 16'b0000_0000_0000_0000;
array[30364] <= 16'b0000_0000_0000_0000;
array[30365] <= 16'b0000_0000_0000_0000;
array[30366] <= 16'b0000_0000_0000_0000;
array[30367] <= 16'b0000_0000_0000_0000;
array[30368] <= 16'b0000_0000_0000_0000;
array[30369] <= 16'b0000_0000_0000_0000;
array[30370] <= 16'b0000_0000_0000_0000;
array[30371] <= 16'b0000_0000_0000_0000;
array[30372] <= 16'b0000_0000_0000_0000;
array[30373] <= 16'b0000_0000_0000_0000;
array[30374] <= 16'b0000_0000_0000_0000;
array[30375] <= 16'b0000_0000_0000_0000;
array[30376] <= 16'b0000_0000_0000_0000;
array[30377] <= 16'b0000_0000_0000_0000;
array[30378] <= 16'b0000_0000_0000_0000;
array[30379] <= 16'b0000_0000_0000_0000;
array[30380] <= 16'b0000_0000_0000_0000;
array[30381] <= 16'b0000_0000_0000_0000;
array[30382] <= 16'b0000_0000_0000_0000;
array[30383] <= 16'b0000_0000_0000_0000;
array[30384] <= 16'b0000_0000_0000_0000;
array[30385] <= 16'b0000_0000_0000_0000;
array[30386] <= 16'b0000_0000_0000_0000;
array[30387] <= 16'b0000_0000_0000_0000;
array[30388] <= 16'b0000_0000_0000_0000;
array[30389] <= 16'b0000_0000_0000_0000;
array[30390] <= 16'b0000_0000_0000_0000;
array[30391] <= 16'b0000_0000_0000_0000;
array[30392] <= 16'b0000_0000_0000_0000;
array[30393] <= 16'b0000_0000_0000_0000;
array[30394] <= 16'b0000_0000_0000_0000;
array[30395] <= 16'b0000_0000_0000_0000;
array[30396] <= 16'b0000_0000_0000_0000;
array[30397] <= 16'b0000_0000_0000_0000;
array[30398] <= 16'b0000_0000_0000_0000;
array[30399] <= 16'b0000_0000_0000_0000;
array[30400] <= 16'b0000_0000_0000_0000;
array[30401] <= 16'b0000_0000_0000_0000;
array[30402] <= 16'b0000_0000_0000_0000;
array[30403] <= 16'b0000_0000_0000_0000;
array[30404] <= 16'b0000_0000_0000_0000;
array[30405] <= 16'b0000_0000_0000_0000;
array[30406] <= 16'b0000_0000_0000_0000;
array[30407] <= 16'b0000_0000_0000_0000;
array[30408] <= 16'b0000_0000_0000_0000;
array[30409] <= 16'b0000_0000_0000_0000;
array[30410] <= 16'b0000_0000_0000_0000;
array[30411] <= 16'b0000_0000_0000_0000;
array[30412] <= 16'b0000_0000_0000_0000;
array[30413] <= 16'b0000_0000_0000_0000;
array[30414] <= 16'b0000_0000_0000_0000;
array[30415] <= 16'b0000_0000_0000_0000;
array[30416] <= 16'b0000_0000_0000_0000;
array[30417] <= 16'b0000_0000_0000_0000;
array[30418] <= 16'b0000_0000_0000_0000;
array[30419] <= 16'b0000_0000_0000_0000;
array[30420] <= 16'b0000_0000_0000_0000;
array[30421] <= 16'b0000_0000_0000_0000;
array[30422] <= 16'b0000_0000_0000_0000;
array[30423] <= 16'b0000_0000_0000_0000;
array[30424] <= 16'b0000_0000_0000_0000;
array[30425] <= 16'b0000_0000_0000_0000;
array[30426] <= 16'b0000_0000_0000_0000;
array[30427] <= 16'b0000_0000_0000_0000;
array[30428] <= 16'b0000_0000_0000_0000;
array[30429] <= 16'b0000_0000_0000_0000;
array[30430] <= 16'b0000_0000_0000_0000;
array[30431] <= 16'b0000_0000_0000_0000;
array[30432] <= 16'b0000_0000_0000_0000;
array[30433] <= 16'b0000_0000_0000_0000;
array[30434] <= 16'b0000_0000_0000_0000;
array[30435] <= 16'b0000_0000_0000_0000;
array[30436] <= 16'b0000_0000_0000_0000;
array[30437] <= 16'b0000_0000_0000_0000;
array[30438] <= 16'b0000_0000_0000_0000;
array[30439] <= 16'b0000_0000_0000_0000;
array[30440] <= 16'b0000_0000_0000_0000;
array[30441] <= 16'b0000_0000_0000_0000;
array[30442] <= 16'b0000_0000_0000_0000;
array[30443] <= 16'b0000_0000_0000_0000;
array[30444] <= 16'b0000_0000_0000_0000;
array[30445] <= 16'b0000_0000_0000_0000;
array[30446] <= 16'b0000_0000_0000_0000;
array[30447] <= 16'b0000_0000_0000_0000;
array[30448] <= 16'b0000_0000_0000_0000;
array[30449] <= 16'b0000_0000_0000_0000;
array[30450] <= 16'b0000_0000_0000_0000;
array[30451] <= 16'b0000_0000_0000_0000;
array[30452] <= 16'b0000_0000_0000_0000;
array[30453] <= 16'b0000_0000_0000_0000;
array[30454] <= 16'b0000_0000_0000_0000;
array[30455] <= 16'b0000_0000_0000_0000;
array[30456] <= 16'b0000_0000_0000_0000;
array[30457] <= 16'b0000_0000_0000_0000;
array[30458] <= 16'b0000_0000_0000_0000;
array[30459] <= 16'b0000_0000_0000_0000;
array[30460] <= 16'b0000_0000_0000_0000;
array[30461] <= 16'b0000_0000_0000_0000;
array[30462] <= 16'b0000_0000_0000_0000;
array[30463] <= 16'b0000_0000_0000_0000;
array[30464] <= 16'b0000_0000_0000_0000;
array[30465] <= 16'b0000_0000_0000_0000;
array[30466] <= 16'b0000_0000_0000_0000;
array[30467] <= 16'b0000_0000_0000_0000;
array[30468] <= 16'b0000_0000_0000_0000;
array[30469] <= 16'b0000_0000_0000_0000;
array[30470] <= 16'b0000_0000_0000_0000;
array[30471] <= 16'b0000_0000_0000_0000;
array[30472] <= 16'b0000_0000_0000_0000;
array[30473] <= 16'b0000_0000_0000_0000;
array[30474] <= 16'b0000_0000_0000_0000;
array[30475] <= 16'b0000_0000_0000_0000;
array[30476] <= 16'b0000_0000_0000_0000;
array[30477] <= 16'b0000_0000_0000_0000;
array[30478] <= 16'b0000_0000_0000_0000;
array[30479] <= 16'b0000_0000_0000_0000;
array[30480] <= 16'b0000_0000_0000_0000;
array[30481] <= 16'b0000_0000_0000_0000;
array[30482] <= 16'b0000_0000_0000_0000;
array[30483] <= 16'b0000_0000_0000_0000;
array[30484] <= 16'b0000_0000_0000_0000;
array[30485] <= 16'b0000_0000_0000_0000;
array[30486] <= 16'b0000_0000_0000_0000;
array[30487] <= 16'b0000_0000_0000_0000;
array[30488] <= 16'b0000_0000_0000_0000;
array[30489] <= 16'b0000_0000_0000_0000;
array[30490] <= 16'b0000_0000_0000_0000;
array[30491] <= 16'b0000_0000_0000_0000;
array[30492] <= 16'b0000_0000_0000_0000;
array[30493] <= 16'b0000_0000_0000_0000;
array[30494] <= 16'b0000_0000_0000_0000;
array[30495] <= 16'b0000_0000_0000_0000;
array[30496] <= 16'b0000_0000_0000_0000;
array[30497] <= 16'b0000_0000_0000_0000;
array[30498] <= 16'b0000_0000_0000_0000;
array[30499] <= 16'b0000_0000_0000_0000;
array[30500] <= 16'b0000_0000_0000_0000;
array[30501] <= 16'b0000_0000_0000_0000;
array[30502] <= 16'b0000_0000_0000_0000;
array[30503] <= 16'b0000_0000_0000_0000;
array[30504] <= 16'b0000_0000_0000_0000;
array[30505] <= 16'b0000_0000_0000_0000;
array[30506] <= 16'b0000_0000_0000_0000;
array[30507] <= 16'b0000_0000_0000_0000;
array[30508] <= 16'b0000_0000_0000_0000;
array[30509] <= 16'b0000_0000_0000_0000;
array[30510] <= 16'b0000_0000_0000_0000;
array[30511] <= 16'b0000_0000_0000_0000;
array[30512] <= 16'b0000_0000_0000_0000;
array[30513] <= 16'b0000_0000_0000_0000;
array[30514] <= 16'b0000_0000_0000_0000;
array[30515] <= 16'b0000_0000_0000_0000;
array[30516] <= 16'b0000_0000_0000_0000;
array[30517] <= 16'b0000_0000_0000_0000;
array[30518] <= 16'b0000_0000_0000_0000;
array[30519] <= 16'b0000_0000_0000_0000;
array[30520] <= 16'b0000_0000_0000_0000;
array[30521] <= 16'b0000_0000_0000_0000;
array[30522] <= 16'b0000_0000_0000_0000;
array[30523] <= 16'b0000_0000_0000_0000;
array[30524] <= 16'b0000_0000_0000_0000;
array[30525] <= 16'b0000_0000_0000_0000;
array[30526] <= 16'b0000_0000_0000_0000;
array[30527] <= 16'b0000_0000_0000_0000;
array[30528] <= 16'b0000_0000_0000_0000;
array[30529] <= 16'b0000_0000_0000_0000;
array[30530] <= 16'b0000_0000_0000_0000;
array[30531] <= 16'b0000_0000_0000_0000;
array[30532] <= 16'b0000_0000_0000_0000;
array[30533] <= 16'b0000_0000_0000_0000;
array[30534] <= 16'b0000_0000_0000_0000;
array[30535] <= 16'b0000_0000_0000_0000;
array[30536] <= 16'b0000_0000_0000_0000;
array[30537] <= 16'b0000_0000_0000_0000;
array[30538] <= 16'b0000_0000_0000_0000;
array[30539] <= 16'b0000_0000_0000_0000;
array[30540] <= 16'b0000_0000_0000_0000;
array[30541] <= 16'b0000_0000_0000_0000;
array[30542] <= 16'b0000_0000_0000_0000;
array[30543] <= 16'b0000_0000_0000_0000;
array[30544] <= 16'b0000_0000_0000_0000;
array[30545] <= 16'b0000_0000_0000_0000;
array[30546] <= 16'b0000_0000_0000_0000;
array[30547] <= 16'b0000_0000_0000_0000;
array[30548] <= 16'b0000_0000_0000_0000;
array[30549] <= 16'b0000_0000_0000_0000;
array[30550] <= 16'b0000_0000_0000_0000;
array[30551] <= 16'b0000_0000_0000_0000;
array[30552] <= 16'b0000_0000_0000_0000;
array[30553] <= 16'b0000_0000_0000_0000;
array[30554] <= 16'b0000_0000_0000_0000;
array[30555] <= 16'b0000_0000_0000_0000;
array[30556] <= 16'b0000_0000_0000_0000;
array[30557] <= 16'b0000_0000_0000_0000;
array[30558] <= 16'b0000_0000_0000_0000;
array[30559] <= 16'b0000_0000_0000_0000;
array[30560] <= 16'b0000_0000_0000_0000;
array[30561] <= 16'b0000_0000_0000_0000;
array[30562] <= 16'b0000_0000_0000_0000;
array[30563] <= 16'b0000_0000_0000_0000;
array[30564] <= 16'b0000_0000_0000_0000;
array[30565] <= 16'b0000_0000_0000_0000;
array[30566] <= 16'b0000_0000_0000_0000;
array[30567] <= 16'b0000_0000_0000_0000;
array[30568] <= 16'b0000_0000_0000_0000;
array[30569] <= 16'b0000_0000_0000_0000;
array[30570] <= 16'b0000_0000_0000_0000;
array[30571] <= 16'b0000_0000_0000_0000;
array[30572] <= 16'b0000_0000_0000_0000;
array[30573] <= 16'b0000_0000_0000_0000;
array[30574] <= 16'b0000_0000_0000_0000;
array[30575] <= 16'b0000_0000_0000_0000;
array[30576] <= 16'b0000_0000_0000_0000;
array[30577] <= 16'b0000_0000_0000_0000;
array[30578] <= 16'b0000_0000_0000_0000;
array[30579] <= 16'b0000_0000_0000_0000;
array[30580] <= 16'b0000_0000_0000_0000;
array[30581] <= 16'b0000_0000_0000_0000;
array[30582] <= 16'b0000_0000_0000_0000;
array[30583] <= 16'b0000_0000_0000_0000;
array[30584] <= 16'b0000_0000_0000_0000;
array[30585] <= 16'b0000_0000_0000_0000;
array[30586] <= 16'b0000_0000_0000_0000;
array[30587] <= 16'b0000_0000_0000_0000;
array[30588] <= 16'b0000_0000_0000_0000;
array[30589] <= 16'b0000_0000_0000_0000;
array[30590] <= 16'b0000_0000_0000_0000;
array[30591] <= 16'b0000_0000_0000_0000;
array[30592] <= 16'b0000_0000_0000_0000;
array[30593] <= 16'b0000_0000_0000_0000;
array[30594] <= 16'b0000_0000_0000_0000;
array[30595] <= 16'b0000_0000_0000_0000;
array[30596] <= 16'b0000_0000_0000_0000;
array[30597] <= 16'b0000_0000_0000_0000;
array[30598] <= 16'b0000_0000_0000_0000;
array[30599] <= 16'b0000_0000_0000_0000;
array[30600] <= 16'b0000_0000_0000_0000;
array[30601] <= 16'b0000_0000_0000_0000;
array[30602] <= 16'b0000_0000_0000_0000;
array[30603] <= 16'b0000_0000_0000_0000;
array[30604] <= 16'b0000_0000_0000_0000;
array[30605] <= 16'b0000_0000_0000_0000;
array[30606] <= 16'b0000_0000_0000_0000;
array[30607] <= 16'b0000_0000_0000_0000;
array[30608] <= 16'b0000_0000_0000_0000;
array[30609] <= 16'b0000_0000_0000_0000;
array[30610] <= 16'b0000_0000_0000_0000;
array[30611] <= 16'b0000_0000_0000_0000;
array[30612] <= 16'b0000_0000_0000_0000;
array[30613] <= 16'b0000_0000_0000_0000;
array[30614] <= 16'b0000_0000_0000_0000;
array[30615] <= 16'b0000_0000_0000_0000;
array[30616] <= 16'b0000_0000_0000_0000;
array[30617] <= 16'b0000_0000_0000_0000;
array[30618] <= 16'b0000_0000_0000_0000;
array[30619] <= 16'b0000_0000_0000_0000;
array[30620] <= 16'b0000_0000_0000_0000;
array[30621] <= 16'b0000_0000_0000_0000;
array[30622] <= 16'b0000_0000_0000_0000;
array[30623] <= 16'b0000_0000_0000_0000;
array[30624] <= 16'b0000_0000_0000_0000;
array[30625] <= 16'b0000_0000_0000_0000;
array[30626] <= 16'b0000_0000_0000_0000;
array[30627] <= 16'b0000_0000_0000_0000;
array[30628] <= 16'b0000_0000_0000_0000;
array[30629] <= 16'b0000_0000_0000_0000;
array[30630] <= 16'b0000_0000_0000_0000;
array[30631] <= 16'b0000_0000_0000_0000;
array[30632] <= 16'b0000_0000_0000_0000;
array[30633] <= 16'b0000_0000_0000_0000;
array[30634] <= 16'b0000_0000_0000_0000;
array[30635] <= 16'b0000_0000_0000_0000;
array[30636] <= 16'b0000_0000_0000_0000;
array[30637] <= 16'b0000_0000_0000_0000;
array[30638] <= 16'b0000_0000_0000_0000;
array[30639] <= 16'b0000_0000_0000_0000;
array[30640] <= 16'b0000_0000_0000_0000;
array[30641] <= 16'b0000_0000_0000_0000;
array[30642] <= 16'b0000_0000_0000_0000;
array[30643] <= 16'b0000_0000_0000_0000;
array[30644] <= 16'b0000_0000_0000_0000;
array[30645] <= 16'b0000_0000_0000_0000;
array[30646] <= 16'b0000_0000_0000_0000;
array[30647] <= 16'b0000_0000_0000_0000;
array[30648] <= 16'b0000_0000_0000_0000;
array[30649] <= 16'b0000_0000_0000_0000;
array[30650] <= 16'b0000_0000_0000_0000;
array[30651] <= 16'b0000_0000_0000_0000;
array[30652] <= 16'b0000_0000_0000_0000;
array[30653] <= 16'b0000_0000_0000_0000;
array[30654] <= 16'b0000_0000_0000_0000;
array[30655] <= 16'b0000_0000_0000_0000;
array[30656] <= 16'b0000_0000_0000_0000;
array[30657] <= 16'b0000_0000_0000_0000;
array[30658] <= 16'b0000_0000_0000_0000;
array[30659] <= 16'b0000_0000_0000_0000;
array[30660] <= 16'b0000_0000_0000_0000;
array[30661] <= 16'b0000_0000_0000_0000;
array[30662] <= 16'b0000_0000_0000_0000;
array[30663] <= 16'b0000_0000_0000_0000;
array[30664] <= 16'b0000_0000_0000_0000;
array[30665] <= 16'b0000_0000_0000_0000;
array[30666] <= 16'b0000_0000_0000_0000;
array[30667] <= 16'b0000_0000_0000_0000;
array[30668] <= 16'b0000_0000_0000_0000;
array[30669] <= 16'b0000_0000_0000_0000;
array[30670] <= 16'b0000_0000_0000_0000;
array[30671] <= 16'b0000_0000_0000_0000;
array[30672] <= 16'b0000_0000_0000_0000;
array[30673] <= 16'b0000_0000_0000_0000;
array[30674] <= 16'b0000_0000_0000_0000;
array[30675] <= 16'b0000_0000_0000_0000;
array[30676] <= 16'b0000_0000_0000_0000;
array[30677] <= 16'b0000_0000_0000_0000;
array[30678] <= 16'b0000_0000_0000_0000;
array[30679] <= 16'b0000_0000_0000_0000;
array[30680] <= 16'b0000_0000_0000_0000;
array[30681] <= 16'b0000_0000_0000_0000;
array[30682] <= 16'b0000_0000_0000_0000;
array[30683] <= 16'b0000_0000_0000_0000;
array[30684] <= 16'b0000_0000_0000_0000;
array[30685] <= 16'b0000_0000_0000_0000;
array[30686] <= 16'b0000_0000_0000_0000;
array[30687] <= 16'b0000_0000_0000_0000;
array[30688] <= 16'b0000_0000_0000_0000;
array[30689] <= 16'b0000_0000_0000_0000;
array[30690] <= 16'b0000_0000_0000_0000;
array[30691] <= 16'b0000_0000_0000_0000;
array[30692] <= 16'b0000_0000_0000_0000;
array[30693] <= 16'b0000_0000_0000_0000;
array[30694] <= 16'b0000_0000_0000_0000;
array[30695] <= 16'b0000_0000_0000_0000;
array[30696] <= 16'b0000_0000_0000_0000;
array[30697] <= 16'b0000_0000_0000_0000;
array[30698] <= 16'b0000_0000_0000_0000;
array[30699] <= 16'b0000_0000_0000_0000;
array[30700] <= 16'b0000_0000_0000_0000;
array[30701] <= 16'b0000_0000_0000_0000;
array[30702] <= 16'b0000_0000_0000_0000;
array[30703] <= 16'b0000_0000_0000_0000;
array[30704] <= 16'b0000_0000_0000_0000;
array[30705] <= 16'b0000_0000_0000_0000;
array[30706] <= 16'b0000_0000_0000_0000;
array[30707] <= 16'b0000_0000_0000_0000;
array[30708] <= 16'b0000_0000_0000_0000;
array[30709] <= 16'b0000_0000_0000_0000;
array[30710] <= 16'b0000_0000_0000_0000;
array[30711] <= 16'b0000_0000_0000_0000;
array[30712] <= 16'b0000_0000_0000_0000;
array[30713] <= 16'b0000_0000_0000_0000;
array[30714] <= 16'b0000_0000_0000_0000;
array[30715] <= 16'b0000_0000_0000_0000;
array[30716] <= 16'b0000_0000_0000_0000;
array[30717] <= 16'b0000_0000_0000_0000;
array[30718] <= 16'b0000_0000_0000_0000;
array[30719] <= 16'b0000_0000_0000_0000;
array[30720] <= 16'b0000_0000_0000_0000;
array[30721] <= 16'b0000_0000_0000_0000;
array[30722] <= 16'b0000_0000_0000_0000;
array[30723] <= 16'b0000_0000_0000_0000;
array[30724] <= 16'b0000_0000_0000_0000;
array[30725] <= 16'b0000_0000_0000_0000;
array[30726] <= 16'b0000_0000_0000_0000;
array[30727] <= 16'b0000_0000_0000_0000;
array[30728] <= 16'b0000_0000_0000_0000;
array[30729] <= 16'b0000_0000_0000_0000;
array[30730] <= 16'b0000_0000_0000_0000;
array[30731] <= 16'b0000_0000_0000_0000;
array[30732] <= 16'b0000_0000_0000_0000;
array[30733] <= 16'b0000_0000_0000_0000;
array[30734] <= 16'b0000_0000_0000_0000;
array[30735] <= 16'b0000_0000_0000_0000;
array[30736] <= 16'b0000_0000_0000_0000;
array[30737] <= 16'b0000_0000_0000_0000;
array[30738] <= 16'b0000_0000_0000_0000;
array[30739] <= 16'b0000_0000_0000_0000;
array[30740] <= 16'b0000_0000_0000_0000;
array[30741] <= 16'b0000_0000_0000_0000;
array[30742] <= 16'b0000_0000_0000_0000;
array[30743] <= 16'b0000_0000_0000_0000;
array[30744] <= 16'b0000_0000_0000_0000;
array[30745] <= 16'b0000_0000_0000_0000;
array[30746] <= 16'b0000_0000_0000_0000;
array[30747] <= 16'b0000_0000_0000_0000;
array[30748] <= 16'b0000_0000_0000_0000;
array[30749] <= 16'b0000_0000_0000_0000;
array[30750] <= 16'b0000_0000_0000_0000;
array[30751] <= 16'b0000_0000_0000_0000;
array[30752] <= 16'b0000_0000_0000_0000;
array[30753] <= 16'b0000_0000_0000_0000;
array[30754] <= 16'b0000_0000_0000_0000;
array[30755] <= 16'b0000_0000_0000_0000;
array[30756] <= 16'b0000_0000_0000_0000;
array[30757] <= 16'b0000_0000_0000_0000;
array[30758] <= 16'b0000_0000_0000_0000;
array[30759] <= 16'b0000_0000_0000_0000;
array[30760] <= 16'b0000_0000_0000_0000;
array[30761] <= 16'b0000_0000_0000_0000;
array[30762] <= 16'b0000_0000_0000_0000;
array[30763] <= 16'b0000_0000_0000_0000;
array[30764] <= 16'b0000_0000_0000_0000;
array[30765] <= 16'b0000_0000_0000_0000;
array[30766] <= 16'b0000_0000_0000_0000;
array[30767] <= 16'b0000_0000_0000_0000;
array[30768] <= 16'b0000_0000_0000_0000;
array[30769] <= 16'b0000_0000_0000_0000;
array[30770] <= 16'b0000_0000_0000_0000;
array[30771] <= 16'b0000_0000_0000_0000;
array[30772] <= 16'b0000_0000_0000_0000;
array[30773] <= 16'b0000_0000_0000_0000;
array[30774] <= 16'b0000_0000_0000_0000;
array[30775] <= 16'b0000_0000_0000_0000;
array[30776] <= 16'b0000_0000_0000_0000;
array[30777] <= 16'b0000_0000_0000_0000;
array[30778] <= 16'b0000_0000_0000_0000;
array[30779] <= 16'b0000_0000_0000_0000;
array[30780] <= 16'b0000_0000_0000_0000;
array[30781] <= 16'b0000_0000_0000_0000;
array[30782] <= 16'b0000_0000_0000_0000;
array[30783] <= 16'b0000_0000_0000_0000;
array[30784] <= 16'b0000_0000_0000_0000;
array[30785] <= 16'b0000_0000_0000_0000;
array[30786] <= 16'b0000_0000_0000_0000;
array[30787] <= 16'b0000_0000_0000_0000;
array[30788] <= 16'b0000_0000_0000_0000;
array[30789] <= 16'b0000_0000_0000_0000;
array[30790] <= 16'b0000_0000_0000_0000;
array[30791] <= 16'b0000_0000_0000_0000;
array[30792] <= 16'b0000_0000_0000_0000;
array[30793] <= 16'b0000_0000_0000_0000;
array[30794] <= 16'b0000_0000_0000_0000;
array[30795] <= 16'b0000_0000_0000_0000;
array[30796] <= 16'b0000_0000_0000_0000;
array[30797] <= 16'b0000_0000_0000_0000;
array[30798] <= 16'b0000_0000_0000_0000;
array[30799] <= 16'b0000_0000_0000_0000;
array[30800] <= 16'b0000_0000_0000_0000;
array[30801] <= 16'b0000_0000_0000_0000;
array[30802] <= 16'b0000_0000_0000_0000;
array[30803] <= 16'b0000_0000_0000_0000;
array[30804] <= 16'b0000_0000_0000_0000;
array[30805] <= 16'b0000_0000_0000_0000;
array[30806] <= 16'b0000_0000_0000_0000;
array[30807] <= 16'b0000_0000_0000_0000;
array[30808] <= 16'b0000_0000_0000_0000;
array[30809] <= 16'b0000_0000_0000_0000;
array[30810] <= 16'b0000_0000_0000_0000;
array[30811] <= 16'b0000_0000_0000_0000;
array[30812] <= 16'b0000_0000_0000_0000;
array[30813] <= 16'b0000_0000_0000_0000;
array[30814] <= 16'b0000_0000_0000_0000;
array[30815] <= 16'b0000_0000_0000_0000;
array[30816] <= 16'b0000_0000_0000_0000;
array[30817] <= 16'b0000_0000_0000_0000;
array[30818] <= 16'b0000_0000_0000_0000;
array[30819] <= 16'b0000_0000_0000_0000;
array[30820] <= 16'b0000_0000_0000_0000;
array[30821] <= 16'b0000_0000_0000_0000;
array[30822] <= 16'b0000_0000_0000_0000;
array[30823] <= 16'b0000_0000_0000_0000;
array[30824] <= 16'b0000_0000_0000_0000;
array[30825] <= 16'b0000_0000_0000_0000;
array[30826] <= 16'b0000_0000_0000_0000;
array[30827] <= 16'b0000_0000_0000_0000;
array[30828] <= 16'b0000_0000_0000_0000;
array[30829] <= 16'b0000_0000_0000_0000;
array[30830] <= 16'b0000_0000_0000_0000;
array[30831] <= 16'b0000_0000_0000_0000;
array[30832] <= 16'b0000_0000_0000_0000;
array[30833] <= 16'b0000_0000_0000_0000;
array[30834] <= 16'b0000_0000_0000_0000;
array[30835] <= 16'b0000_0000_0000_0000;
array[30836] <= 16'b0000_0000_0000_0000;
array[30837] <= 16'b0000_0000_0000_0000;
array[30838] <= 16'b0000_0000_0000_0000;
array[30839] <= 16'b0000_0000_0000_0000;
array[30840] <= 16'b0000_0000_0000_0000;
array[30841] <= 16'b0000_0000_0000_0000;
array[30842] <= 16'b0000_0000_0000_0000;
array[30843] <= 16'b0000_0000_0000_0000;
array[30844] <= 16'b0000_0000_0000_0000;
array[30845] <= 16'b0000_0000_0000_0000;
array[30846] <= 16'b0000_0000_0000_0000;
array[30847] <= 16'b0000_0000_0000_0000;
array[30848] <= 16'b0000_0000_0000_0000;
array[30849] <= 16'b0000_0000_0000_0000;
array[30850] <= 16'b0000_0000_0000_0000;
array[30851] <= 16'b0000_0000_0000_0000;
array[30852] <= 16'b0000_0000_0000_0000;
array[30853] <= 16'b0000_0000_0000_0000;
array[30854] <= 16'b0000_0000_0000_0000;
array[30855] <= 16'b0000_0000_0000_0000;
array[30856] <= 16'b0000_0000_0000_0000;
array[30857] <= 16'b0000_0000_0000_0000;
array[30858] <= 16'b0000_0000_0000_0000;
array[30859] <= 16'b0000_0000_0000_0000;
array[30860] <= 16'b0000_0000_0000_0000;
array[30861] <= 16'b0000_0000_0000_0000;
array[30862] <= 16'b0000_0000_0000_0000;
array[30863] <= 16'b0000_0000_0000_0000;
array[30864] <= 16'b0000_0000_0000_0000;
array[30865] <= 16'b0000_0000_0000_0000;
array[30866] <= 16'b0000_0000_0000_0000;
array[30867] <= 16'b0000_0000_0000_0000;
array[30868] <= 16'b0000_0000_0000_0000;
array[30869] <= 16'b0000_0000_0000_0000;
array[30870] <= 16'b0000_0000_0000_0000;
array[30871] <= 16'b0000_0000_0000_0000;
array[30872] <= 16'b0000_0000_0000_0000;
array[30873] <= 16'b0000_0000_0000_0000;
array[30874] <= 16'b0000_0000_0000_0000;
array[30875] <= 16'b0000_0000_0000_0000;
array[30876] <= 16'b0000_0000_0000_0000;
array[30877] <= 16'b0000_0000_0000_0000;
array[30878] <= 16'b0000_0000_0000_0000;
array[30879] <= 16'b0000_0000_0000_0000;
array[30880] <= 16'b0000_0000_0000_0000;
array[30881] <= 16'b0000_0000_0000_0000;
array[30882] <= 16'b0000_0000_0000_0000;
array[30883] <= 16'b0000_0000_0000_0000;
array[30884] <= 16'b0000_0000_0000_0000;
array[30885] <= 16'b0000_0000_0000_0000;
array[30886] <= 16'b0000_0000_0000_0000;
array[30887] <= 16'b0000_0000_0000_0000;
array[30888] <= 16'b0000_0000_0000_0000;
array[30889] <= 16'b0000_0000_0000_0000;
array[30890] <= 16'b0000_0000_0000_0000;
array[30891] <= 16'b0000_0000_0000_0000;
array[30892] <= 16'b0000_0000_0000_0000;
array[30893] <= 16'b0000_0000_0000_0000;
array[30894] <= 16'b0000_0000_0000_0000;
array[30895] <= 16'b0000_0000_0000_0000;
array[30896] <= 16'b0000_0000_0000_0000;
array[30897] <= 16'b0000_0000_0000_0000;
array[30898] <= 16'b0000_0000_0000_0000;
array[30899] <= 16'b0000_0000_0000_0000;
array[30900] <= 16'b0000_0000_0000_0000;
array[30901] <= 16'b0000_0000_0000_0000;
array[30902] <= 16'b0000_0000_0000_0000;
array[30903] <= 16'b0000_0000_0000_0000;
array[30904] <= 16'b0000_0000_0000_0000;
array[30905] <= 16'b0000_0000_0000_0000;
array[30906] <= 16'b0000_0000_0000_0000;
array[30907] <= 16'b0000_0000_0000_0000;
array[30908] <= 16'b0000_0000_0000_0000;
array[30909] <= 16'b0000_0000_0000_0000;
array[30910] <= 16'b0000_0000_0000_0000;
array[30911] <= 16'b0000_0000_0000_0000;
array[30912] <= 16'b0000_0000_0000_0000;
array[30913] <= 16'b0000_0000_0000_0000;
array[30914] <= 16'b0000_0000_0000_0000;
array[30915] <= 16'b0000_0000_0000_0000;
array[30916] <= 16'b0000_0000_0000_0000;
array[30917] <= 16'b0000_0000_0000_0000;
array[30918] <= 16'b0000_0000_0000_0000;
array[30919] <= 16'b0000_0000_0000_0000;
array[30920] <= 16'b0000_0000_0000_0000;
array[30921] <= 16'b0000_0000_0000_0000;
array[30922] <= 16'b0000_0000_0000_0000;
array[30923] <= 16'b0000_0000_0000_0000;
array[30924] <= 16'b0000_0000_0000_0000;
array[30925] <= 16'b0000_0000_0000_0000;
array[30926] <= 16'b0000_0000_0000_0000;
array[30927] <= 16'b0000_0000_0000_0000;
array[30928] <= 16'b0000_0000_0000_0000;
array[30929] <= 16'b0000_0000_0000_0000;
array[30930] <= 16'b0000_0000_0000_0000;
array[30931] <= 16'b0000_0000_0000_0000;
array[30932] <= 16'b0000_0000_0000_0000;
array[30933] <= 16'b0000_0000_0000_0000;
array[30934] <= 16'b0000_0000_0000_0000;
array[30935] <= 16'b0000_0000_0000_0000;
array[30936] <= 16'b0000_0000_0000_0000;
array[30937] <= 16'b0000_0000_0000_0000;
array[30938] <= 16'b0000_0000_0000_0000;
array[30939] <= 16'b0000_0000_0000_0000;
array[30940] <= 16'b0000_0000_0000_0000;
array[30941] <= 16'b0000_0000_0000_0000;
array[30942] <= 16'b0000_0000_0000_0000;
array[30943] <= 16'b0000_0000_0000_0000;
array[30944] <= 16'b0000_0000_0000_0000;
array[30945] <= 16'b0000_0000_0000_0000;
array[30946] <= 16'b0000_0000_0000_0000;
array[30947] <= 16'b0000_0000_0000_0000;
array[30948] <= 16'b0000_0000_0000_0000;
array[30949] <= 16'b0000_0000_0000_0000;
array[30950] <= 16'b0000_0000_0000_0000;
array[30951] <= 16'b0000_0000_0000_0000;
array[30952] <= 16'b0000_0000_0000_0000;
array[30953] <= 16'b0000_0000_0000_0000;
array[30954] <= 16'b0000_0000_0000_0000;
array[30955] <= 16'b0000_0000_0000_0000;
array[30956] <= 16'b0000_0000_0000_0000;
array[30957] <= 16'b0000_0000_0000_0000;
array[30958] <= 16'b0000_0000_0000_0000;
array[30959] <= 16'b0000_0000_0000_0000;
array[30960] <= 16'b0000_0000_0000_0000;
array[30961] <= 16'b0000_0000_0000_0000;
array[30962] <= 16'b0000_0000_0000_0000;
array[30963] <= 16'b0000_0000_0000_0000;
array[30964] <= 16'b0000_0000_0000_0000;
array[30965] <= 16'b0000_0000_0000_0000;
array[30966] <= 16'b0000_0000_0000_0000;
array[30967] <= 16'b0000_0000_0000_0000;
array[30968] <= 16'b0000_0000_0000_0000;
array[30969] <= 16'b0000_0000_0000_0000;
array[30970] <= 16'b0000_0000_0000_0000;
array[30971] <= 16'b0000_0000_0000_0000;
array[30972] <= 16'b0000_0000_0000_0000;
array[30973] <= 16'b0000_0000_0000_0000;
array[30974] <= 16'b0000_0000_0000_0000;
array[30975] <= 16'b0000_0000_0000_0000;
array[30976] <= 16'b0000_0000_0000_0000;
array[30977] <= 16'b0000_0000_0000_0000;
array[30978] <= 16'b0000_0000_0000_0000;
array[30979] <= 16'b0000_0000_0000_0000;
array[30980] <= 16'b0000_0000_0000_0000;
array[30981] <= 16'b0000_0000_0000_0000;
array[30982] <= 16'b0000_0000_0000_0000;
array[30983] <= 16'b0000_0000_0000_0000;
array[30984] <= 16'b0000_0000_0000_0000;
array[30985] <= 16'b0000_0000_0000_0000;
array[30986] <= 16'b0000_0000_0000_0000;
array[30987] <= 16'b0000_0000_0000_0000;
array[30988] <= 16'b0000_0000_0000_0000;
array[30989] <= 16'b0000_0000_0000_0000;
array[30990] <= 16'b0000_0000_0000_0000;
array[30991] <= 16'b0000_0000_0000_0000;
array[30992] <= 16'b0000_0000_0000_0000;
array[30993] <= 16'b0000_0000_0000_0000;
array[30994] <= 16'b0000_0000_0000_0000;
array[30995] <= 16'b0000_0000_0000_0000;
array[30996] <= 16'b0000_0000_0000_0000;
array[30997] <= 16'b0000_0000_0000_0000;
array[30998] <= 16'b0000_0000_0000_0000;
array[30999] <= 16'b0000_0000_0000_0000;
array[31000] <= 16'b0000_0000_0000_0000;
array[31001] <= 16'b0000_0000_0000_0000;
array[31002] <= 16'b0000_0000_0000_0000;
array[31003] <= 16'b0000_0000_0000_0000;
array[31004] <= 16'b0000_0000_0000_0000;
array[31005] <= 16'b0000_0000_0000_0000;
array[31006] <= 16'b0000_0000_0000_0000;
array[31007] <= 16'b0000_0000_0000_0000;
array[31008] <= 16'b0000_0000_0000_0000;
array[31009] <= 16'b0000_0000_0000_0000;
array[31010] <= 16'b0000_0000_0000_0000;
array[31011] <= 16'b0000_0000_0000_0000;
array[31012] <= 16'b0000_0000_0000_0000;
array[31013] <= 16'b0000_0000_0000_0000;
array[31014] <= 16'b0000_0000_0000_0000;
array[31015] <= 16'b0000_0000_0000_0000;
array[31016] <= 16'b0000_0000_0000_0000;
array[31017] <= 16'b0000_0000_0000_0000;
array[31018] <= 16'b0000_0000_0000_0000;
array[31019] <= 16'b0000_0000_0000_0000;
array[31020] <= 16'b0000_0000_0000_0000;
array[31021] <= 16'b0000_0000_0000_0000;
array[31022] <= 16'b0000_0000_0000_0000;
array[31023] <= 16'b0000_0000_0000_0000;
array[31024] <= 16'b0000_0000_0000_0000;
array[31025] <= 16'b0000_0000_0000_0000;
array[31026] <= 16'b0000_0000_0000_0000;
array[31027] <= 16'b0000_0000_0000_0000;
array[31028] <= 16'b0000_0000_0000_0000;
array[31029] <= 16'b0000_0000_0000_0000;
array[31030] <= 16'b0000_0000_0000_0000;
array[31031] <= 16'b0000_0000_0000_0000;
array[31032] <= 16'b0000_0000_0000_0000;
array[31033] <= 16'b0000_0000_0000_0000;
array[31034] <= 16'b0000_0000_0000_0000;
array[31035] <= 16'b0000_0000_0000_0000;
array[31036] <= 16'b0000_0000_0000_0000;
array[31037] <= 16'b0000_0000_0000_0000;
array[31038] <= 16'b0000_0000_0000_0000;
array[31039] <= 16'b0000_0000_0000_0000;
array[31040] <= 16'b0000_0000_0000_0000;
array[31041] <= 16'b0000_0000_0000_0000;
array[31042] <= 16'b0000_0000_0000_0000;
array[31043] <= 16'b0000_0000_0000_0000;
array[31044] <= 16'b0000_0000_0000_0000;
array[31045] <= 16'b0000_0000_0000_0000;
array[31046] <= 16'b0000_0000_0000_0000;
array[31047] <= 16'b0000_0000_0000_0000;
array[31048] <= 16'b0000_0000_0000_0000;
array[31049] <= 16'b0000_0000_0000_0000;
array[31050] <= 16'b0000_0000_0000_0000;
array[31051] <= 16'b0000_0000_0000_0000;
array[31052] <= 16'b0000_0000_0000_0000;
array[31053] <= 16'b0000_0000_0000_0000;
array[31054] <= 16'b0000_0000_0000_0000;
array[31055] <= 16'b0000_0000_0000_0000;
array[31056] <= 16'b0000_0000_0000_0000;
array[31057] <= 16'b0000_0000_0000_0000;
array[31058] <= 16'b0000_0000_0000_0000;
array[31059] <= 16'b0000_0000_0000_0000;
array[31060] <= 16'b0000_0000_0000_0000;
array[31061] <= 16'b0000_0000_0000_0000;
array[31062] <= 16'b0000_0000_0000_0000;
array[31063] <= 16'b0000_0000_0000_0000;
array[31064] <= 16'b0000_0000_0000_0000;
array[31065] <= 16'b0000_0000_0000_0000;
array[31066] <= 16'b0000_0000_0000_0000;
array[31067] <= 16'b0000_0000_0000_0000;
array[31068] <= 16'b0000_0000_0000_0000;
array[31069] <= 16'b0000_0000_0000_0000;
array[31070] <= 16'b0000_0000_0000_0000;
array[31071] <= 16'b0000_0000_0000_0000;
array[31072] <= 16'b0000_0000_0000_0000;
array[31073] <= 16'b0000_0000_0000_0000;
array[31074] <= 16'b0000_0000_0000_0000;
array[31075] <= 16'b0000_0000_0000_0000;
array[31076] <= 16'b0000_0000_0000_0000;
array[31077] <= 16'b0000_0000_0000_0000;
array[31078] <= 16'b0000_0000_0000_0000;
array[31079] <= 16'b0000_0000_0000_0000;
array[31080] <= 16'b0000_0000_0000_0000;
array[31081] <= 16'b0000_0000_0000_0000;
array[31082] <= 16'b0000_0000_0000_0000;
array[31083] <= 16'b0000_0000_0000_0000;
array[31084] <= 16'b0000_0000_0000_0000;
array[31085] <= 16'b0000_0000_0000_0000;
array[31086] <= 16'b0000_0000_0000_0000;
array[31087] <= 16'b0000_0000_0000_0000;
array[31088] <= 16'b0000_0000_0000_0000;
array[31089] <= 16'b0000_0000_0000_0000;
array[31090] <= 16'b0000_0000_0000_0000;
array[31091] <= 16'b0000_0000_0000_0000;
array[31092] <= 16'b0000_0000_0000_0000;
array[31093] <= 16'b0000_0000_0000_0000;
array[31094] <= 16'b0000_0000_0000_0000;
array[31095] <= 16'b0000_0000_0000_0000;
array[31096] <= 16'b0000_0000_0000_0000;
array[31097] <= 16'b0000_0000_0000_0000;
array[31098] <= 16'b0000_0000_0000_0000;
array[31099] <= 16'b0000_0000_0000_0000;
array[31100] <= 16'b0000_0000_0000_0000;
array[31101] <= 16'b0000_0000_0000_0000;
array[31102] <= 16'b0000_0000_0000_0000;
array[31103] <= 16'b0000_0000_0000_0000;
array[31104] <= 16'b0000_0000_0000_0000;
array[31105] <= 16'b0000_0000_0000_0000;
array[31106] <= 16'b0000_0000_0000_0000;
array[31107] <= 16'b0000_0000_0000_0000;
array[31108] <= 16'b0000_0000_0000_0000;
array[31109] <= 16'b0000_0000_0000_0000;
array[31110] <= 16'b0000_0000_0000_0000;
array[31111] <= 16'b0000_0000_0000_0000;
array[31112] <= 16'b0000_0000_0000_0000;
array[31113] <= 16'b0000_0000_0000_0000;
array[31114] <= 16'b0000_0000_0000_0000;
array[31115] <= 16'b0000_0000_0000_0000;
array[31116] <= 16'b0000_0000_0000_0000;
array[31117] <= 16'b0000_0000_0000_0000;
array[31118] <= 16'b0000_0000_0000_0000;
array[31119] <= 16'b0000_0000_0000_0000;
array[31120] <= 16'b0000_0000_0000_0000;
array[31121] <= 16'b0000_0000_0000_0000;
array[31122] <= 16'b0000_0000_0000_0000;
array[31123] <= 16'b0000_0000_0000_0000;
array[31124] <= 16'b0000_0000_0000_0000;
array[31125] <= 16'b0000_0000_0000_0000;
array[31126] <= 16'b0000_0000_0000_0000;
array[31127] <= 16'b0000_0000_0000_0000;
array[31128] <= 16'b0000_0000_0000_0000;
array[31129] <= 16'b0000_0000_0000_0000;
array[31130] <= 16'b0000_0000_0000_0000;
array[31131] <= 16'b0000_0000_0000_0000;
array[31132] <= 16'b0000_0000_0000_0000;
array[31133] <= 16'b0000_0000_0000_0000;
array[31134] <= 16'b0000_0000_0000_0000;
array[31135] <= 16'b0000_0000_0000_0000;
array[31136] <= 16'b0000_0000_0000_0000;
array[31137] <= 16'b0000_0000_0000_0000;
array[31138] <= 16'b0000_0000_0000_0000;
array[31139] <= 16'b0000_0000_0000_0000;
array[31140] <= 16'b0000_0000_0000_0000;
array[31141] <= 16'b0000_0000_0000_0000;
array[31142] <= 16'b0000_0000_0000_0000;
array[31143] <= 16'b0000_0000_0000_0000;
array[31144] <= 16'b0000_0000_0000_0000;
array[31145] <= 16'b0000_0000_0000_0000;
array[31146] <= 16'b0000_0000_0000_0000;
array[31147] <= 16'b0000_0000_0000_0000;
array[31148] <= 16'b0000_0000_0000_0000;
array[31149] <= 16'b0000_0000_0000_0000;
array[31150] <= 16'b0000_0000_0000_0000;
array[31151] <= 16'b0000_0000_0000_0000;
array[31152] <= 16'b0000_0000_0000_0000;
array[31153] <= 16'b0000_0000_0000_0000;
array[31154] <= 16'b0000_0000_0000_0000;
array[31155] <= 16'b0000_0000_0000_0000;
array[31156] <= 16'b0000_0000_0000_0000;
array[31157] <= 16'b0000_0000_0000_0000;
array[31158] <= 16'b0000_0000_0000_0000;
array[31159] <= 16'b0000_0000_0000_0000;
array[31160] <= 16'b0000_0000_0000_0000;
array[31161] <= 16'b0000_0000_0000_0000;
array[31162] <= 16'b0000_0000_0000_0000;
array[31163] <= 16'b0000_0000_0000_0000;
array[31164] <= 16'b0000_0000_0000_0000;
array[31165] <= 16'b0000_0000_0000_0000;
array[31166] <= 16'b0000_0000_0000_0000;
array[31167] <= 16'b0000_0000_0000_0000;
array[31168] <= 16'b0000_0000_0000_0000;
array[31169] <= 16'b0000_0000_0000_0000;
array[31170] <= 16'b0000_0000_0000_0000;
array[31171] <= 16'b0000_0000_0000_0000;
array[31172] <= 16'b0000_0000_0000_0000;
array[31173] <= 16'b0000_0000_0000_0000;
array[31174] <= 16'b0000_0000_0000_0000;
array[31175] <= 16'b0000_0000_0000_0000;
array[31176] <= 16'b0000_0000_0000_0000;
array[31177] <= 16'b0000_0000_0000_0000;
array[31178] <= 16'b0000_0000_0000_0000;
array[31179] <= 16'b0000_0000_0000_0000;
array[31180] <= 16'b0000_0000_0000_0000;
array[31181] <= 16'b0000_0000_0000_0000;
array[31182] <= 16'b0000_0000_0000_0000;
array[31183] <= 16'b0000_0000_0000_0000;
array[31184] <= 16'b0000_0000_0000_0000;
array[31185] <= 16'b0000_0000_0000_0000;
array[31186] <= 16'b0000_0000_0000_0000;
array[31187] <= 16'b0000_0000_0000_0000;
array[31188] <= 16'b0000_0000_0000_0000;
array[31189] <= 16'b0000_0000_0000_0000;
array[31190] <= 16'b0000_0000_0000_0000;
array[31191] <= 16'b0000_0000_0000_0000;
array[31192] <= 16'b0000_0000_0000_0000;
array[31193] <= 16'b0000_0000_0000_0000;
array[31194] <= 16'b0000_0000_0000_0000;
array[31195] <= 16'b0000_0000_0000_0000;
array[31196] <= 16'b0000_0000_0000_0000;
array[31197] <= 16'b0000_0000_0000_0000;
array[31198] <= 16'b0000_0000_0000_0000;
array[31199] <= 16'b0000_0000_0000_0000;
array[31200] <= 16'b0000_0000_0000_0000;
array[31201] <= 16'b0000_0000_0000_0000;
array[31202] <= 16'b0000_0000_0000_0000;
array[31203] <= 16'b0000_0000_0000_0000;
array[31204] <= 16'b0000_0000_0000_0000;
array[31205] <= 16'b0000_0000_0000_0000;
array[31206] <= 16'b0000_0000_0000_0000;
array[31207] <= 16'b0000_0000_0000_0000;
array[31208] <= 16'b0000_0000_0000_0000;
array[31209] <= 16'b0000_0000_0000_0000;
array[31210] <= 16'b0000_0000_0000_0000;
array[31211] <= 16'b0000_0000_0000_0000;
array[31212] <= 16'b0000_0000_0000_0000;
array[31213] <= 16'b0000_0000_0000_0000;
array[31214] <= 16'b0000_0000_0000_0000;
array[31215] <= 16'b0000_0000_0000_0000;
array[31216] <= 16'b0000_0000_0000_0000;
array[31217] <= 16'b0000_0000_0000_0000;
array[31218] <= 16'b0000_0000_0000_0000;
array[31219] <= 16'b0000_0000_0000_0000;
array[31220] <= 16'b0000_0000_0000_0000;
array[31221] <= 16'b0000_0000_0000_0000;
array[31222] <= 16'b0000_0000_0000_0000;
array[31223] <= 16'b0000_0000_0000_0000;
array[31224] <= 16'b0000_0000_0000_0000;
array[31225] <= 16'b0000_0000_0000_0000;
array[31226] <= 16'b0000_0000_0000_0000;
array[31227] <= 16'b0000_0000_0000_0000;
array[31228] <= 16'b0000_0000_0000_0000;
array[31229] <= 16'b0000_0000_0000_0000;
array[31230] <= 16'b0000_0000_0000_0000;
array[31231] <= 16'b0000_0000_0000_0000;
array[31232] <= 16'b0000_0000_0000_0000;
array[31233] <= 16'b0000_0000_0000_0000;
array[31234] <= 16'b0000_0000_0000_0000;
array[31235] <= 16'b0000_0000_0000_0000;
array[31236] <= 16'b0000_0000_0000_0000;
array[31237] <= 16'b0000_0000_0000_0000;
array[31238] <= 16'b0000_0000_0000_0000;
array[31239] <= 16'b0000_0000_0000_0000;
array[31240] <= 16'b0000_0000_0000_0000;
array[31241] <= 16'b0000_0000_0000_0000;
array[31242] <= 16'b0000_0000_0000_0000;
array[31243] <= 16'b0000_0000_0000_0000;
array[31244] <= 16'b0000_0000_0000_0000;
array[31245] <= 16'b0000_0000_0000_0000;
array[31246] <= 16'b0000_0000_0000_0000;
array[31247] <= 16'b0000_0000_0000_0000;
array[31248] <= 16'b0000_0000_0000_0000;
array[31249] <= 16'b0000_0000_0000_0000;
array[31250] <= 16'b0000_0000_0000_0000;
array[31251] <= 16'b0000_0000_0000_0000;
array[31252] <= 16'b0000_0000_0000_0000;
array[31253] <= 16'b0000_0000_0000_0000;
array[31254] <= 16'b0000_0000_0000_0000;
array[31255] <= 16'b0000_0000_0000_0000;
array[31256] <= 16'b0000_0000_0000_0000;
array[31257] <= 16'b0000_0000_0000_0000;
array[31258] <= 16'b0000_0000_0000_0000;
array[31259] <= 16'b0000_0000_0000_0000;
array[31260] <= 16'b0000_0000_0000_0000;
array[31261] <= 16'b0000_0000_0000_0000;
array[31262] <= 16'b0000_0000_0000_0000;
array[31263] <= 16'b0000_0000_0000_0000;
array[31264] <= 16'b0000_0000_0000_0000;
array[31265] <= 16'b0000_0000_0000_0000;
array[31266] <= 16'b0000_0000_0000_0000;
array[31267] <= 16'b0000_0000_0000_0000;
array[31268] <= 16'b0000_0000_0000_0000;
array[31269] <= 16'b0000_0000_0000_0000;
array[31270] <= 16'b0000_0000_0000_0000;
array[31271] <= 16'b0000_0000_0000_0000;
array[31272] <= 16'b0000_0000_0000_0000;
array[31273] <= 16'b0000_0000_0000_0000;
array[31274] <= 16'b0000_0000_0000_0000;
array[31275] <= 16'b0000_0000_0000_0000;
array[31276] <= 16'b0000_0000_0000_0000;
array[31277] <= 16'b0000_0000_0000_0000;
array[31278] <= 16'b0000_0000_0000_0000;
array[31279] <= 16'b0000_0000_0000_0000;
array[31280] <= 16'b0000_0000_0000_0000;
array[31281] <= 16'b0000_0000_0000_0000;
array[31282] <= 16'b0000_0000_0000_0000;
array[31283] <= 16'b0000_0000_0000_0000;
array[31284] <= 16'b0000_0000_0000_0000;
array[31285] <= 16'b0000_0000_0000_0000;
array[31286] <= 16'b0000_0000_0000_0000;
array[31287] <= 16'b0000_0000_0000_0000;
array[31288] <= 16'b0000_0000_0000_0000;
array[31289] <= 16'b0000_0000_0000_0000;
array[31290] <= 16'b0000_0000_0000_0000;
array[31291] <= 16'b0000_0000_0000_0000;
array[31292] <= 16'b0000_0000_0000_0000;
array[31293] <= 16'b0000_0000_0000_0000;
array[31294] <= 16'b0000_0000_0000_0000;
array[31295] <= 16'b0000_0000_0000_0000;
array[31296] <= 16'b0000_0000_0000_0000;
array[31297] <= 16'b0000_0000_0000_0000;
array[31298] <= 16'b0000_0000_0000_0000;
array[31299] <= 16'b0000_0000_0000_0000;
array[31300] <= 16'b0000_0000_0000_0000;
array[31301] <= 16'b0000_0000_0000_0000;
array[31302] <= 16'b0000_0000_0000_0000;
array[31303] <= 16'b0000_0000_0000_0000;
array[31304] <= 16'b0000_0000_0000_0000;
array[31305] <= 16'b0000_0000_0000_0000;
array[31306] <= 16'b0000_0000_0000_0000;
array[31307] <= 16'b0000_0000_0000_0000;
array[31308] <= 16'b0000_0000_0000_0000;
array[31309] <= 16'b0000_0000_0000_0000;
array[31310] <= 16'b0000_0000_0000_0000;
array[31311] <= 16'b0000_0000_0000_0000;
array[31312] <= 16'b0000_0000_0000_0000;
array[31313] <= 16'b0000_0000_0000_0000;
array[31314] <= 16'b0000_0000_0000_0000;
array[31315] <= 16'b0000_0000_0000_0000;
array[31316] <= 16'b0000_0000_0000_0000;
array[31317] <= 16'b0000_0000_0000_0000;
array[31318] <= 16'b0000_0000_0000_0000;
array[31319] <= 16'b0000_0000_0000_0000;
array[31320] <= 16'b0000_0000_0000_0000;
array[31321] <= 16'b0000_0000_0000_0000;
array[31322] <= 16'b0000_0000_0000_0000;
array[31323] <= 16'b0000_0000_0000_0000;
array[31324] <= 16'b0000_0000_0000_0000;
array[31325] <= 16'b0000_0000_0000_0000;
array[31326] <= 16'b0000_0000_0000_0000;
array[31327] <= 16'b0000_0000_0000_0000;
array[31328] <= 16'b0000_0000_0000_0000;
array[31329] <= 16'b0000_0000_0000_0000;
array[31330] <= 16'b0000_0000_0000_0000;
array[31331] <= 16'b0000_0000_0000_0000;
array[31332] <= 16'b0000_0000_0000_0000;
array[31333] <= 16'b0000_0000_0000_0000;
array[31334] <= 16'b0000_0000_0000_0000;
array[31335] <= 16'b0000_0000_0000_0000;
array[31336] <= 16'b0000_0000_0000_0000;
array[31337] <= 16'b0000_0000_0000_0000;
array[31338] <= 16'b0000_0000_0000_0000;
array[31339] <= 16'b0000_0000_0000_0000;
array[31340] <= 16'b0000_0000_0000_0000;
array[31341] <= 16'b0000_0000_0000_0000;
array[31342] <= 16'b0000_0000_0000_0000;
array[31343] <= 16'b0000_0000_0000_0000;
array[31344] <= 16'b0000_0000_0000_0000;
array[31345] <= 16'b0000_0000_0000_0000;
array[31346] <= 16'b0000_0000_0000_0000;
array[31347] <= 16'b0000_0000_0000_0000;
array[31348] <= 16'b0000_0000_0000_0000;
array[31349] <= 16'b0000_0000_0000_0000;
array[31350] <= 16'b0000_0000_0000_0000;
array[31351] <= 16'b0000_0000_0000_0000;
array[31352] <= 16'b0000_0000_0000_0000;
array[31353] <= 16'b0000_0000_0000_0000;
array[31354] <= 16'b0000_0000_0000_0000;
array[31355] <= 16'b0000_0000_0000_0000;
array[31356] <= 16'b0000_0000_0000_0000;
array[31357] <= 16'b0000_0000_0000_0000;
array[31358] <= 16'b0000_0000_0000_0000;
array[31359] <= 16'b0000_0000_0000_0000;
array[31360] <= 16'b0000_0000_0000_0000;
array[31361] <= 16'b0000_0000_0000_0000;
array[31362] <= 16'b0000_0000_0000_0000;
array[31363] <= 16'b0000_0000_0000_0000;
array[31364] <= 16'b0000_0000_0000_0000;
array[31365] <= 16'b0000_0000_0000_0000;
array[31366] <= 16'b0000_0000_0000_0000;
array[31367] <= 16'b0000_0000_0000_0000;
array[31368] <= 16'b0000_0000_0000_0000;
array[31369] <= 16'b0000_0000_0000_0000;
array[31370] <= 16'b0000_0000_0000_0000;
array[31371] <= 16'b0000_0000_0000_0000;
array[31372] <= 16'b0000_0000_0000_0000;
array[31373] <= 16'b0000_0000_0000_0000;
array[31374] <= 16'b0000_0000_0000_0000;
array[31375] <= 16'b0000_0000_0000_0000;
array[31376] <= 16'b0000_0000_0000_0000;
array[31377] <= 16'b0000_0000_0000_0000;
array[31378] <= 16'b0000_0000_0000_0000;
array[31379] <= 16'b0000_0000_0000_0000;
array[31380] <= 16'b0000_0000_0000_0000;
array[31381] <= 16'b0000_0000_0000_0000;
array[31382] <= 16'b0000_0000_0000_0000;
array[31383] <= 16'b0000_0000_0000_0000;
array[31384] <= 16'b0000_0000_0000_0000;
array[31385] <= 16'b0000_0000_0000_0000;
array[31386] <= 16'b0000_0000_0000_0000;
array[31387] <= 16'b0000_0000_0000_0000;
array[31388] <= 16'b0000_0000_0000_0000;
array[31389] <= 16'b0000_0000_0000_0000;
array[31390] <= 16'b0000_0000_0000_0000;
array[31391] <= 16'b0000_0000_0000_0000;
array[31392] <= 16'b0000_0000_0000_0000;
array[31393] <= 16'b0000_0000_0000_0000;
array[31394] <= 16'b0000_0000_0000_0000;
array[31395] <= 16'b0000_0000_0000_0000;
array[31396] <= 16'b0000_0000_0000_0000;
array[31397] <= 16'b0000_0000_0000_0000;
array[31398] <= 16'b0000_0000_0000_0000;
array[31399] <= 16'b0000_0000_0000_0000;
array[31400] <= 16'b0000_0000_0000_0000;
array[31401] <= 16'b0000_0000_0000_0000;
array[31402] <= 16'b0000_0000_0000_0000;
array[31403] <= 16'b0000_0000_0000_0000;
array[31404] <= 16'b0000_0000_0000_0000;
array[31405] <= 16'b0000_0000_0000_0000;
array[31406] <= 16'b0000_0000_0000_0000;
array[31407] <= 16'b0000_0000_0000_0000;
array[31408] <= 16'b0000_0000_0000_0000;
array[31409] <= 16'b0000_0000_0000_0000;
array[31410] <= 16'b0000_0000_0000_0000;
array[31411] <= 16'b0000_0000_0000_0000;
array[31412] <= 16'b0000_0000_0000_0000;
array[31413] <= 16'b0000_0000_0000_0000;
array[31414] <= 16'b0000_0000_0000_0000;
array[31415] <= 16'b0000_0000_0000_0000;
array[31416] <= 16'b0000_0000_0000_0000;
array[31417] <= 16'b0000_0000_0000_0000;
array[31418] <= 16'b0000_0000_0000_0000;
array[31419] <= 16'b0000_0000_0000_0000;
array[31420] <= 16'b0000_0000_0000_0000;
array[31421] <= 16'b0000_0000_0000_0000;
array[31422] <= 16'b0000_0000_0000_0000;
array[31423] <= 16'b0000_0000_0000_0000;
array[31424] <= 16'b0000_0000_0000_0000;
array[31425] <= 16'b0000_0000_0000_0000;
array[31426] <= 16'b0000_0000_0000_0000;
array[31427] <= 16'b0000_0000_0000_0000;
array[31428] <= 16'b0000_0000_0000_0000;
array[31429] <= 16'b0000_0000_0000_0000;
array[31430] <= 16'b0000_0000_0000_0000;
array[31431] <= 16'b0000_0000_0000_0000;
array[31432] <= 16'b0000_0000_0000_0000;
array[31433] <= 16'b0000_0000_0000_0000;
array[31434] <= 16'b0000_0000_0000_0000;
array[31435] <= 16'b0000_0000_0000_0000;
array[31436] <= 16'b0000_0000_0000_0000;
array[31437] <= 16'b0000_0000_0000_0000;
array[31438] <= 16'b0000_0000_0000_0000;
array[31439] <= 16'b0000_0000_0000_0000;
array[31440] <= 16'b0000_0000_0000_0000;
array[31441] <= 16'b0000_0000_0000_0000;
array[31442] <= 16'b0000_0000_0000_0000;
array[31443] <= 16'b0000_0000_0000_0000;
array[31444] <= 16'b0000_0000_0000_0000;
array[31445] <= 16'b0000_0000_0000_0000;
array[31446] <= 16'b0000_0000_0000_0000;
array[31447] <= 16'b0000_0000_0000_0000;
array[31448] <= 16'b0000_0000_0000_0000;
array[31449] <= 16'b0000_0000_0000_0000;
array[31450] <= 16'b0000_0000_0000_0000;
array[31451] <= 16'b0000_0000_0000_0000;
array[31452] <= 16'b0000_0000_0000_0000;
array[31453] <= 16'b0000_0000_0000_0000;
array[31454] <= 16'b0000_0000_0000_0000;
array[31455] <= 16'b0000_0000_0000_0000;
array[31456] <= 16'b0000_0000_0000_0000;
array[31457] <= 16'b0000_0000_0000_0000;
array[31458] <= 16'b0000_0000_0000_0000;
array[31459] <= 16'b0000_0000_0000_0000;
array[31460] <= 16'b0000_0000_0000_0000;
array[31461] <= 16'b0000_0000_0000_0000;
array[31462] <= 16'b0000_0000_0000_0000;
array[31463] <= 16'b0000_0000_0000_0000;
array[31464] <= 16'b0000_0000_0000_0000;
array[31465] <= 16'b0000_0000_0000_0000;
array[31466] <= 16'b0000_0000_0000_0000;
array[31467] <= 16'b0000_0000_0000_0000;
array[31468] <= 16'b0000_0000_0000_0000;
array[31469] <= 16'b0000_0000_0000_0000;
array[31470] <= 16'b0000_0000_0000_0000;
array[31471] <= 16'b0000_0000_0000_0000;
array[31472] <= 16'b0000_0000_0000_0000;
array[31473] <= 16'b0000_0000_0000_0000;
array[31474] <= 16'b0000_0000_0000_0000;
array[31475] <= 16'b0000_0000_0000_0000;
array[31476] <= 16'b0000_0000_0000_0000;
array[31477] <= 16'b0000_0000_0000_0000;
array[31478] <= 16'b0000_0000_0000_0000;
array[31479] <= 16'b0000_0000_0000_0000;
array[31480] <= 16'b0000_0000_0000_0000;
array[31481] <= 16'b0000_0000_0000_0000;
array[31482] <= 16'b0000_0000_0000_0000;
array[31483] <= 16'b0000_0000_0000_0000;
array[31484] <= 16'b0000_0000_0000_0000;
array[31485] <= 16'b0000_0000_0000_0000;
array[31486] <= 16'b0000_0000_0000_0000;
array[31487] <= 16'b0000_0000_0000_0000;
array[31488] <= 16'b0000_0000_0000_0000;
array[31489] <= 16'b0000_0000_0000_0000;
array[31490] <= 16'b0000_0000_0000_0000;
array[31491] <= 16'b0000_0000_0000_0000;
array[31492] <= 16'b0000_0000_0000_0000;
array[31493] <= 16'b0000_0000_0000_0000;
array[31494] <= 16'b0000_0000_0000_0000;
array[31495] <= 16'b0000_0000_0000_0000;
array[31496] <= 16'b0000_0000_0000_0000;
array[31497] <= 16'b0000_0000_0000_0000;
array[31498] <= 16'b0000_0000_0000_0000;
array[31499] <= 16'b0000_0000_0000_0000;
array[31500] <= 16'b0000_0000_0000_0000;
array[31501] <= 16'b0000_0000_0000_0000;
array[31502] <= 16'b0000_0000_0000_0000;
array[31503] <= 16'b0000_0000_0000_0000;
array[31504] <= 16'b0000_0000_0000_0000;
array[31505] <= 16'b0000_0000_0000_0000;
array[31506] <= 16'b0000_0000_0000_0000;
array[31507] <= 16'b0000_0000_0000_0000;
array[31508] <= 16'b0000_0000_0000_0000;
array[31509] <= 16'b0000_0000_0000_0000;
array[31510] <= 16'b0000_0000_0000_0000;
array[31511] <= 16'b0000_0000_0000_0000;
array[31512] <= 16'b0000_0000_0000_0000;
array[31513] <= 16'b0000_0000_0000_0000;
array[31514] <= 16'b0000_0000_0000_0000;
array[31515] <= 16'b0000_0000_0000_0000;
array[31516] <= 16'b0000_0000_0000_0000;
array[31517] <= 16'b0000_0000_0000_0000;
array[31518] <= 16'b0000_0000_0000_0000;
array[31519] <= 16'b0000_0000_0000_0000;
array[31520] <= 16'b0000_0000_0000_0000;
array[31521] <= 16'b0000_0000_0000_0000;
array[31522] <= 16'b0000_0000_0000_0000;
array[31523] <= 16'b0000_0000_0000_0000;
array[31524] <= 16'b0000_0000_0000_0000;
array[31525] <= 16'b0000_0000_0000_0000;
array[31526] <= 16'b0000_0000_0000_0000;
array[31527] <= 16'b0000_0000_0000_0000;
array[31528] <= 16'b0000_0000_0000_0000;
array[31529] <= 16'b0000_0000_0000_0000;
array[31530] <= 16'b0000_0000_0000_0000;
array[31531] <= 16'b0000_0000_0000_0000;
array[31532] <= 16'b0000_0000_0000_0000;
array[31533] <= 16'b0000_0000_0000_0000;
array[31534] <= 16'b0000_0000_0000_0000;
array[31535] <= 16'b0000_0000_0000_0000;
array[31536] <= 16'b0000_0000_0000_0000;
array[31537] <= 16'b0000_0000_0000_0000;
array[31538] <= 16'b0000_0000_0000_0000;
array[31539] <= 16'b0000_0000_0000_0000;
array[31540] <= 16'b0000_0000_0000_0000;
array[31541] <= 16'b0000_0000_0000_0000;
array[31542] <= 16'b0000_0000_0000_0000;
array[31543] <= 16'b0000_0000_0000_0000;
array[31544] <= 16'b0000_0000_0000_0000;
array[31545] <= 16'b0000_0000_0000_0000;
array[31546] <= 16'b0000_0000_0000_0000;
array[31547] <= 16'b0000_0000_0000_0000;
array[31548] <= 16'b0000_0000_0000_0000;
array[31549] <= 16'b0000_0000_0000_0000;
array[31550] <= 16'b0000_0000_0000_0000;
array[31551] <= 16'b0000_0000_0000_0000;
array[31552] <= 16'b0000_0000_0000_0000;
array[31553] <= 16'b0000_0000_0000_0000;
array[31554] <= 16'b0000_0000_0000_0000;
array[31555] <= 16'b0000_0000_0000_0000;
array[31556] <= 16'b0000_0000_0000_0000;
array[31557] <= 16'b0000_0000_0000_0000;
array[31558] <= 16'b0000_0000_0000_0000;
array[31559] <= 16'b0000_0000_0000_0000;
array[31560] <= 16'b0000_0000_0000_0000;
array[31561] <= 16'b0000_0000_0000_0000;
array[31562] <= 16'b0000_0000_0000_0000;
array[31563] <= 16'b0000_0000_0000_0000;
array[31564] <= 16'b0000_0000_0000_0000;
array[31565] <= 16'b0000_0000_0000_0000;
array[31566] <= 16'b0000_0000_0000_0000;
array[31567] <= 16'b0000_0000_0000_0000;
array[31568] <= 16'b0000_0000_0000_0000;
array[31569] <= 16'b0000_0000_0000_0000;
array[31570] <= 16'b0000_0000_0000_0000;
array[31571] <= 16'b0000_0000_0000_0000;
array[31572] <= 16'b0000_0000_0000_0000;
array[31573] <= 16'b0000_0000_0000_0000;
array[31574] <= 16'b0000_0000_0000_0000;
array[31575] <= 16'b0000_0000_0000_0000;
array[31576] <= 16'b0000_0000_0000_0000;
array[31577] <= 16'b0000_0000_0000_0000;
array[31578] <= 16'b0000_0000_0000_0000;
array[31579] <= 16'b0000_0000_0000_0000;
array[31580] <= 16'b0000_0000_0000_0000;
array[31581] <= 16'b0000_0000_0000_0000;
array[31582] <= 16'b0000_0000_0000_0000;
array[31583] <= 16'b0000_0000_0000_0000;
array[31584] <= 16'b0000_0000_0000_0000;
array[31585] <= 16'b0000_0000_0000_0000;
array[31586] <= 16'b0000_0000_0000_0000;
array[31587] <= 16'b0000_0000_0000_0000;
array[31588] <= 16'b0000_0000_0000_0000;
array[31589] <= 16'b0000_0000_0000_0000;
array[31590] <= 16'b0000_0000_0000_0000;
array[31591] <= 16'b0000_0000_0000_0000;
array[31592] <= 16'b0000_0000_0000_0000;
array[31593] <= 16'b0000_0000_0000_0000;
array[31594] <= 16'b0000_0000_0000_0000;
array[31595] <= 16'b0000_0000_0000_0000;
array[31596] <= 16'b0000_0000_0000_0000;
array[31597] <= 16'b0000_0000_0000_0000;
array[31598] <= 16'b0000_0000_0000_0000;
array[31599] <= 16'b0000_0000_0000_0000;
array[31600] <= 16'b0000_0000_0000_0000;
array[31601] <= 16'b0000_0000_0000_0000;
array[31602] <= 16'b0000_0000_0000_0000;
array[31603] <= 16'b0000_0000_0000_0000;
array[31604] <= 16'b0000_0000_0000_0000;
array[31605] <= 16'b0000_0000_0000_0000;
array[31606] <= 16'b0000_0000_0000_0000;
array[31607] <= 16'b0000_0000_0000_0000;
array[31608] <= 16'b0000_0000_0000_0000;
array[31609] <= 16'b0000_0000_0000_0000;
array[31610] <= 16'b0000_0000_0000_0000;
array[31611] <= 16'b0000_0000_0000_0000;
array[31612] <= 16'b0000_0000_0000_0000;
array[31613] <= 16'b0000_0000_0000_0000;
array[31614] <= 16'b0000_0000_0000_0000;
array[31615] <= 16'b0000_0000_0000_0000;
array[31616] <= 16'b0000_0000_0000_0000;
array[31617] <= 16'b0000_0000_0000_0000;
array[31618] <= 16'b0000_0000_0000_0000;
array[31619] <= 16'b0000_0000_0000_0000;
array[31620] <= 16'b0000_0000_0000_0000;
array[31621] <= 16'b0000_0000_0000_0000;
array[31622] <= 16'b0000_0000_0000_0000;
array[31623] <= 16'b0000_0000_0000_0000;
array[31624] <= 16'b0000_0000_0000_0000;
array[31625] <= 16'b0000_0000_0000_0000;
array[31626] <= 16'b0000_0000_0000_0000;
array[31627] <= 16'b0000_0000_0000_0000;
array[31628] <= 16'b0000_0000_0000_0000;
array[31629] <= 16'b0000_0000_0000_0000;
array[31630] <= 16'b0000_0000_0000_0000;
array[31631] <= 16'b0000_0000_0000_0000;
array[31632] <= 16'b0000_0000_0000_0000;
array[31633] <= 16'b0000_0000_0000_0000;
array[31634] <= 16'b0000_0000_0000_0000;
array[31635] <= 16'b0000_0000_0000_0000;
array[31636] <= 16'b0000_0000_0000_0000;
array[31637] <= 16'b0000_0000_0000_0000;
array[31638] <= 16'b0000_0000_0000_0000;
array[31639] <= 16'b0000_0000_0000_0000;
array[31640] <= 16'b0000_0000_0000_0000;
array[31641] <= 16'b0000_0000_0000_0000;
array[31642] <= 16'b0000_0000_0000_0000;
array[31643] <= 16'b0000_0000_0000_0000;
array[31644] <= 16'b0000_0000_0000_0000;
array[31645] <= 16'b0000_0000_0000_0000;
array[31646] <= 16'b0000_0000_0000_0000;
array[31647] <= 16'b0000_0000_0000_0000;
array[31648] <= 16'b0000_0000_0000_0000;
array[31649] <= 16'b0000_0000_0000_0000;
array[31650] <= 16'b0000_0000_0000_0000;
array[31651] <= 16'b0000_0000_0000_0000;
array[31652] <= 16'b0000_0000_0000_0000;
array[31653] <= 16'b0000_0000_0000_0000;
array[31654] <= 16'b0000_0000_0000_0000;
array[31655] <= 16'b0000_0000_0000_0000;
array[31656] <= 16'b0000_0000_0000_0000;
array[31657] <= 16'b0000_0000_0000_0000;
array[31658] <= 16'b0000_0000_0000_0000;
array[31659] <= 16'b0000_0000_0000_0000;
array[31660] <= 16'b0000_0000_0000_0000;
array[31661] <= 16'b0000_0000_0000_0000;
array[31662] <= 16'b0000_0000_0000_0000;
array[31663] <= 16'b0000_0000_0000_0000;
array[31664] <= 16'b0000_0000_0000_0000;
array[31665] <= 16'b0000_0000_0000_0000;
array[31666] <= 16'b0000_0000_0000_0000;
array[31667] <= 16'b0000_0000_0000_0000;
array[31668] <= 16'b0000_0000_0000_0000;
array[31669] <= 16'b0000_0000_0000_0000;
array[31670] <= 16'b0000_0000_0000_0000;
array[31671] <= 16'b0000_0000_0000_0000;
array[31672] <= 16'b0000_0000_0000_0000;
array[31673] <= 16'b0000_0000_0000_0000;
array[31674] <= 16'b0000_0000_0000_0000;
array[31675] <= 16'b0000_0000_0000_0000;
array[31676] <= 16'b0000_0000_0000_0000;
array[31677] <= 16'b0000_0000_0000_0000;
array[31678] <= 16'b0000_0000_0000_0000;
array[31679] <= 16'b0000_0000_0000_0000;
array[31680] <= 16'b0000_0000_0000_0000;
array[31681] <= 16'b0000_0000_0000_0000;
array[31682] <= 16'b0000_0000_0000_0000;
array[31683] <= 16'b0000_0000_0000_0000;
array[31684] <= 16'b0000_0000_0000_0000;
array[31685] <= 16'b0000_0000_0000_0000;
array[31686] <= 16'b0000_0000_0000_0000;
array[31687] <= 16'b0000_0000_0000_0000;
array[31688] <= 16'b0000_0000_0000_0000;
array[31689] <= 16'b0000_0000_0000_0000;
array[31690] <= 16'b0000_0000_0000_0000;
array[31691] <= 16'b0000_0000_0000_0000;
array[31692] <= 16'b0000_0000_0000_0000;
array[31693] <= 16'b0000_0000_0000_0000;
array[31694] <= 16'b0000_0000_0000_0000;
array[31695] <= 16'b0000_0000_0000_0000;
array[31696] <= 16'b0000_0000_0000_0000;
array[31697] <= 16'b0000_0000_0000_0000;
array[31698] <= 16'b0000_0000_0000_0000;
array[31699] <= 16'b0000_0000_0000_0000;
array[31700] <= 16'b0000_0000_0000_0000;
array[31701] <= 16'b0000_0000_0000_0000;
array[31702] <= 16'b0000_0000_0000_0000;
array[31703] <= 16'b0000_0000_0000_0000;
array[31704] <= 16'b0000_0000_0000_0000;
array[31705] <= 16'b0000_0000_0000_0000;
array[31706] <= 16'b0000_0000_0000_0000;
array[31707] <= 16'b0000_0000_0000_0000;
array[31708] <= 16'b0000_0000_0000_0000;
array[31709] <= 16'b0000_0000_0000_0000;
array[31710] <= 16'b0000_0000_0000_0000;
array[31711] <= 16'b0000_0000_0000_0000;
array[31712] <= 16'b0000_0000_0000_0000;
array[31713] <= 16'b0000_0000_0000_0000;
array[31714] <= 16'b0000_0000_0000_0000;
array[31715] <= 16'b0000_0000_0000_0000;
array[31716] <= 16'b0000_0000_0000_0000;
array[31717] <= 16'b0000_0000_0000_0000;
array[31718] <= 16'b0000_0000_0000_0000;
array[31719] <= 16'b0000_0000_0000_0000;
array[31720] <= 16'b0000_0000_0000_0000;
array[31721] <= 16'b0000_0000_0000_0000;
array[31722] <= 16'b0000_0000_0000_0000;
array[31723] <= 16'b0000_0000_0000_0000;
array[31724] <= 16'b0000_0000_0000_0000;
array[31725] <= 16'b0000_0000_0000_0000;
array[31726] <= 16'b0000_0000_0000_0000;
array[31727] <= 16'b0000_0000_0000_0000;
array[31728] <= 16'b0000_0000_0000_0000;
array[31729] <= 16'b0000_0000_0000_0000;
array[31730] <= 16'b0000_0000_0000_0000;
array[31731] <= 16'b0000_0000_0000_0000;
array[31732] <= 16'b0000_0000_0000_0000;
array[31733] <= 16'b0000_0000_0000_0000;
array[31734] <= 16'b0000_0000_0000_0000;
array[31735] <= 16'b0000_0000_0000_0000;
array[31736] <= 16'b0000_0000_0000_0000;
array[31737] <= 16'b0000_0000_0000_0000;
array[31738] <= 16'b0000_0000_0000_0000;
array[31739] <= 16'b0000_0000_0000_0000;
array[31740] <= 16'b0000_0000_0000_0000;
array[31741] <= 16'b0000_0000_0000_0000;
array[31742] <= 16'b0000_0000_0000_0000;
array[31743] <= 16'b0000_0000_0000_0000;
array[31744] <= 16'b0000_0000_0000_0000;
array[31745] <= 16'b0000_0000_0000_0000;
array[31746] <= 16'b0000_0000_0000_0000;
array[31747] <= 16'b0000_0000_0000_0000;
array[31748] <= 16'b0000_0000_0000_0000;
array[31749] <= 16'b0000_0000_0000_0000;
array[31750] <= 16'b0000_0000_0000_0000;
array[31751] <= 16'b0000_0000_0000_0000;
array[31752] <= 16'b0000_0000_0000_0000;
array[31753] <= 16'b0000_0000_0000_0000;
array[31754] <= 16'b0000_0000_0000_0000;
array[31755] <= 16'b0000_0000_0000_0000;
array[31756] <= 16'b0000_0000_0000_0000;
array[31757] <= 16'b0000_0000_0000_0000;
array[31758] <= 16'b0000_0000_0000_0000;
array[31759] <= 16'b0000_0000_0000_0000;
array[31760] <= 16'b0000_0000_0000_0000;
array[31761] <= 16'b0000_0000_0000_0000;
array[31762] <= 16'b0000_0000_0000_0000;
array[31763] <= 16'b0000_0000_0000_0000;
array[31764] <= 16'b0000_0000_0000_0000;
array[31765] <= 16'b0000_0000_0000_0000;
array[31766] <= 16'b0000_0000_0000_0000;
array[31767] <= 16'b0000_0000_0000_0000;
array[31768] <= 16'b0000_0000_0000_0000;
array[31769] <= 16'b0000_0000_0000_0000;
array[31770] <= 16'b0000_0000_0000_0000;
array[31771] <= 16'b0000_0000_0000_0000;
array[31772] <= 16'b0000_0000_0000_0000;
array[31773] <= 16'b0000_0000_0000_0000;
array[31774] <= 16'b0000_0000_0000_0000;
array[31775] <= 16'b0000_0000_0000_0000;
array[31776] <= 16'b0000_0000_0000_0000;
array[31777] <= 16'b0000_0000_0000_0000;
array[31778] <= 16'b0000_0000_0000_0000;
array[31779] <= 16'b0000_0000_0000_0000;
array[31780] <= 16'b0000_0000_0000_0000;
array[31781] <= 16'b0000_0000_0000_0000;
array[31782] <= 16'b0000_0000_0000_0000;
array[31783] <= 16'b0000_0000_0000_0000;
array[31784] <= 16'b0000_0000_0000_0000;
array[31785] <= 16'b0000_0000_0000_0000;
array[31786] <= 16'b0000_0000_0000_0000;
array[31787] <= 16'b0000_0000_0000_0000;
array[31788] <= 16'b0000_0000_0000_0000;
array[31789] <= 16'b0000_0000_0000_0000;
array[31790] <= 16'b0000_0000_0000_0000;
array[31791] <= 16'b0000_0000_0000_0000;
array[31792] <= 16'b0000_0000_0000_0000;
array[31793] <= 16'b0000_0000_0000_0000;
array[31794] <= 16'b0000_0000_0000_0000;
array[31795] <= 16'b0000_0000_0000_0000;
array[31796] <= 16'b0000_0000_0000_0000;
array[31797] <= 16'b0000_0000_0000_0000;
array[31798] <= 16'b0000_0000_0000_0000;
array[31799] <= 16'b0000_0000_0000_0000;
array[31800] <= 16'b0000_0000_0000_0000;
array[31801] <= 16'b0000_0000_0000_0000;
array[31802] <= 16'b0000_0000_0000_0000;
array[31803] <= 16'b0000_0000_0000_0000;
array[31804] <= 16'b0000_0000_0000_0000;
array[31805] <= 16'b0000_0000_0000_0000;
array[31806] <= 16'b0000_0000_0000_0000;
array[31807] <= 16'b0000_0000_0000_0000;
array[31808] <= 16'b0000_0000_0000_0000;
array[31809] <= 16'b0000_0000_0000_0000;
array[31810] <= 16'b0000_0000_0000_0000;
array[31811] <= 16'b0000_0000_0000_0000;
array[31812] <= 16'b0000_0000_0000_0000;
array[31813] <= 16'b0000_0000_0000_0000;
array[31814] <= 16'b0000_0000_0000_0000;
array[31815] <= 16'b0000_0000_0000_0000;
array[31816] <= 16'b0000_0000_0000_0000;
array[31817] <= 16'b0000_0000_0000_0000;
array[31818] <= 16'b0000_0000_0000_0000;
array[31819] <= 16'b0000_0000_0000_0000;
array[31820] <= 16'b0000_0000_0000_0000;
array[31821] <= 16'b0000_0000_0000_0000;
array[31822] <= 16'b0000_0000_0000_0000;
array[31823] <= 16'b0000_0000_0000_0000;
array[31824] <= 16'b0000_0000_0000_0000;
array[31825] <= 16'b0000_0000_0000_0000;
array[31826] <= 16'b0000_0000_0000_0000;
array[31827] <= 16'b0000_0000_0000_0000;
array[31828] <= 16'b0000_0000_0000_0000;
array[31829] <= 16'b0000_0000_0000_0000;
array[31830] <= 16'b0000_0000_0000_0000;
array[31831] <= 16'b0000_0000_0000_0000;
array[31832] <= 16'b0000_0000_0000_0000;
array[31833] <= 16'b0000_0000_0000_0000;
array[31834] <= 16'b0000_0000_0000_0000;
array[31835] <= 16'b0000_0000_0000_0000;
array[31836] <= 16'b0000_0000_0000_0000;
array[31837] <= 16'b0000_0000_0000_0000;
array[31838] <= 16'b0000_0000_0000_0000;
array[31839] <= 16'b0000_0000_0000_0000;
array[31840] <= 16'b0000_0000_0000_0000;
array[31841] <= 16'b0000_0000_0000_0000;
array[31842] <= 16'b0000_0000_0000_0000;
array[31843] <= 16'b0000_0000_0000_0000;
array[31844] <= 16'b0000_0000_0000_0000;
array[31845] <= 16'b0000_0000_0000_0000;
array[31846] <= 16'b0000_0000_0000_0000;
array[31847] <= 16'b0000_0000_0000_0000;
array[31848] <= 16'b0000_0000_0000_0000;
array[31849] <= 16'b0000_0000_0000_0000;
array[31850] <= 16'b0000_0000_0000_0000;
array[31851] <= 16'b0000_0000_0000_0000;
array[31852] <= 16'b0000_0000_0000_0000;
array[31853] <= 16'b0000_0000_0000_0000;
array[31854] <= 16'b0000_0000_0000_0000;
array[31855] <= 16'b0000_0000_0000_0000;
array[31856] <= 16'b0000_0000_0000_0000;
array[31857] <= 16'b0000_0000_0000_0000;
array[31858] <= 16'b0000_0000_0000_0000;
array[31859] <= 16'b0000_0000_0000_0000;
array[31860] <= 16'b0000_0000_0000_0000;
array[31861] <= 16'b0000_0000_0000_0000;
array[31862] <= 16'b0000_0000_0000_0000;
array[31863] <= 16'b0000_0000_0000_0000;
array[31864] <= 16'b0000_0000_0000_0000;
array[31865] <= 16'b0000_0000_0000_0000;
array[31866] <= 16'b0000_0000_0000_0000;
array[31867] <= 16'b0000_0000_0000_0000;
array[31868] <= 16'b0000_0000_0000_0000;
array[31869] <= 16'b0000_0000_0000_0000;
array[31870] <= 16'b0000_0000_0000_0000;
array[31871] <= 16'b0000_0000_0000_0000;
array[31872] <= 16'b0000_0000_0000_0000;
array[31873] <= 16'b0000_0000_0000_0000;
array[31874] <= 16'b0000_0000_0000_0000;
array[31875] <= 16'b0000_0000_0000_0000;
array[31876] <= 16'b0000_0000_0000_0000;
array[31877] <= 16'b0000_0000_0000_0000;
array[31878] <= 16'b0000_0000_0000_0000;
array[31879] <= 16'b0000_0000_0000_0000;
array[31880] <= 16'b0000_0000_0000_0000;
array[31881] <= 16'b0000_0000_0000_0000;
array[31882] <= 16'b0000_0000_0000_0000;
array[31883] <= 16'b0000_0000_0000_0000;
array[31884] <= 16'b0000_0000_0000_0000;
array[31885] <= 16'b0000_0000_0000_0000;
array[31886] <= 16'b0000_0000_0000_0000;
array[31887] <= 16'b0000_0000_0000_0000;
array[31888] <= 16'b0000_0000_0000_0000;
array[31889] <= 16'b0000_0000_0000_0000;
array[31890] <= 16'b0000_0000_0000_0000;
array[31891] <= 16'b0000_0000_0000_0000;
array[31892] <= 16'b0000_0000_0000_0000;
array[31893] <= 16'b0000_0000_0000_0000;
array[31894] <= 16'b0000_0000_0000_0000;
array[31895] <= 16'b0000_0000_0000_0000;
array[31896] <= 16'b0000_0000_0000_0000;
array[31897] <= 16'b0000_0000_0000_0000;
array[31898] <= 16'b0000_0000_0000_0000;
array[31899] <= 16'b0000_0000_0000_0000;
array[31900] <= 16'b0000_0000_0000_0000;
array[31901] <= 16'b0000_0000_0000_0000;
array[31902] <= 16'b0000_0000_0000_0000;
array[31903] <= 16'b0000_0000_0000_0000;
array[31904] <= 16'b0000_0000_0000_0000;
array[31905] <= 16'b0000_0000_0000_0000;
array[31906] <= 16'b0000_0000_0000_0000;
array[31907] <= 16'b0000_0000_0000_0000;
array[31908] <= 16'b0000_0000_0000_0000;
array[31909] <= 16'b0000_0000_0000_0000;
array[31910] <= 16'b0000_0000_0000_0000;
array[31911] <= 16'b0000_0000_0000_0000;
array[31912] <= 16'b0000_0000_0000_0000;
array[31913] <= 16'b0000_0000_0000_0000;
array[31914] <= 16'b0000_0000_0000_0000;
array[31915] <= 16'b0000_0000_0000_0000;
array[31916] <= 16'b0000_0000_0000_0000;
array[31917] <= 16'b0000_0000_0000_0000;
array[31918] <= 16'b0000_0000_0000_0000;
array[31919] <= 16'b0000_0000_0000_0000;
array[31920] <= 16'b0000_0000_0000_0000;
array[31921] <= 16'b0000_0000_0000_0000;
array[31922] <= 16'b0000_0000_0000_0000;
array[31923] <= 16'b0000_0000_0000_0000;
array[31924] <= 16'b0000_0000_0000_0000;
array[31925] <= 16'b0000_0000_0000_0000;
array[31926] <= 16'b0000_0000_0000_0000;
array[31927] <= 16'b0000_0000_0000_0000;
array[31928] <= 16'b0000_0000_0000_0000;
array[31929] <= 16'b0000_0000_0000_0000;
array[31930] <= 16'b0000_0000_0000_0000;
array[31931] <= 16'b0000_0000_0000_0000;
array[31932] <= 16'b0000_0000_0000_0000;
array[31933] <= 16'b0000_0000_0000_0000;
array[31934] <= 16'b0000_0000_0000_0000;
array[31935] <= 16'b0000_0000_0000_0000;
array[31936] <= 16'b0000_0000_0000_0000;
array[31937] <= 16'b0000_0000_0000_0000;
array[31938] <= 16'b0000_0000_0000_0000;
array[31939] <= 16'b0000_0000_0000_0000;
array[31940] <= 16'b0000_0000_0000_0000;
array[31941] <= 16'b0000_0000_0000_0000;
array[31942] <= 16'b0000_0000_0000_0000;
array[31943] <= 16'b0000_0000_0000_0000;
array[31944] <= 16'b0000_0000_0000_0000;
array[31945] <= 16'b0000_0000_0000_0000;
array[31946] <= 16'b0000_0000_0000_0000;
array[31947] <= 16'b0000_0000_0000_0000;
array[31948] <= 16'b0000_0000_0000_0000;
array[31949] <= 16'b0000_0000_0000_0000;
array[31950] <= 16'b0000_0000_0000_0000;
array[31951] <= 16'b0000_0000_0000_0000;
array[31952] <= 16'b0000_0000_0000_0000;
array[31953] <= 16'b0000_0000_0000_0000;
array[31954] <= 16'b0000_0000_0000_0000;
array[31955] <= 16'b0000_0000_0000_0000;
array[31956] <= 16'b0000_0000_0000_0000;
array[31957] <= 16'b0000_0000_0000_0000;
array[31958] <= 16'b0000_0000_0000_0000;
array[31959] <= 16'b0000_0000_0000_0000;
array[31960] <= 16'b0000_0000_0000_0000;
array[31961] <= 16'b0000_0000_0000_0000;
array[31962] <= 16'b0000_0000_0000_0000;
array[31963] <= 16'b0000_0000_0000_0000;
array[31964] <= 16'b0000_0000_0000_0000;
array[31965] <= 16'b0000_0000_0000_0000;
array[31966] <= 16'b0000_0000_0000_0000;
array[31967] <= 16'b0000_0000_0000_0000;
array[31968] <= 16'b0000_0000_0000_0000;
array[31969] <= 16'b0000_0000_0000_0000;
array[31970] <= 16'b0000_0000_0000_0000;
array[31971] <= 16'b0000_0000_0000_0000;
array[31972] <= 16'b0000_0000_0000_0000;
array[31973] <= 16'b0000_0000_0000_0000;
array[31974] <= 16'b0000_0000_0000_0000;
array[31975] <= 16'b0000_0000_0000_0000;
array[31976] <= 16'b0000_0000_0000_0000;
array[31977] <= 16'b0000_0000_0000_0000;
array[31978] <= 16'b0000_0000_0000_0000;
array[31979] <= 16'b0000_0000_0000_0000;
array[31980] <= 16'b0000_0000_0000_0000;
array[31981] <= 16'b0000_0000_0000_0000;
array[31982] <= 16'b0000_0000_0000_0000;
array[31983] <= 16'b0000_0000_0000_0000;
array[31984] <= 16'b0000_0000_0000_0000;
array[31985] <= 16'b0000_0000_0000_0000;
array[31986] <= 16'b0000_0000_0000_0000;
array[31987] <= 16'b0000_0000_0000_0000;
array[31988] <= 16'b0000_0000_0000_0000;
array[31989] <= 16'b0000_0000_0000_0000;
array[31990] <= 16'b0000_0000_0000_0000;
array[31991] <= 16'b0000_0000_0000_0000;
array[31992] <= 16'b0000_0000_0000_0000;
array[31993] <= 16'b0000_0000_0000_0000;
array[31994] <= 16'b0000_0000_0000_0000;
array[31995] <= 16'b0000_0000_0000_0000;
array[31996] <= 16'b0000_0000_0000_0000;
array[31997] <= 16'b0000_0000_0000_0000;
array[31998] <= 16'b0000_0000_0000_0000;
array[31999] <= 16'b0000_0000_0000_0000;
array[32000] <= 16'b0000_0000_0000_0000;
array[32001] <= 16'b0000_0000_0000_0000;
array[32002] <= 16'b0000_0000_0000_0000;
array[32003] <= 16'b0000_0000_0000_0000;
array[32004] <= 16'b0000_0000_0000_0000;
array[32005] <= 16'b0000_0000_0000_0000;
array[32006] <= 16'b0000_0000_0000_0000;
array[32007] <= 16'b0000_0000_0000_0000;
array[32008] <= 16'b0000_0000_0000_0000;
array[32009] <= 16'b0000_0000_0000_0000;
array[32010] <= 16'b0000_0000_0000_0000;
array[32011] <= 16'b0000_0000_0000_0000;
array[32012] <= 16'b0000_0000_0000_0000;
array[32013] <= 16'b0000_0000_0000_0000;
array[32014] <= 16'b0000_0000_0000_0000;
array[32015] <= 16'b0000_0000_0000_0000;
array[32016] <= 16'b0000_0000_0000_0000;
array[32017] <= 16'b0000_0000_0000_0000;
array[32018] <= 16'b0000_0000_0000_0000;
array[32019] <= 16'b0000_0000_0000_0000;
array[32020] <= 16'b0000_0000_0000_0000;
array[32021] <= 16'b0000_0000_0000_0000;
array[32022] <= 16'b0000_0000_0000_0000;
array[32023] <= 16'b0000_0000_0000_0000;
array[32024] <= 16'b0000_0000_0000_0000;
array[32025] <= 16'b0000_0000_0000_0000;
array[32026] <= 16'b0000_0000_0000_0000;
array[32027] <= 16'b0000_0000_0000_0000;
array[32028] <= 16'b0000_0000_0000_0000;
array[32029] <= 16'b0000_0000_0000_0000;
array[32030] <= 16'b0000_0000_0000_0000;
array[32031] <= 16'b0000_0000_0000_0000;
array[32032] <= 16'b0000_0000_0000_0000;
array[32033] <= 16'b0000_0000_0000_0000;
array[32034] <= 16'b0000_0000_0000_0000;
array[32035] <= 16'b0000_0000_0000_0000;
array[32036] <= 16'b0000_0000_0000_0000;
array[32037] <= 16'b0000_0000_0000_0000;
array[32038] <= 16'b0000_0000_0000_0000;
array[32039] <= 16'b0000_0000_0000_0000;
array[32040] <= 16'b0000_0000_0000_0000;
array[32041] <= 16'b0000_0000_0000_0000;
array[32042] <= 16'b0000_0000_0000_0000;
array[32043] <= 16'b0000_0000_0000_0000;
array[32044] <= 16'b0000_0000_0000_0000;
array[32045] <= 16'b0000_0000_0000_0000;
array[32046] <= 16'b0000_0000_0000_0000;
array[32047] <= 16'b0000_0000_0000_0000;
array[32048] <= 16'b0000_0000_0000_0000;
array[32049] <= 16'b0000_0000_0000_0000;
array[32050] <= 16'b0000_0000_0000_0000;
array[32051] <= 16'b0000_0000_0000_0000;
array[32052] <= 16'b0000_0000_0000_0000;
array[32053] <= 16'b0000_0000_0000_0000;
array[32054] <= 16'b0000_0000_0000_0000;
array[32055] <= 16'b0000_0000_0000_0000;
array[32056] <= 16'b0000_0000_0000_0000;
array[32057] <= 16'b0000_0000_0000_0000;
array[32058] <= 16'b0000_0000_0000_0000;
array[32059] <= 16'b0000_0000_0000_0000;
array[32060] <= 16'b0000_0000_0000_0000;
array[32061] <= 16'b0000_0000_0000_0000;
array[32062] <= 16'b0000_0000_0000_0000;
array[32063] <= 16'b0000_0000_0000_0000;
array[32064] <= 16'b0000_0000_0000_0000;
array[32065] <= 16'b0000_0000_0000_0000;
array[32066] <= 16'b0000_0000_0000_0000;
array[32067] <= 16'b0000_0000_0000_0000;
array[32068] <= 16'b0000_0000_0000_0000;
array[32069] <= 16'b0000_0000_0000_0000;
array[32070] <= 16'b0000_0000_0000_0000;
array[32071] <= 16'b0000_0000_0000_0000;
array[32072] <= 16'b0000_0000_0000_0000;
array[32073] <= 16'b0000_0000_0000_0000;
array[32074] <= 16'b0000_0000_0000_0000;
array[32075] <= 16'b0000_0000_0000_0000;
array[32076] <= 16'b0000_0000_0000_0000;
array[32077] <= 16'b0000_0000_0000_0000;
array[32078] <= 16'b0000_0000_0000_0000;
array[32079] <= 16'b0000_0000_0000_0000;
array[32080] <= 16'b0000_0000_0000_0000;
array[32081] <= 16'b0000_0000_0000_0000;
array[32082] <= 16'b0000_0000_0000_0000;
array[32083] <= 16'b0000_0000_0000_0000;
array[32084] <= 16'b0000_0000_0000_0000;
array[32085] <= 16'b0000_0000_0000_0000;
array[32086] <= 16'b0000_0000_0000_0000;
array[32087] <= 16'b0000_0000_0000_0000;
array[32088] <= 16'b0000_0000_0000_0000;
array[32089] <= 16'b0000_0000_0000_0000;
array[32090] <= 16'b0000_0000_0000_0000;
array[32091] <= 16'b0000_0000_0000_0000;
array[32092] <= 16'b0000_0000_0000_0000;
array[32093] <= 16'b0000_0000_0000_0000;
array[32094] <= 16'b0000_0000_0000_0000;
array[32095] <= 16'b0000_0000_0000_0000;
array[32096] <= 16'b0000_0000_0000_0000;
array[32097] <= 16'b0000_0000_0000_0000;
array[32098] <= 16'b0000_0000_0000_0000;
array[32099] <= 16'b0000_0000_0000_0000;
array[32100] <= 16'b0000_0000_0000_0000;
array[32101] <= 16'b0000_0000_0000_0000;
array[32102] <= 16'b0000_0000_0000_0000;
array[32103] <= 16'b0000_0000_0000_0000;
array[32104] <= 16'b0000_0000_0000_0000;
array[32105] <= 16'b0000_0000_0000_0000;
array[32106] <= 16'b0000_0000_0000_0000;
array[32107] <= 16'b0000_0000_0000_0000;
array[32108] <= 16'b0000_0000_0000_0000;
array[32109] <= 16'b0000_0000_0000_0000;
array[32110] <= 16'b0000_0000_0000_0000;
array[32111] <= 16'b0000_0000_0000_0000;
array[32112] <= 16'b0000_0000_0000_0000;
array[32113] <= 16'b0000_0000_0000_0000;
array[32114] <= 16'b0000_0000_0000_0000;
array[32115] <= 16'b0000_0000_0000_0000;
array[32116] <= 16'b0000_0000_0000_0000;
array[32117] <= 16'b0000_0000_0000_0000;
array[32118] <= 16'b0000_0000_0000_0000;
array[32119] <= 16'b0000_0000_0000_0000;
array[32120] <= 16'b0000_0000_0000_0000;
array[32121] <= 16'b0000_0000_0000_0000;
array[32122] <= 16'b0000_0000_0000_0000;
array[32123] <= 16'b0000_0000_0000_0000;
array[32124] <= 16'b0000_0000_0000_0000;
array[32125] <= 16'b0000_0000_0000_0000;
array[32126] <= 16'b0000_0000_0000_0000;
array[32127] <= 16'b0000_0000_0000_0000;
array[32128] <= 16'b0000_0000_0000_0000;
array[32129] <= 16'b0000_0000_0000_0000;
array[32130] <= 16'b0000_0000_0000_0000;
array[32131] <= 16'b0000_0000_0000_0000;
array[32132] <= 16'b0000_0000_0000_0000;
array[32133] <= 16'b0000_0000_0000_0000;
array[32134] <= 16'b0000_0000_0000_0000;
array[32135] <= 16'b0000_0000_0000_0000;
array[32136] <= 16'b0000_0000_0000_0000;
array[32137] <= 16'b0000_0000_0000_0000;
array[32138] <= 16'b0000_0000_0000_0000;
array[32139] <= 16'b0000_0000_0000_0000;
array[32140] <= 16'b0000_0000_0000_0000;
array[32141] <= 16'b0000_0000_0000_0000;
array[32142] <= 16'b0000_0000_0000_0000;
array[32143] <= 16'b0000_0000_0000_0000;
array[32144] <= 16'b0000_0000_0000_0000;
array[32145] <= 16'b0000_0000_0000_0000;
array[32146] <= 16'b0000_0000_0000_0000;
array[32147] <= 16'b0000_0000_0000_0000;
array[32148] <= 16'b0000_0000_0000_0000;
array[32149] <= 16'b0000_0000_0000_0000;
array[32150] <= 16'b0000_0000_0000_0000;
array[32151] <= 16'b0000_0000_0000_0000;
array[32152] <= 16'b0000_0000_0000_0000;
array[32153] <= 16'b0000_0000_0000_0000;
array[32154] <= 16'b0000_0000_0000_0000;
array[32155] <= 16'b0000_0000_0000_0000;
array[32156] <= 16'b0000_0000_0000_0000;
array[32157] <= 16'b0000_0000_0000_0000;
array[32158] <= 16'b0000_0000_0000_0000;
array[32159] <= 16'b0000_0000_0000_0000;
array[32160] <= 16'b0000_0000_0000_0000;
array[32161] <= 16'b0000_0000_0000_0000;
array[32162] <= 16'b0000_0000_0000_0000;
array[32163] <= 16'b0000_0000_0000_0000;
array[32164] <= 16'b0000_0000_0000_0000;
array[32165] <= 16'b0000_0000_0000_0000;
array[32166] <= 16'b0000_0000_0000_0000;
array[32167] <= 16'b0000_0000_0000_0000;
array[32168] <= 16'b0000_0000_0000_0000;
array[32169] <= 16'b0000_0000_0000_0000;
array[32170] <= 16'b0000_0000_0000_0000;
array[32171] <= 16'b0000_0000_0000_0000;
array[32172] <= 16'b0000_0000_0000_0000;
array[32173] <= 16'b0000_0000_0000_0000;
array[32174] <= 16'b0000_0000_0000_0000;
array[32175] <= 16'b0000_0000_0000_0000;
array[32176] <= 16'b0000_0000_0000_0000;
array[32177] <= 16'b0000_0000_0000_0000;
array[32178] <= 16'b0000_0000_0000_0000;
array[32179] <= 16'b0000_0000_0000_0000;
array[32180] <= 16'b0000_0000_0000_0000;
array[32181] <= 16'b0000_0000_0000_0000;
array[32182] <= 16'b0000_0000_0000_0000;
array[32183] <= 16'b0000_0000_0000_0000;
array[32184] <= 16'b0000_0000_0000_0000;
array[32185] <= 16'b0000_0000_0000_0000;
array[32186] <= 16'b0000_0000_0000_0000;
array[32187] <= 16'b0000_0000_0000_0000;
array[32188] <= 16'b0000_0000_0000_0000;
array[32189] <= 16'b0000_0000_0000_0000;
array[32190] <= 16'b0000_0000_0000_0000;
array[32191] <= 16'b0000_0000_0000_0000;
array[32192] <= 16'b0000_0000_0000_0000;
array[32193] <= 16'b0000_0000_0000_0000;
array[32194] <= 16'b0000_0000_0000_0000;
array[32195] <= 16'b0000_0000_0000_0000;
array[32196] <= 16'b0000_0000_0000_0000;
array[32197] <= 16'b0000_0000_0000_0000;
array[32198] <= 16'b0000_0000_0000_0000;
array[32199] <= 16'b0000_0000_0000_0000;
array[32200] <= 16'b0000_0000_0000_0000;
array[32201] <= 16'b0000_0000_0000_0000;
array[32202] <= 16'b0000_0000_0000_0000;
array[32203] <= 16'b0000_0000_0000_0000;
array[32204] <= 16'b0000_0000_0000_0000;
array[32205] <= 16'b0000_0000_0000_0000;
array[32206] <= 16'b0000_0000_0000_0000;
array[32207] <= 16'b0000_0000_0000_0000;
array[32208] <= 16'b0000_0000_0000_0000;
array[32209] <= 16'b0000_0000_0000_0000;
array[32210] <= 16'b0000_0000_0000_0000;
array[32211] <= 16'b0000_0000_0000_0000;
array[32212] <= 16'b0000_0000_0000_0000;
array[32213] <= 16'b0000_0000_0000_0000;
array[32214] <= 16'b0000_0000_0000_0000;
array[32215] <= 16'b0000_0000_0000_0000;
array[32216] <= 16'b0000_0000_0000_0000;
array[32217] <= 16'b0000_0000_0000_0000;
array[32218] <= 16'b0000_0000_0000_0000;
array[32219] <= 16'b0000_0000_0000_0000;
array[32220] <= 16'b0000_0000_0000_0000;
array[32221] <= 16'b0000_0000_0000_0000;
array[32222] <= 16'b0000_0000_0000_0000;
array[32223] <= 16'b0000_0000_0000_0000;
array[32224] <= 16'b0000_0000_0000_0000;
array[32225] <= 16'b0000_0000_0000_0000;
array[32226] <= 16'b0000_0000_0000_0000;
array[32227] <= 16'b0000_0000_0000_0000;
array[32228] <= 16'b0000_0000_0000_0000;
array[32229] <= 16'b0000_0000_0000_0000;
array[32230] <= 16'b0000_0000_0000_0000;
array[32231] <= 16'b0000_0000_0000_0000;
array[32232] <= 16'b0000_0000_0000_0000;
array[32233] <= 16'b0000_0000_0000_0000;
array[32234] <= 16'b0000_0000_0000_0000;
array[32235] <= 16'b0000_0000_0000_0000;
array[32236] <= 16'b0000_0000_0000_0000;
array[32237] <= 16'b0000_0000_0000_0000;
array[32238] <= 16'b0000_0000_0000_0000;
array[32239] <= 16'b0000_0000_0000_0000;
array[32240] <= 16'b0000_0000_0000_0000;
array[32241] <= 16'b0000_0000_0000_0000;
array[32242] <= 16'b0000_0000_0000_0000;
array[32243] <= 16'b0000_0000_0000_0000;
array[32244] <= 16'b0000_0000_0000_0000;
array[32245] <= 16'b0000_0000_0000_0000;
array[32246] <= 16'b0000_0000_0000_0000;
array[32247] <= 16'b0000_0000_0000_0000;
array[32248] <= 16'b0000_0000_0000_0000;
array[32249] <= 16'b0000_0000_0000_0000;
array[32250] <= 16'b0000_0000_0000_0000;
array[32251] <= 16'b0000_0000_0000_0000;
array[32252] <= 16'b0000_0000_0000_0000;
array[32253] <= 16'b0000_0000_0000_0000;
array[32254] <= 16'b0000_0000_0000_0000;
array[32255] <= 16'b0000_0000_0000_0000;
array[32256] <= 16'b0000_0000_0000_0000;
array[32257] <= 16'b0000_0000_0000_0000;
array[32258] <= 16'b0000_0000_0000_0000;
array[32259] <= 16'b0000_0000_0000_0000;
array[32260] <= 16'b0000_0000_0000_0000;
array[32261] <= 16'b0000_0000_0000_0000;
array[32262] <= 16'b0000_0000_0000_0000;
array[32263] <= 16'b0000_0000_0000_0000;
array[32264] <= 16'b0000_0000_0000_0000;
array[32265] <= 16'b0000_0000_0000_0000;
array[32266] <= 16'b0000_0000_0000_0000;
array[32267] <= 16'b0000_0000_0000_0000;
array[32268] <= 16'b0000_0000_0000_0000;
array[32269] <= 16'b0000_0000_0000_0000;
array[32270] <= 16'b0000_0000_0000_0000;
array[32271] <= 16'b0000_0000_0000_0000;
array[32272] <= 16'b0000_0000_0000_0000;
array[32273] <= 16'b0000_0000_0000_0000;
array[32274] <= 16'b0000_0000_0000_0000;
array[32275] <= 16'b0000_0000_0000_0000;
array[32276] <= 16'b0000_0000_0000_0000;
array[32277] <= 16'b0000_0000_0000_0000;
array[32278] <= 16'b0000_0000_0000_0000;
array[32279] <= 16'b0000_0000_0000_0000;
array[32280] <= 16'b0000_0000_0000_0000;
array[32281] <= 16'b0000_0000_0000_0000;
array[32282] <= 16'b0000_0000_0000_0000;
array[32283] <= 16'b0000_0000_0000_0000;
array[32284] <= 16'b0000_0000_0000_0000;
array[32285] <= 16'b0000_0000_0000_0000;
array[32286] <= 16'b0000_0000_0000_0000;
array[32287] <= 16'b0000_0000_0000_0000;
array[32288] <= 16'b0000_0000_0000_0000;
array[32289] <= 16'b0000_0000_0000_0000;
array[32290] <= 16'b0000_0000_0000_0000;
array[32291] <= 16'b0000_0000_0000_0000;
array[32292] <= 16'b0000_0000_0000_0000;
array[32293] <= 16'b0000_0000_0000_0000;
array[32294] <= 16'b0000_0000_0000_0000;
array[32295] <= 16'b0000_0000_0000_0000;
array[32296] <= 16'b0000_0000_0000_0000;
array[32297] <= 16'b0000_0000_0000_0000;
array[32298] <= 16'b0000_0000_0000_0000;
array[32299] <= 16'b0000_0000_0000_0000;
array[32300] <= 16'b0000_0000_0000_0000;
array[32301] <= 16'b0000_0000_0000_0000;
array[32302] <= 16'b0000_0000_0000_0000;
array[32303] <= 16'b0000_0000_0000_0000;
array[32304] <= 16'b0000_0000_0000_0000;
array[32305] <= 16'b0000_0000_0000_0000;
array[32306] <= 16'b0000_0000_0000_0000;
array[32307] <= 16'b0000_0000_0000_0000;
array[32308] <= 16'b0000_0000_0000_0000;
array[32309] <= 16'b0000_0000_0000_0000;
array[32310] <= 16'b0000_0000_0000_0000;
array[32311] <= 16'b0000_0000_0000_0000;
array[32312] <= 16'b0000_0000_0000_0000;
array[32313] <= 16'b0000_0000_0000_0000;
array[32314] <= 16'b0000_0000_0000_0000;
array[32315] <= 16'b0000_0000_0000_0000;
array[32316] <= 16'b0000_0000_0000_0000;
array[32317] <= 16'b0000_0000_0000_0000;
array[32318] <= 16'b0000_0000_0000_0000;
array[32319] <= 16'b0000_0000_0000_0000;
array[32320] <= 16'b0000_0000_0000_0000;
array[32321] <= 16'b0000_0000_0000_0000;
array[32322] <= 16'b0000_0000_0000_0000;
array[32323] <= 16'b0000_0000_0000_0000;
array[32324] <= 16'b0000_0000_0000_0000;
array[32325] <= 16'b0000_0000_0000_0000;
array[32326] <= 16'b0000_0000_0000_0000;
array[32327] <= 16'b0000_0000_0000_0000;
array[32328] <= 16'b0000_0000_0000_0000;
array[32329] <= 16'b0000_0000_0000_0000;
array[32330] <= 16'b0000_0000_0000_0000;
array[32331] <= 16'b0000_0000_0000_0000;
array[32332] <= 16'b0000_0000_0000_0000;
array[32333] <= 16'b0000_0000_0000_0000;
array[32334] <= 16'b0000_0000_0000_0000;
array[32335] <= 16'b0000_0000_0000_0000;
array[32336] <= 16'b0000_0000_0000_0000;
array[32337] <= 16'b0000_0000_0000_0000;
array[32338] <= 16'b0000_0000_0000_0000;
array[32339] <= 16'b0000_0000_0000_0000;
array[32340] <= 16'b0000_0000_0000_0000;
array[32341] <= 16'b0000_0000_0000_0000;
array[32342] <= 16'b0000_0000_0000_0000;
array[32343] <= 16'b0000_0000_0000_0000;
array[32344] <= 16'b0000_0000_0000_0000;
array[32345] <= 16'b0000_0000_0000_0000;
array[32346] <= 16'b0000_0000_0000_0000;
array[32347] <= 16'b0000_0000_0000_0000;
array[32348] <= 16'b0000_0000_0000_0000;
array[32349] <= 16'b0000_0000_0000_0000;
array[32350] <= 16'b0000_0000_0000_0000;
array[32351] <= 16'b0000_0000_0000_0000;
array[32352] <= 16'b0000_0000_0000_0000;
array[32353] <= 16'b0000_0000_0000_0000;
array[32354] <= 16'b0000_0000_0000_0000;
array[32355] <= 16'b0000_0000_0000_0000;
array[32356] <= 16'b0000_0000_0000_0000;
array[32357] <= 16'b0000_0000_0000_0000;
array[32358] <= 16'b0000_0000_0000_0000;
array[32359] <= 16'b0000_0000_0000_0000;
array[32360] <= 16'b0000_0000_0000_0000;
array[32361] <= 16'b0000_0000_0000_0000;
array[32362] <= 16'b0000_0000_0000_0000;
array[32363] <= 16'b0000_0000_0000_0000;
array[32364] <= 16'b0000_0000_0000_0000;
array[32365] <= 16'b0000_0000_0000_0000;
array[32366] <= 16'b0000_0000_0000_0000;
array[32367] <= 16'b0000_0000_0000_0000;
array[32368] <= 16'b0000_0000_0000_0000;
array[32369] <= 16'b0000_0000_0000_0000;
array[32370] <= 16'b0000_0000_0000_0000;
array[32371] <= 16'b0000_0000_0000_0000;
array[32372] <= 16'b0000_0000_0000_0000;
array[32373] <= 16'b0000_0000_0000_0000;
array[32374] <= 16'b0000_0000_0000_0000;
array[32375] <= 16'b0000_0000_0000_0000;
array[32376] <= 16'b0000_0000_0000_0000;
array[32377] <= 16'b0000_0000_0000_0000;
array[32378] <= 16'b0000_0000_0000_0000;
array[32379] <= 16'b0000_0000_0000_0000;
array[32380] <= 16'b0000_0000_0000_0000;
array[32381] <= 16'b0000_0000_0000_0000;
array[32382] <= 16'b0000_0000_0000_0000;
array[32383] <= 16'b0000_0000_0000_0000;
array[32384] <= 16'b0000_0000_0000_0000;
array[32385] <= 16'b0000_0000_0000_0000;
array[32386] <= 16'b0000_0000_0000_0000;
array[32387] <= 16'b0000_0000_0000_0000;
array[32388] <= 16'b0000_0000_0000_0000;
array[32389] <= 16'b0000_0000_0000_0000;
array[32390] <= 16'b0000_0000_0000_0000;
array[32391] <= 16'b0000_0000_0000_0000;
array[32392] <= 16'b0000_0000_0000_0000;
array[32393] <= 16'b0000_0000_0000_0000;
array[32394] <= 16'b0000_0000_0000_0000;
array[32395] <= 16'b0000_0000_0000_0000;
array[32396] <= 16'b0000_0000_0000_0000;
array[32397] <= 16'b0000_0000_0000_0000;
array[32398] <= 16'b0000_0000_0000_0000;
array[32399] <= 16'b0000_0000_0000_0000;
array[32400] <= 16'b0000_0000_0000_0000;
array[32401] <= 16'b0000_0000_0000_0000;
array[32402] <= 16'b0000_0000_0000_0000;
array[32403] <= 16'b0000_0000_0000_0000;
array[32404] <= 16'b0000_0000_0000_0000;
array[32405] <= 16'b0000_0000_0000_0000;
array[32406] <= 16'b0000_0000_0000_0000;
array[32407] <= 16'b0000_0000_0000_0000;
array[32408] <= 16'b0000_0000_0000_0000;
array[32409] <= 16'b0000_0000_0000_0000;
array[32410] <= 16'b0000_0000_0000_0000;
array[32411] <= 16'b0000_0000_0000_0000;
array[32412] <= 16'b0000_0000_0000_0000;
array[32413] <= 16'b0000_0000_0000_0000;
array[32414] <= 16'b0000_0000_0000_0000;
array[32415] <= 16'b0000_0000_0000_0000;
array[32416] <= 16'b0000_0000_0000_0000;
array[32417] <= 16'b0000_0000_0000_0000;
array[32418] <= 16'b0000_0000_0000_0000;
array[32419] <= 16'b0000_0000_0000_0000;
array[32420] <= 16'b0000_0000_0000_0000;
array[32421] <= 16'b0000_0000_0000_0000;
array[32422] <= 16'b0000_0000_0000_0000;
array[32423] <= 16'b0000_0000_0000_0000;
array[32424] <= 16'b0000_0000_0000_0000;
array[32425] <= 16'b0000_0000_0000_0000;
array[32426] <= 16'b0000_0000_0000_0000;
array[32427] <= 16'b0000_0000_0000_0000;
array[32428] <= 16'b0000_0000_0000_0000;
array[32429] <= 16'b0000_0000_0000_0000;
array[32430] <= 16'b0000_0000_0000_0000;
array[32431] <= 16'b0000_0000_0000_0000;
array[32432] <= 16'b0000_0000_0000_0000;
array[32433] <= 16'b0000_0000_0000_0000;
array[32434] <= 16'b0000_0000_0000_0000;
array[32435] <= 16'b0000_0000_0000_0000;
array[32436] <= 16'b0000_0000_0000_0000;
array[32437] <= 16'b0000_0000_0000_0000;
array[32438] <= 16'b0000_0000_0000_0000;
array[32439] <= 16'b0000_0000_0000_0000;
array[32440] <= 16'b0000_0000_0000_0000;
array[32441] <= 16'b0000_0000_0000_0000;
array[32442] <= 16'b0000_0000_0000_0000;
array[32443] <= 16'b0000_0000_0000_0000;
array[32444] <= 16'b0000_0000_0000_0000;
array[32445] <= 16'b0000_0000_0000_0000;
array[32446] <= 16'b0000_0000_0000_0000;
array[32447] <= 16'b0000_0000_0000_0000;
array[32448] <= 16'b0000_0000_0000_0000;
array[32449] <= 16'b0000_0000_0000_0000;
array[32450] <= 16'b0000_0000_0000_0000;
array[32451] <= 16'b0000_0000_0000_0000;
array[32452] <= 16'b0000_0000_0000_0000;
array[32453] <= 16'b0000_0000_0000_0000;
array[32454] <= 16'b0000_0000_0000_0000;
array[32455] <= 16'b0000_0000_0000_0000;
array[32456] <= 16'b0000_0000_0000_0000;
array[32457] <= 16'b0000_0000_0000_0000;
array[32458] <= 16'b0000_0000_0000_0000;
array[32459] <= 16'b0000_0000_0000_0000;
array[32460] <= 16'b0000_0000_0000_0000;
array[32461] <= 16'b0000_0000_0000_0000;
array[32462] <= 16'b0000_0000_0000_0000;
array[32463] <= 16'b0000_0000_0000_0000;
array[32464] <= 16'b0000_0000_0000_0000;
array[32465] <= 16'b0000_0000_0000_0000;
array[32466] <= 16'b0000_0000_0000_0000;
array[32467] <= 16'b0000_0000_0000_0000;
array[32468] <= 16'b0000_0000_0000_0000;
array[32469] <= 16'b0000_0000_0000_0000;
array[32470] <= 16'b0000_0000_0000_0000;
array[32471] <= 16'b0000_0000_0000_0000;
array[32472] <= 16'b0000_0000_0000_0000;
array[32473] <= 16'b0000_0000_0000_0000;
array[32474] <= 16'b0000_0000_0000_0000;
array[32475] <= 16'b0000_0000_0000_0000;
array[32476] <= 16'b0000_0000_0000_0000;
array[32477] <= 16'b0000_0000_0000_0000;
array[32478] <= 16'b0000_0000_0000_0000;
array[32479] <= 16'b0000_0000_0000_0000;
array[32480] <= 16'b0000_0000_0000_0000;
array[32481] <= 16'b0000_0000_0000_0000;
array[32482] <= 16'b0000_0000_0000_0000;
array[32483] <= 16'b0000_0000_0000_0000;
array[32484] <= 16'b0000_0000_0000_0000;
array[32485] <= 16'b0000_0000_0000_0000;
array[32486] <= 16'b0000_0000_0000_0000;
array[32487] <= 16'b0000_0000_0000_0000;
array[32488] <= 16'b0000_0000_0000_0000;
array[32489] <= 16'b0000_0000_0000_0000;
array[32490] <= 16'b0000_0000_0000_0000;
array[32491] <= 16'b0000_0000_0000_0000;
array[32492] <= 16'b0000_0000_0000_0000;
array[32493] <= 16'b0000_0000_0000_0000;
array[32494] <= 16'b0000_0000_0000_0000;
array[32495] <= 16'b0000_0000_0000_0000;
array[32496] <= 16'b0000_0000_0000_0000;
array[32497] <= 16'b0000_0000_0000_0000;
array[32498] <= 16'b0000_0000_0000_0000;
array[32499] <= 16'b0000_0000_0000_0000;
array[32500] <= 16'b0000_0000_0000_0000;
array[32501] <= 16'b0000_0000_0000_0000;
array[32502] <= 16'b0000_0000_0000_0000;
array[32503] <= 16'b0000_0000_0000_0000;
array[32504] <= 16'b0000_0000_0000_0000;
array[32505] <= 16'b0000_0000_0000_0000;
array[32506] <= 16'b0000_0000_0000_0000;
array[32507] <= 16'b0000_0000_0000_0000;
array[32508] <= 16'b0000_0000_0000_0000;
array[32509] <= 16'b0000_0000_0000_0000;
array[32510] <= 16'b0000_0000_0000_0000;
array[32511] <= 16'b0000_0000_0000_0000;
array[32512] <= 16'b0000_0000_0000_0000;
array[32513] <= 16'b0000_0000_0000_0000;
array[32514] <= 16'b0000_0000_0000_0000;
array[32515] <= 16'b0000_0000_0000_0000;
array[32516] <= 16'b0000_0000_0000_0000;
array[32517] <= 16'b0000_0000_0000_0000;
array[32518] <= 16'b0000_0000_0000_0000;
array[32519] <= 16'b0000_0000_0000_0000;
array[32520] <= 16'b0000_0000_0000_0000;
array[32521] <= 16'b0000_0000_0000_0000;
array[32522] <= 16'b0000_0000_0000_0000;
array[32523] <= 16'b0000_0000_0000_0000;
array[32524] <= 16'b0000_0000_0000_0000;
array[32525] <= 16'b0000_0000_0000_0000;
array[32526] <= 16'b0000_0000_0000_0000;
array[32527] <= 16'b0000_0000_0000_0000;
array[32528] <= 16'b0000_0000_0000_0000;
array[32529] <= 16'b0000_0000_0000_0000;
array[32530] <= 16'b0000_0000_0000_0000;
array[32531] <= 16'b0000_0000_0000_0000;
array[32532] <= 16'b0000_0000_0000_0000;
array[32533] <= 16'b0000_0000_0000_0000;
array[32534] <= 16'b0000_0000_0000_0000;
array[32535] <= 16'b0000_0000_0000_0000;
array[32536] <= 16'b0000_0000_0000_0000;
array[32537] <= 16'b0000_0000_0000_0000;
array[32538] <= 16'b0000_0000_0000_0000;
array[32539] <= 16'b0000_0000_0000_0000;
array[32540] <= 16'b0000_0000_0000_0000;
array[32541] <= 16'b0000_0000_0000_0000;
array[32542] <= 16'b0000_0000_0000_0000;
array[32543] <= 16'b0000_0000_0000_0000;
array[32544] <= 16'b0000_0000_0000_0000;
array[32545] <= 16'b0000_0000_0000_0000;
array[32546] <= 16'b0000_0000_0000_0000;
array[32547] <= 16'b0000_0000_0000_0000;
array[32548] <= 16'b0000_0000_0000_0000;
array[32549] <= 16'b0000_0000_0000_0000;
array[32550] <= 16'b0000_0000_0000_0000;
array[32551] <= 16'b0000_0000_0000_0000;
array[32552] <= 16'b0000_0000_0000_0000;
array[32553] <= 16'b0000_0000_0000_0000;
array[32554] <= 16'b0000_0000_0000_0000;
array[32555] <= 16'b0000_0000_0000_0000;
array[32556] <= 16'b0000_0000_0000_0000;
array[32557] <= 16'b0000_0000_0000_0000;
array[32558] <= 16'b0000_0000_0000_0000;
array[32559] <= 16'b0000_0000_0000_0000;
array[32560] <= 16'b0000_0000_0000_0000;
array[32561] <= 16'b0000_0000_0000_0000;
array[32562] <= 16'b0000_0000_0000_0000;
array[32563] <= 16'b0000_0000_0000_0000;
array[32564] <= 16'b0000_0000_0000_0000;
array[32565] <= 16'b0000_0000_0000_0000;
array[32566] <= 16'b0000_0000_0000_0000;
array[32567] <= 16'b0000_0000_0000_0000;
array[32568] <= 16'b0000_0000_0000_0000;
array[32569] <= 16'b0000_0000_0000_0000;
array[32570] <= 16'b0000_0000_0000_0000;
array[32571] <= 16'b0000_0000_0000_0000;
array[32572] <= 16'b0000_0000_0000_0000;
array[32573] <= 16'b0000_0000_0000_0000;
array[32574] <= 16'b0000_0000_0000_0000;
array[32575] <= 16'b0000_0000_0000_0000;
array[32576] <= 16'b0000_0000_0000_0000;
array[32577] <= 16'b0000_0000_0000_0000;
array[32578] <= 16'b0000_0000_0000_0000;
array[32579] <= 16'b0000_0000_0000_0000;
array[32580] <= 16'b0000_0000_0000_0000;
array[32581] <= 16'b0000_0000_0000_0000;
array[32582] <= 16'b0000_0000_0000_0000;
array[32583] <= 16'b0000_0000_0000_0000;
array[32584] <= 16'b0000_0000_0000_0000;
array[32585] <= 16'b0000_0000_0000_0000;
array[32586] <= 16'b0000_0000_0000_0000;
array[32587] <= 16'b0000_0000_0000_0000;
array[32588] <= 16'b0000_0000_0000_0000;
array[32589] <= 16'b0000_0000_0000_0000;
array[32590] <= 16'b0000_0000_0000_0000;
array[32591] <= 16'b0000_0000_0000_0000;
array[32592] <= 16'b0000_0000_0000_0000;
array[32593] <= 16'b0000_0000_0000_0000;
array[32594] <= 16'b0000_0000_0000_0000;
array[32595] <= 16'b0000_0000_0000_0000;
array[32596] <= 16'b0000_0000_0000_0000;
array[32597] <= 16'b0000_0000_0000_0000;
array[32598] <= 16'b0000_0000_0000_0000;
array[32599] <= 16'b0000_0000_0000_0000;
array[32600] <= 16'b0000_0000_0000_0000;
array[32601] <= 16'b0000_0000_0000_0000;
array[32602] <= 16'b0000_0000_0000_0000;
array[32603] <= 16'b0000_0000_0000_0000;
array[32604] <= 16'b0000_0000_0000_0000;
array[32605] <= 16'b0000_0000_0000_0000;
array[32606] <= 16'b0000_0000_0000_0000;
array[32607] <= 16'b0000_0000_0000_0000;
array[32608] <= 16'b0000_0000_0000_0000;
array[32609] <= 16'b0000_0000_0000_0000;
array[32610] <= 16'b0000_0000_0000_0000;
array[32611] <= 16'b0000_0000_0000_0000;
array[32612] <= 16'b0000_0000_0000_0000;
array[32613] <= 16'b0000_0000_0000_0000;
array[32614] <= 16'b0000_0000_0000_0000;
array[32615] <= 16'b0000_0000_0000_0000;
array[32616] <= 16'b0000_0000_0000_0000;
array[32617] <= 16'b0000_0000_0000_0000;
array[32618] <= 16'b0000_0000_0000_0000;
array[32619] <= 16'b0000_0000_0000_0000;
array[32620] <= 16'b0000_0000_0000_0000;
array[32621] <= 16'b0000_0000_0000_0000;
array[32622] <= 16'b0000_0000_0000_0000;
array[32623] <= 16'b0000_0000_0000_0000;
array[32624] <= 16'b0000_0000_0000_0000;
array[32625] <= 16'b0000_0000_0000_0000;
array[32626] <= 16'b0000_0000_0000_0000;
array[32627] <= 16'b0000_0000_0000_0000;
array[32628] <= 16'b0000_0000_0000_0000;
array[32629] <= 16'b0000_0000_0000_0000;
array[32630] <= 16'b0000_0000_0000_0000;
array[32631] <= 16'b0000_0000_0000_0000;
array[32632] <= 16'b0000_0000_0000_0000;
array[32633] <= 16'b0000_0000_0000_0000;
array[32634] <= 16'b0000_0000_0000_0000;
array[32635] <= 16'b0000_0000_0000_0000;
array[32636] <= 16'b0000_0000_0000_0000;
array[32637] <= 16'b0000_0000_0000_0000;
array[32638] <= 16'b0000_0000_0000_0000;
array[32639] <= 16'b0000_0000_0000_0000;
array[32640] <= 16'b0000_0000_0000_0000;
array[32641] <= 16'b0000_0000_0000_0000;
array[32642] <= 16'b0000_0000_0000_0000;
array[32643] <= 16'b0000_0000_0000_0000;
array[32644] <= 16'b0000_0000_0000_0000;
array[32645] <= 16'b0000_0000_0000_0000;
array[32646] <= 16'b0000_0000_0000_0000;
array[32647] <= 16'b0000_0000_0000_0000;
array[32648] <= 16'b0000_0000_0000_0000;
array[32649] <= 16'b0000_0000_0000_0000;
array[32650] <= 16'b0000_0000_0000_0000;
array[32651] <= 16'b0000_0000_0000_0000;
array[32652] <= 16'b0000_0000_0000_0000;
array[32653] <= 16'b0000_0000_0000_0000;
array[32654] <= 16'b0000_0000_0000_0000;
array[32655] <= 16'b0000_0000_0000_0000;
array[32656] <= 16'b0000_0000_0000_0000;
array[32657] <= 16'b0000_0000_0000_0000;
array[32658] <= 16'b0000_0000_0000_0000;
array[32659] <= 16'b0000_0000_0000_0000;
array[32660] <= 16'b0000_0000_0000_0000;
array[32661] <= 16'b0000_0000_0000_0000;
array[32662] <= 16'b0000_0000_0000_0000;
array[32663] <= 16'b0000_0000_0000_0000;
array[32664] <= 16'b0000_0000_0000_0000;
array[32665] <= 16'b0000_0000_0000_0000;
array[32666] <= 16'b0000_0000_0000_0000;
array[32667] <= 16'b0000_0000_0000_0000;
array[32668] <= 16'b0000_0000_0000_0000;
array[32669] <= 16'b0000_0000_0000_0000;
array[32670] <= 16'b0000_0000_0000_0000;
array[32671] <= 16'b0000_0000_0000_0000;
array[32672] <= 16'b0000_0000_0000_0000;
array[32673] <= 16'b0000_0000_0000_0000;
array[32674] <= 16'b0000_0000_0000_0000;
array[32675] <= 16'b0000_0000_0000_0000;
array[32676] <= 16'b0000_0000_0000_0000;
array[32677] <= 16'b0000_0000_0000_0000;
array[32678] <= 16'b0000_0000_0000_0000;
array[32679] <= 16'b0000_0000_0000_0000;
array[32680] <= 16'b0000_0000_0000_0000;
array[32681] <= 16'b0000_0000_0000_0000;
array[32682] <= 16'b0000_0000_0000_0000;
array[32683] <= 16'b0000_0000_0000_0000;
array[32684] <= 16'b0000_0000_0000_0000;
array[32685] <= 16'b0000_0000_0000_0000;
array[32686] <= 16'b0000_0000_0000_0000;
array[32687] <= 16'b0000_0000_0000_0000;
array[32688] <= 16'b0000_0000_0000_0000;
array[32689] <= 16'b0000_0000_0000_0000;
array[32690] <= 16'b0000_0000_0000_0000;
array[32691] <= 16'b0000_0000_0000_0000;
array[32692] <= 16'b0000_0000_0000_0000;
array[32693] <= 16'b0000_0000_0000_0000;
array[32694] <= 16'b0000_0000_0000_0000;
array[32695] <= 16'b0000_0000_0000_0000;
array[32696] <= 16'b0000_0000_0000_0000;
array[32697] <= 16'b0000_0000_0000_0000;
array[32698] <= 16'b0000_0000_0000_0000;
array[32699] <= 16'b0000_0000_0000_0000;
array[32700] <= 16'b0000_0000_0000_0000;
array[32701] <= 16'b0000_0000_0000_0000;
array[32702] <= 16'b0000_0000_0000_0000;
array[32703] <= 16'b0000_0000_0000_0000;
array[32704] <= 16'b0000_0000_0000_0000;
array[32705] <= 16'b0000_0000_0000_0000;
array[32706] <= 16'b0000_0000_0000_0000;
array[32707] <= 16'b0000_0000_0000_0000;
array[32708] <= 16'b0000_0000_0000_0000;
array[32709] <= 16'b0000_0000_0000_0000;
array[32710] <= 16'b0000_0000_0000_0000;
array[32711] <= 16'b0000_0000_0000_0000;
array[32712] <= 16'b0000_0000_0000_0000;
array[32713] <= 16'b0000_0000_0000_0000;
array[32714] <= 16'b0000_0000_0000_0000;
array[32715] <= 16'b0000_0000_0000_0000;
array[32716] <= 16'b0000_0000_0000_0000;
array[32717] <= 16'b0000_0000_0000_0000;
array[32718] <= 16'b0000_0000_0000_0000;
array[32719] <= 16'b0000_0000_0000_0000;
array[32720] <= 16'b0000_0000_0000_0000;
array[32721] <= 16'b0000_0000_0000_0000;
array[32722] <= 16'b0000_0000_0000_0000;
array[32723] <= 16'b0000_0000_0000_0000;
array[32724] <= 16'b0000_0000_0000_0000;
array[32725] <= 16'b0000_0000_0000_0000;
array[32726] <= 16'b0000_0000_0000_0000;
array[32727] <= 16'b0000_0000_0000_0000;
array[32728] <= 16'b0000_0000_0000_0000;
array[32729] <= 16'b0000_0000_0000_0000;
array[32730] <= 16'b0000_0000_0000_0000;
array[32731] <= 16'b0000_0000_0000_0000;
array[32732] <= 16'b0000_0000_0000_0000;
array[32733] <= 16'b0000_0000_0000_0000;
array[32734] <= 16'b0000_0000_0000_0000;
array[32735] <= 16'b0000_0000_0000_0000;
array[32736] <= 16'b0000_0000_0000_0000;
array[32737] <= 16'b0000_0000_0000_0000;
array[32738] <= 16'b0000_0000_0000_0000;
array[32739] <= 16'b0000_0000_0000_0000;
array[32740] <= 16'b0000_0000_0000_0000;
array[32741] <= 16'b0000_0000_0000_0000;
array[32742] <= 16'b0000_0000_0000_0000;
array[32743] <= 16'b0000_0000_0000_0000;
array[32744] <= 16'b0000_0000_0000_0000;
array[32745] <= 16'b0000_0000_0000_0000;
array[32746] <= 16'b0000_0000_0000_0000;
array[32747] <= 16'b0000_0000_0000_0000;
array[32748] <= 16'b0000_0000_0000_0000;
array[32749] <= 16'b0000_0000_0000_0000;
array[32750] <= 16'b0000_0000_0000_0000;
array[32751] <= 16'b0000_0000_0000_0000;
array[32752] <= 16'b0000_0000_0000_0000;
array[32753] <= 16'b0000_0000_0000_0000;
array[32754] <= 16'b0000_0000_0000_0000;
array[32755] <= 16'b0000_0000_0000_0000;
array[32756] <= 16'b0000_0000_0000_0000;
array[32757] <= 16'b0000_0000_0000_0000;
array[32758] <= 16'b0000_0000_0000_0000;
array[32759] <= 16'b0000_0000_0000_0000;
array[32760] <= 16'b0000_0000_0000_0000;
array[32761] <= 16'b0000_0000_0000_0000;
array[32762] <= 16'b0000_0000_0000_0000;
array[32763] <= 16'b0000_0000_0000_0000;
array[32764] <= 16'b0000_0000_0000_0000;
array[32765] <= 16'b0000_0000_0000_0000;
array[32766] <= 16'b0000_0000_0000_0000;
array[32767] <= 16'b0000_0000_0000_0000;
array[32768] <= 16'b0000_0000_0000_0000;
array[32769] <= 16'b0000_0000_0000_0000;
array[32770] <= 16'b0000_0000_0000_0000;
array[32771] <= 16'b0000_0000_0000_0000;
array[32772] <= 16'b0000_0000_0000_0000;
array[32773] <= 16'b0000_0000_0000_0000;
array[32774] <= 16'b0000_0000_0000_0000;
array[32775] <= 16'b0000_0000_0000_0000;
array[32776] <= 16'b0000_0000_0000_0000;
array[32777] <= 16'b0000_0000_0000_0000;
array[32778] <= 16'b0000_0000_0000_0000;
array[32779] <= 16'b0000_0000_0000_0000;
array[32780] <= 16'b0000_0000_0000_0000;
array[32781] <= 16'b0000_0000_0000_0000;
array[32782] <= 16'b0000_0000_0000_0000;
array[32783] <= 16'b0000_0000_0000_0000;
array[32784] <= 16'b0000_0000_0000_0000;
array[32785] <= 16'b0000_0000_0000_0000;
array[32786] <= 16'b0000_0000_0000_0000;
array[32787] <= 16'b0000_0000_0000_0000;
array[32788] <= 16'b0000_0000_0000_0000;
array[32789] <= 16'b0000_0000_0000_0000;
array[32790] <= 16'b0000_0000_0000_0000;
array[32791] <= 16'b0000_0000_0000_0000;
array[32792] <= 16'b0000_0000_0000_0000;
array[32793] <= 16'b0000_0000_0000_0000;
array[32794] <= 16'b0000_0000_0000_0000;
array[32795] <= 16'b0000_0000_0000_0000;
array[32796] <= 16'b0000_0000_0000_0000;
array[32797] <= 16'b0000_0000_0000_0000;
array[32798] <= 16'b0000_0000_0000_0000;
array[32799] <= 16'b0000_0000_0000_0000;
array[32800] <= 16'b0000_0000_0000_0000;
array[32801] <= 16'b0000_0000_0000_0000;
array[32802] <= 16'b0000_0000_0000_0000;
array[32803] <= 16'b0000_0000_0000_0000;
array[32804] <= 16'b0000_0000_0000_0000;
array[32805] <= 16'b0000_0000_0000_0000;
array[32806] <= 16'b0000_0000_0000_0000;
array[32807] <= 16'b0000_0000_0000_0000;
array[32808] <= 16'b0000_0000_0000_0000;
array[32809] <= 16'b0000_0000_0000_0000;
array[32810] <= 16'b0000_0000_0000_0000;
array[32811] <= 16'b0000_0000_0000_0000;
array[32812] <= 16'b0000_0000_0000_0000;
array[32813] <= 16'b0000_0000_0000_0000;
array[32814] <= 16'b0000_0000_0000_0000;
array[32815] <= 16'b0000_0000_0000_0000;
array[32816] <= 16'b0000_0000_0000_0000;
array[32817] <= 16'b0000_0000_0000_0000;
array[32818] <= 16'b0000_0000_0000_0000;
array[32819] <= 16'b0000_0000_0000_0000;
array[32820] <= 16'b0000_0000_0000_0000;
array[32821] <= 16'b0000_0000_0000_0000;
array[32822] <= 16'b0000_0000_0000_0000;
array[32823] <= 16'b0000_0000_0000_0000;
array[32824] <= 16'b0000_0000_0000_0000;
array[32825] <= 16'b0000_0000_0000_0000;
array[32826] <= 16'b0000_0000_0000_0000;
array[32827] <= 16'b0000_0000_0000_0000;
array[32828] <= 16'b0000_0000_0000_0000;
array[32829] <= 16'b0000_0000_0000_0000;
array[32830] <= 16'b0000_0000_0000_0000;
array[32831] <= 16'b0000_0000_0000_0000;
array[32832] <= 16'b0000_0000_0000_0000;
array[32833] <= 16'b0000_0000_0000_0000;
array[32834] <= 16'b0000_0000_0000_0000;
array[32835] <= 16'b0000_0000_0000_0000;
array[32836] <= 16'b0000_0000_0000_0000;
array[32837] <= 16'b0000_0000_0000_0000;
array[32838] <= 16'b0000_0000_0000_0000;
array[32839] <= 16'b0000_0000_0000_0000;
array[32840] <= 16'b0000_0000_0000_0000;
array[32841] <= 16'b0000_0000_0000_0000;
array[32842] <= 16'b0000_0000_0000_0000;
array[32843] <= 16'b0000_0000_0000_0000;
array[32844] <= 16'b0000_0000_0000_0000;
array[32845] <= 16'b0000_0000_0000_0000;
array[32846] <= 16'b0000_0000_0000_0000;
array[32847] <= 16'b0000_0000_0000_0000;
array[32848] <= 16'b0000_0000_0000_0000;
array[32849] <= 16'b0000_0000_0000_0000;
array[32850] <= 16'b0000_0000_0000_0000;
array[32851] <= 16'b0000_0000_0000_0000;
array[32852] <= 16'b0000_0000_0000_0000;
array[32853] <= 16'b0000_0000_0000_0000;
array[32854] <= 16'b0000_0000_0000_0000;
array[32855] <= 16'b0000_0000_0000_0000;
array[32856] <= 16'b0000_0000_0000_0000;
array[32857] <= 16'b0000_0000_0000_0000;
array[32858] <= 16'b0000_0000_0000_0000;
array[32859] <= 16'b0000_0000_0000_0000;
array[32860] <= 16'b0000_0000_0000_0000;
array[32861] <= 16'b0000_0000_0000_0000;
array[32862] <= 16'b0000_0000_0000_0000;
array[32863] <= 16'b0000_0000_0000_0000;
array[32864] <= 16'b0000_0000_0000_0000;
array[32865] <= 16'b0000_0000_0000_0000;
array[32866] <= 16'b0000_0000_0000_0000;
array[32867] <= 16'b0000_0000_0000_0000;
array[32868] <= 16'b0000_0000_0000_0000;
array[32869] <= 16'b0000_0000_0000_0000;
array[32870] <= 16'b0000_0000_0000_0000;
array[32871] <= 16'b0000_0000_0000_0000;
array[32872] <= 16'b0000_0000_0000_0000;
array[32873] <= 16'b0000_0000_0000_0000;
array[32874] <= 16'b0000_0000_0000_0000;
array[32875] <= 16'b0000_0000_0000_0000;
array[32876] <= 16'b0000_0000_0000_0000;
array[32877] <= 16'b0000_0000_0000_0000;
array[32878] <= 16'b0000_0000_0000_0000;
array[32879] <= 16'b0000_0000_0000_0000;
array[32880] <= 16'b0000_0000_0000_0000;
array[32881] <= 16'b0000_0000_0000_0000;
array[32882] <= 16'b0000_0000_0000_0000;
array[32883] <= 16'b0000_0000_0000_0000;
array[32884] <= 16'b0000_0000_0000_0000;
array[32885] <= 16'b0000_0000_0000_0000;
array[32886] <= 16'b0000_0000_0000_0000;
array[32887] <= 16'b0000_0000_0000_0000;
array[32888] <= 16'b0000_0000_0000_0000;
array[32889] <= 16'b0000_0000_0000_0000;
array[32890] <= 16'b0000_0000_0000_0000;
array[32891] <= 16'b0000_0000_0000_0000;
array[32892] <= 16'b0000_0000_0000_0000;
array[32893] <= 16'b0000_0000_0000_0000;
array[32894] <= 16'b0000_0000_0000_0000;
array[32895] <= 16'b0000_0000_0000_0000;
array[32896] <= 16'b0000_0000_0000_0000;
array[32897] <= 16'b0000_0000_0000_0000;
array[32898] <= 16'b0000_0000_0000_0000;
array[32899] <= 16'b0000_0000_0000_0000;
array[32900] <= 16'b0000_0000_0000_0000;
array[32901] <= 16'b0000_0000_0000_0000;
array[32902] <= 16'b0000_0000_0000_0000;
array[32903] <= 16'b0000_0000_0000_0000;
array[32904] <= 16'b0000_0000_0000_0000;
array[32905] <= 16'b0000_0000_0000_0000;
array[32906] <= 16'b0000_0000_0000_0000;
array[32907] <= 16'b0000_0000_0000_0000;
array[32908] <= 16'b0000_0000_0000_0000;
array[32909] <= 16'b0000_0000_0000_0000;
array[32910] <= 16'b0000_0000_0000_0000;
array[32911] <= 16'b0000_0000_0000_0000;
array[32912] <= 16'b0000_0000_0000_0000;
array[32913] <= 16'b0000_0000_0000_0000;
array[32914] <= 16'b0000_0000_0000_0000;
array[32915] <= 16'b0000_0000_0000_0000;
array[32916] <= 16'b0000_0000_0000_0000;
array[32917] <= 16'b0000_0000_0000_0000;
array[32918] <= 16'b0000_0000_0000_0000;
array[32919] <= 16'b0000_0000_0000_0000;
array[32920] <= 16'b0000_0000_0000_0000;
array[32921] <= 16'b0000_0000_0000_0000;
array[32922] <= 16'b0000_0000_0000_0000;
array[32923] <= 16'b0000_0000_0000_0000;
array[32924] <= 16'b0000_0000_0000_0000;
array[32925] <= 16'b0000_0000_0000_0000;
array[32926] <= 16'b0000_0000_0000_0000;
array[32927] <= 16'b0000_0000_0000_0000;
array[32928] <= 16'b0000_0000_0000_0000;
array[32929] <= 16'b0000_0000_0000_0000;
array[32930] <= 16'b0000_0000_0000_0000;
array[32931] <= 16'b0000_0000_0000_0000;
array[32932] <= 16'b0000_0000_0000_0000;
array[32933] <= 16'b0000_0000_0000_0000;
array[32934] <= 16'b0000_0000_0000_0000;
array[32935] <= 16'b0000_0000_0000_0000;
array[32936] <= 16'b0000_0000_0000_0000;
array[32937] <= 16'b0000_0000_0000_0000;
array[32938] <= 16'b0000_0000_0000_0000;
array[32939] <= 16'b0000_0000_0000_0000;
array[32940] <= 16'b0000_0000_0000_0000;
array[32941] <= 16'b0000_0000_0000_0000;
array[32942] <= 16'b0000_0000_0000_0000;
array[32943] <= 16'b0000_0000_0000_0000;
array[32944] <= 16'b0000_0000_0000_0000;
array[32945] <= 16'b0000_0000_0000_0000;
array[32946] <= 16'b0000_0000_0000_0000;
array[32947] <= 16'b0000_0000_0000_0000;
array[32948] <= 16'b0000_0000_0000_0000;
array[32949] <= 16'b0000_0000_0000_0000;
array[32950] <= 16'b0000_0000_0000_0000;
array[32951] <= 16'b0000_0000_0000_0000;
array[32952] <= 16'b0000_0000_0000_0000;
array[32953] <= 16'b0000_0000_0000_0000;
array[32954] <= 16'b0000_0000_0000_0000;
array[32955] <= 16'b0000_0000_0000_0000;
array[32956] <= 16'b0000_0000_0000_0000;
array[32957] <= 16'b0000_0000_0000_0000;
array[32958] <= 16'b0000_0000_0000_0000;
array[32959] <= 16'b0000_0000_0000_0000;
array[32960] <= 16'b0000_0000_0000_0000;
array[32961] <= 16'b0000_0000_0000_0000;
array[32962] <= 16'b0000_0000_0000_0000;
array[32963] <= 16'b0000_0000_0000_0000;
array[32964] <= 16'b0000_0000_0000_0000;
array[32965] <= 16'b0000_0000_0000_0000;
array[32966] <= 16'b0000_0000_0000_0000;
array[32967] <= 16'b0000_0000_0000_0000;
array[32968] <= 16'b0000_0000_0000_0000;
array[32969] <= 16'b0000_0000_0000_0000;
array[32970] <= 16'b0000_0000_0000_0000;
array[32971] <= 16'b0000_0000_0000_0000;
array[32972] <= 16'b0000_0000_0000_0000;
array[32973] <= 16'b0000_0000_0000_0000;
array[32974] <= 16'b0000_0000_0000_0000;
array[32975] <= 16'b0000_0000_0000_0000;
array[32976] <= 16'b0000_0000_0000_0000;
array[32977] <= 16'b0000_0000_0000_0000;
array[32978] <= 16'b0000_0000_0000_0000;
array[32979] <= 16'b0000_0000_0000_0000;
array[32980] <= 16'b0000_0000_0000_0000;
array[32981] <= 16'b0000_0000_0000_0000;
array[32982] <= 16'b0000_0000_0000_0000;
array[32983] <= 16'b0000_0000_0000_0000;
array[32984] <= 16'b0000_0000_0000_0000;
array[32985] <= 16'b0000_0000_0000_0000;
array[32986] <= 16'b0000_0000_0000_0000;
array[32987] <= 16'b0000_0000_0000_0000;
array[32988] <= 16'b0000_0000_0000_0000;
array[32989] <= 16'b0000_0000_0000_0000;
array[32990] <= 16'b0000_0000_0000_0000;
array[32991] <= 16'b0000_0000_0000_0000;
array[32992] <= 16'b0000_0000_0000_0000;
array[32993] <= 16'b0000_0000_0000_0000;
array[32994] <= 16'b0000_0000_0000_0000;
array[32995] <= 16'b0000_0000_0000_0000;
array[32996] <= 16'b0000_0000_0000_0000;
array[32997] <= 16'b0000_0000_0000_0000;
array[32998] <= 16'b0000_0000_0000_0000;
array[32999] <= 16'b0000_0000_0000_0000;
array[33000] <= 16'b0000_0000_0000_0000;
array[33001] <= 16'b0000_0000_0000_0000;
array[33002] <= 16'b0000_0000_0000_0000;
array[33003] <= 16'b0000_0000_0000_0000;
array[33004] <= 16'b0000_0000_0000_0000;
array[33005] <= 16'b0000_0000_0000_0000;
array[33006] <= 16'b0000_0000_0000_0000;
array[33007] <= 16'b0000_0000_0000_0000;
array[33008] <= 16'b0000_0000_0000_0000;
array[33009] <= 16'b0000_0000_0000_0000;
array[33010] <= 16'b0000_0000_0000_0000;
array[33011] <= 16'b0000_0000_0000_0000;
array[33012] <= 16'b0000_0000_0000_0000;
array[33013] <= 16'b0000_0000_0000_0000;
array[33014] <= 16'b0000_0000_0000_0000;
array[33015] <= 16'b0000_0000_0000_0000;
array[33016] <= 16'b0000_0000_0000_0000;
array[33017] <= 16'b0000_0000_0000_0000;
array[33018] <= 16'b0000_0000_0000_0000;
array[33019] <= 16'b0000_0000_0000_0000;
array[33020] <= 16'b0000_0000_0000_0000;
array[33021] <= 16'b0000_0000_0000_0000;
array[33022] <= 16'b0000_0000_0000_0000;
array[33023] <= 16'b0000_0000_0000_0000;
array[33024] <= 16'b0000_0000_0000_0000;
array[33025] <= 16'b0000_0000_0000_0000;
array[33026] <= 16'b0000_0000_0000_0000;
array[33027] <= 16'b0000_0000_0000_0000;
array[33028] <= 16'b0000_0000_0000_0000;
array[33029] <= 16'b0000_0000_0000_0000;
array[33030] <= 16'b0000_0000_0000_0000;
array[33031] <= 16'b0000_0000_0000_0000;
array[33032] <= 16'b0000_0000_0000_0000;
array[33033] <= 16'b0000_0000_0000_0000;
array[33034] <= 16'b0000_0000_0000_0000;
array[33035] <= 16'b0000_0000_0000_0000;
array[33036] <= 16'b0000_0000_0000_0000;
array[33037] <= 16'b0000_0000_0000_0000;
array[33038] <= 16'b0000_0000_0000_0000;
array[33039] <= 16'b0000_0000_0000_0000;
array[33040] <= 16'b0000_0000_0000_0000;
array[33041] <= 16'b0000_0000_0000_0000;
array[33042] <= 16'b0000_0000_0000_0000;
array[33043] <= 16'b0000_0000_0000_0000;
array[33044] <= 16'b0000_0000_0000_0000;
array[33045] <= 16'b0000_0000_0000_0000;
array[33046] <= 16'b0000_0000_0000_0000;
array[33047] <= 16'b0000_0000_0000_0000;
array[33048] <= 16'b0000_0000_0000_0000;
array[33049] <= 16'b0000_0000_0000_0000;
array[33050] <= 16'b0000_0000_0000_0000;
array[33051] <= 16'b0000_0000_0000_0000;
array[33052] <= 16'b0000_0000_0000_0000;
array[33053] <= 16'b0000_0000_0000_0000;
array[33054] <= 16'b0000_0000_0000_0000;
array[33055] <= 16'b0000_0000_0000_0000;
array[33056] <= 16'b0000_0000_0000_0000;
array[33057] <= 16'b0000_0000_0000_0000;
array[33058] <= 16'b0000_0000_0000_0000;
array[33059] <= 16'b0000_0000_0000_0000;
array[33060] <= 16'b0000_0000_0000_0000;
array[33061] <= 16'b0000_0000_0000_0000;
array[33062] <= 16'b0000_0000_0000_0000;
array[33063] <= 16'b0000_0000_0000_0000;
array[33064] <= 16'b0000_0000_0000_0000;
array[33065] <= 16'b0000_0000_0000_0000;
array[33066] <= 16'b0000_0000_0000_0000;
array[33067] <= 16'b0000_0000_0000_0000;
array[33068] <= 16'b0000_0000_0000_0000;
array[33069] <= 16'b0000_0000_0000_0000;
array[33070] <= 16'b0000_0000_0000_0000;
array[33071] <= 16'b0000_0000_0000_0000;
array[33072] <= 16'b0000_0000_0000_0000;
array[33073] <= 16'b0000_0000_0000_0000;
array[33074] <= 16'b0000_0000_0000_0000;
array[33075] <= 16'b0000_0000_0000_0000;
array[33076] <= 16'b0000_0000_0000_0000;
array[33077] <= 16'b0000_0000_0000_0000;
array[33078] <= 16'b0000_0000_0000_0000;
array[33079] <= 16'b0000_0000_0000_0000;
array[33080] <= 16'b0000_0000_0000_0000;
array[33081] <= 16'b0000_0000_0000_0000;
array[33082] <= 16'b0000_0000_0000_0000;
array[33083] <= 16'b0000_0000_0000_0000;
array[33084] <= 16'b0000_0000_0000_0000;
array[33085] <= 16'b0000_0000_0000_0000;
array[33086] <= 16'b0000_0000_0000_0000;
array[33087] <= 16'b0000_0000_0000_0000;
array[33088] <= 16'b0000_0000_0000_0000;
array[33089] <= 16'b0000_0000_0000_0000;
array[33090] <= 16'b0000_0000_0000_0000;
array[33091] <= 16'b0000_0000_0000_0000;
array[33092] <= 16'b0000_0000_0000_0000;
array[33093] <= 16'b0000_0000_0000_0000;
array[33094] <= 16'b0000_0000_0000_0000;
array[33095] <= 16'b0000_0000_0000_0000;
array[33096] <= 16'b0000_0000_0000_0000;
array[33097] <= 16'b0000_0000_0000_0000;
array[33098] <= 16'b0000_0000_0000_0000;
array[33099] <= 16'b0000_0000_0000_0000;
array[33100] <= 16'b0000_0000_0000_0000;
array[33101] <= 16'b0000_0000_0000_0000;
array[33102] <= 16'b0000_0000_0000_0000;
array[33103] <= 16'b0000_0000_0000_0000;
array[33104] <= 16'b0000_0000_0000_0000;
array[33105] <= 16'b0000_0000_0000_0000;
array[33106] <= 16'b0000_0000_0000_0000;
array[33107] <= 16'b0000_0000_0000_0000;
array[33108] <= 16'b0000_0000_0000_0000;
array[33109] <= 16'b0000_0000_0000_0000;
array[33110] <= 16'b0000_0000_0000_0000;
array[33111] <= 16'b0000_0000_0000_0000;
array[33112] <= 16'b0000_0000_0000_0000;
array[33113] <= 16'b0000_0000_0000_0000;
array[33114] <= 16'b0000_0000_0000_0000;
array[33115] <= 16'b0000_0000_0000_0000;
array[33116] <= 16'b0000_0000_0000_0000;
array[33117] <= 16'b0000_0000_0000_0000;
array[33118] <= 16'b0000_0000_0000_0000;
array[33119] <= 16'b0000_0000_0000_0000;
array[33120] <= 16'b0000_0000_0000_0000;
array[33121] <= 16'b0000_0000_0000_0000;
array[33122] <= 16'b0000_0000_0000_0000;
array[33123] <= 16'b0000_0000_0000_0000;
array[33124] <= 16'b0000_0000_0000_0000;
array[33125] <= 16'b0000_0000_0000_0000;
array[33126] <= 16'b0000_0000_0000_0000;
array[33127] <= 16'b0000_0000_0000_0000;
array[33128] <= 16'b0000_0000_0000_0000;
array[33129] <= 16'b0000_0000_0000_0000;
array[33130] <= 16'b0000_0000_0000_0000;
array[33131] <= 16'b0000_0000_0000_0000;
array[33132] <= 16'b0000_0000_0000_0000;
array[33133] <= 16'b0000_0000_0000_0000;
array[33134] <= 16'b0000_0000_0000_0000;
array[33135] <= 16'b0000_0000_0000_0000;
array[33136] <= 16'b0000_0000_0000_0000;
array[33137] <= 16'b0000_0000_0000_0000;
array[33138] <= 16'b0000_0000_0000_0000;
array[33139] <= 16'b0000_0000_0000_0000;
array[33140] <= 16'b0000_0000_0000_0000;
array[33141] <= 16'b0000_0000_0000_0000;
array[33142] <= 16'b0000_0000_0000_0000;
array[33143] <= 16'b0000_0000_0000_0000;
array[33144] <= 16'b0000_0000_0000_0000;
array[33145] <= 16'b0000_0000_0000_0000;
array[33146] <= 16'b0000_0000_0000_0000;
array[33147] <= 16'b0000_0000_0000_0000;
array[33148] <= 16'b0000_0000_0000_0000;
array[33149] <= 16'b0000_0000_0000_0000;
array[33150] <= 16'b0000_0000_0000_0000;
array[33151] <= 16'b0000_0000_0000_0000;
array[33152] <= 16'b0000_0000_0000_0000;
array[33153] <= 16'b0000_0000_0000_0000;
array[33154] <= 16'b0000_0000_0000_0000;
array[33155] <= 16'b0000_0000_0000_0000;
array[33156] <= 16'b0000_0000_0000_0000;
array[33157] <= 16'b0000_0000_0000_0000;
array[33158] <= 16'b0000_0000_0000_0000;
array[33159] <= 16'b0000_0000_0000_0000;
array[33160] <= 16'b0000_0000_0000_0000;
array[33161] <= 16'b0000_0000_0000_0000;
array[33162] <= 16'b0000_0000_0000_0000;
array[33163] <= 16'b0000_0000_0000_0000;
array[33164] <= 16'b0000_0000_0000_0000;
array[33165] <= 16'b0000_0000_0000_0000;
array[33166] <= 16'b0000_0000_0000_0000;
array[33167] <= 16'b0000_0000_0000_0000;
array[33168] <= 16'b0000_0000_0000_0000;
array[33169] <= 16'b0000_0000_0000_0000;
array[33170] <= 16'b0000_0000_0000_0000;
array[33171] <= 16'b0000_0000_0000_0000;
array[33172] <= 16'b0000_0000_0000_0000;
array[33173] <= 16'b0000_0000_0000_0000;
array[33174] <= 16'b0000_0000_0000_0000;
array[33175] <= 16'b0000_0000_0000_0000;
array[33176] <= 16'b0000_0000_0000_0000;
array[33177] <= 16'b0000_0000_0000_0000;
array[33178] <= 16'b0000_0000_0000_0000;
array[33179] <= 16'b0000_0000_0000_0000;
array[33180] <= 16'b0000_0000_0000_0000;
array[33181] <= 16'b0000_0000_0000_0000;
array[33182] <= 16'b0000_0000_0000_0000;
array[33183] <= 16'b0000_0000_0000_0000;
array[33184] <= 16'b0000_0000_0000_0000;
array[33185] <= 16'b0000_0000_0000_0000;
array[33186] <= 16'b0000_0000_0000_0000;
array[33187] <= 16'b0000_0000_0000_0000;
array[33188] <= 16'b0000_0000_0000_0000;
array[33189] <= 16'b0000_0000_0000_0000;
array[33190] <= 16'b0000_0000_0000_0000;
array[33191] <= 16'b0000_0000_0000_0000;
array[33192] <= 16'b0000_0000_0000_0000;
array[33193] <= 16'b0000_0000_0000_0000;
array[33194] <= 16'b0000_0000_0000_0000;
array[33195] <= 16'b0000_0000_0000_0000;
array[33196] <= 16'b0000_0000_0000_0000;
array[33197] <= 16'b0000_0000_0000_0000;
array[33198] <= 16'b0000_0000_0000_0000;
array[33199] <= 16'b0000_0000_0000_0000;
array[33200] <= 16'b0000_0000_0000_0000;
array[33201] <= 16'b0000_0000_0000_0000;
array[33202] <= 16'b0000_0000_0000_0000;
array[33203] <= 16'b0000_0000_0000_0000;
array[33204] <= 16'b0000_0000_0000_0000;
array[33205] <= 16'b0000_0000_0000_0000;
array[33206] <= 16'b0000_0000_0000_0000;
array[33207] <= 16'b0000_0000_0000_0000;
array[33208] <= 16'b0000_0000_0000_0000;
array[33209] <= 16'b0000_0000_0000_0000;
array[33210] <= 16'b0000_0000_0000_0000;
array[33211] <= 16'b0000_0000_0000_0000;
array[33212] <= 16'b0000_0000_0000_0000;
array[33213] <= 16'b0000_0000_0000_0000;
array[33214] <= 16'b0000_0000_0000_0000;
array[33215] <= 16'b0000_0000_0000_0000;
array[33216] <= 16'b0000_0000_0000_0000;
array[33217] <= 16'b0000_0000_0000_0000;
array[33218] <= 16'b0000_0000_0000_0000;
array[33219] <= 16'b0000_0000_0000_0000;
array[33220] <= 16'b0000_0000_0000_0000;
array[33221] <= 16'b0000_0000_0000_0000;
array[33222] <= 16'b0000_0000_0000_0000;
array[33223] <= 16'b0000_0000_0000_0000;
array[33224] <= 16'b0000_0000_0000_0000;
array[33225] <= 16'b0000_0000_0000_0000;
array[33226] <= 16'b0000_0000_0000_0000;
array[33227] <= 16'b0000_0000_0000_0000;
array[33228] <= 16'b0000_0000_0000_0000;
array[33229] <= 16'b0000_0000_0000_0000;
array[33230] <= 16'b0000_0000_0000_0000;
array[33231] <= 16'b0000_0000_0000_0000;
array[33232] <= 16'b0000_0000_0000_0000;
array[33233] <= 16'b0000_0000_0000_0000;
array[33234] <= 16'b0000_0000_0000_0000;
array[33235] <= 16'b0000_0000_0000_0000;
array[33236] <= 16'b0000_0000_0000_0000;
array[33237] <= 16'b0000_0000_0000_0000;
array[33238] <= 16'b0000_0000_0000_0000;
array[33239] <= 16'b0000_0000_0000_0000;
array[33240] <= 16'b0000_0000_0000_0000;
array[33241] <= 16'b0000_0000_0000_0000;
array[33242] <= 16'b0000_0000_0000_0000;
array[33243] <= 16'b0000_0000_0000_0000;
array[33244] <= 16'b0000_0000_0000_0000;
array[33245] <= 16'b0000_0000_0000_0000;
array[33246] <= 16'b0000_0000_0000_0000;
array[33247] <= 16'b0000_0000_0000_0000;
array[33248] <= 16'b0000_0000_0000_0000;
array[33249] <= 16'b0000_0000_0000_0000;
array[33250] <= 16'b0000_0000_0000_0000;
array[33251] <= 16'b0000_0000_0000_0000;
array[33252] <= 16'b0000_0000_0000_0000;
array[33253] <= 16'b0000_0000_0000_0000;
array[33254] <= 16'b0000_0000_0000_0000;
array[33255] <= 16'b0000_0000_0000_0000;
array[33256] <= 16'b0000_0000_0000_0000;
array[33257] <= 16'b0000_0000_0000_0000;
array[33258] <= 16'b0000_0000_0000_0000;
array[33259] <= 16'b0000_0000_0000_0000;
array[33260] <= 16'b0000_0000_0000_0000;
array[33261] <= 16'b0000_0000_0000_0000;
array[33262] <= 16'b0000_0000_0000_0000;
array[33263] <= 16'b0000_0000_0000_0000;
array[33264] <= 16'b0000_0000_0000_0000;
array[33265] <= 16'b0000_0000_0000_0000;
array[33266] <= 16'b0000_0000_0000_0000;
array[33267] <= 16'b0000_0000_0000_0000;
array[33268] <= 16'b0000_0000_0000_0000;
array[33269] <= 16'b0000_0000_0000_0000;
array[33270] <= 16'b0000_0000_0000_0000;
array[33271] <= 16'b0000_0000_0000_0000;
array[33272] <= 16'b0000_0000_0000_0000;
array[33273] <= 16'b0000_0000_0000_0000;
array[33274] <= 16'b0000_0000_0000_0000;
array[33275] <= 16'b0000_0000_0000_0000;
array[33276] <= 16'b0000_0000_0000_0000;
array[33277] <= 16'b0000_0000_0000_0000;
array[33278] <= 16'b0000_0000_0000_0000;
array[33279] <= 16'b0000_0000_0000_0000;
array[33280] <= 16'b0000_0000_0000_0000;
array[33281] <= 16'b0000_0000_0000_0000;
array[33282] <= 16'b0000_0000_0000_0000;
array[33283] <= 16'b0000_0000_0000_0000;
array[33284] <= 16'b0000_0000_0000_0000;
array[33285] <= 16'b0000_0000_0000_0000;
array[33286] <= 16'b0000_0000_0000_0000;
array[33287] <= 16'b0000_0000_0000_0000;
array[33288] <= 16'b0000_0000_0000_0000;
array[33289] <= 16'b0000_0000_0000_0000;
array[33290] <= 16'b0000_0000_0000_0000;
array[33291] <= 16'b0000_0000_0000_0000;
array[33292] <= 16'b0000_0000_0000_0000;
array[33293] <= 16'b0000_0000_0000_0000;
array[33294] <= 16'b0000_0000_0000_0000;
array[33295] <= 16'b0000_0000_0000_0000;
array[33296] <= 16'b0000_0000_0000_0000;
array[33297] <= 16'b0000_0000_0000_0000;
array[33298] <= 16'b0000_0000_0000_0000;
array[33299] <= 16'b0000_0000_0000_0000;
array[33300] <= 16'b0000_0000_0000_0000;
array[33301] <= 16'b0000_0000_0000_0000;
array[33302] <= 16'b0000_0000_0000_0000;
array[33303] <= 16'b0000_0000_0000_0000;
array[33304] <= 16'b0000_0000_0000_0000;
array[33305] <= 16'b0000_0000_0000_0000;
array[33306] <= 16'b0000_0000_0000_0000;
array[33307] <= 16'b0000_0000_0000_0000;
array[33308] <= 16'b0000_0000_0000_0000;
array[33309] <= 16'b0000_0000_0000_0000;
array[33310] <= 16'b0000_0000_0000_0000;
array[33311] <= 16'b0000_0000_0000_0000;
array[33312] <= 16'b0000_0000_0000_0000;
array[33313] <= 16'b0000_0000_0000_0000;
array[33314] <= 16'b0000_0000_0000_0000;
array[33315] <= 16'b0000_0000_0000_0000;
array[33316] <= 16'b0000_0000_0000_0000;
array[33317] <= 16'b0000_0000_0000_0000;
array[33318] <= 16'b0000_0000_0000_0000;
array[33319] <= 16'b0000_0000_0000_0000;
array[33320] <= 16'b0000_0000_0000_0000;
array[33321] <= 16'b0000_0000_0000_0000;
array[33322] <= 16'b0000_0000_0000_0000;
array[33323] <= 16'b0000_0000_0000_0000;
array[33324] <= 16'b0000_0000_0000_0000;
array[33325] <= 16'b0000_0000_0000_0000;
array[33326] <= 16'b0000_0000_0000_0000;
array[33327] <= 16'b0000_0000_0000_0000;
array[33328] <= 16'b0000_0000_0000_0000;
array[33329] <= 16'b0000_0000_0000_0000;
array[33330] <= 16'b0000_0000_0000_0000;
array[33331] <= 16'b0000_0000_0000_0000;
array[33332] <= 16'b0000_0000_0000_0000;
array[33333] <= 16'b0000_0000_0000_0000;
array[33334] <= 16'b0000_0000_0000_0000;
array[33335] <= 16'b0000_0000_0000_0000;
array[33336] <= 16'b0000_0000_0000_0000;
array[33337] <= 16'b0000_0000_0000_0000;
array[33338] <= 16'b0000_0000_0000_0000;
array[33339] <= 16'b0000_0000_0000_0000;
array[33340] <= 16'b0000_0000_0000_0000;
array[33341] <= 16'b0000_0000_0000_0000;
array[33342] <= 16'b0000_0000_0000_0000;
array[33343] <= 16'b0000_0000_0000_0000;
array[33344] <= 16'b0000_0000_0000_0000;
array[33345] <= 16'b0000_0000_0000_0000;
array[33346] <= 16'b0000_0000_0000_0000;
array[33347] <= 16'b0000_0000_0000_0000;
array[33348] <= 16'b0000_0000_0000_0000;
array[33349] <= 16'b0000_0000_0000_0000;
array[33350] <= 16'b0000_0000_0000_0000;
array[33351] <= 16'b0000_0000_0000_0000;
array[33352] <= 16'b0000_0000_0000_0000;
array[33353] <= 16'b0000_0000_0000_0000;
array[33354] <= 16'b0000_0000_0000_0000;
array[33355] <= 16'b0000_0000_0000_0000;
array[33356] <= 16'b0000_0000_0000_0000;
array[33357] <= 16'b0000_0000_0000_0000;
array[33358] <= 16'b0000_0000_0000_0000;
array[33359] <= 16'b0000_0000_0000_0000;
array[33360] <= 16'b0000_0000_0000_0000;
array[33361] <= 16'b0000_0000_0000_0000;
array[33362] <= 16'b0000_0000_0000_0000;
array[33363] <= 16'b0000_0000_0000_0000;
array[33364] <= 16'b0000_0000_0000_0000;
array[33365] <= 16'b0000_0000_0000_0000;
array[33366] <= 16'b0000_0000_0000_0000;
array[33367] <= 16'b0000_0000_0000_0000;
array[33368] <= 16'b0000_0000_0000_0000;
array[33369] <= 16'b0000_0000_0000_0000;
array[33370] <= 16'b0000_0000_0000_0000;
array[33371] <= 16'b0000_0000_0000_0000;
array[33372] <= 16'b0000_0000_0000_0000;
array[33373] <= 16'b0000_0000_0000_0000;
array[33374] <= 16'b0000_0000_0000_0000;
array[33375] <= 16'b0000_0000_0000_0000;
array[33376] <= 16'b0000_0000_0000_0000;
array[33377] <= 16'b0000_0000_0000_0000;
array[33378] <= 16'b0000_0000_0000_0000;
array[33379] <= 16'b0000_0000_0000_0000;
array[33380] <= 16'b0000_0000_0000_0000;
array[33381] <= 16'b0000_0000_0000_0000;
array[33382] <= 16'b0000_0000_0000_0000;
array[33383] <= 16'b0000_0000_0000_0000;
array[33384] <= 16'b0000_0000_0000_0000;
array[33385] <= 16'b0000_0000_0000_0000;
array[33386] <= 16'b0000_0000_0000_0000;
array[33387] <= 16'b0000_0000_0000_0000;
array[33388] <= 16'b0000_0000_0000_0000;
array[33389] <= 16'b0000_0000_0000_0000;
array[33390] <= 16'b0000_0000_0000_0000;
array[33391] <= 16'b0000_0000_0000_0000;
array[33392] <= 16'b0000_0000_0000_0000;
array[33393] <= 16'b0000_0000_0000_0000;
array[33394] <= 16'b0000_0000_0000_0000;
array[33395] <= 16'b0000_0000_0000_0000;
array[33396] <= 16'b0000_0000_0000_0000;
array[33397] <= 16'b0000_0000_0000_0000;
array[33398] <= 16'b0000_0000_0000_0000;
array[33399] <= 16'b0000_0000_0000_0000;
array[33400] <= 16'b0000_0000_0000_0000;
array[33401] <= 16'b0000_0000_0000_0000;
array[33402] <= 16'b0000_0000_0000_0000;
array[33403] <= 16'b0000_0000_0000_0000;
array[33404] <= 16'b0000_0000_0000_0000;
array[33405] <= 16'b0000_0000_0000_0000;
array[33406] <= 16'b0000_0000_0000_0000;
array[33407] <= 16'b0000_0000_0000_0000;
array[33408] <= 16'b0000_0000_0000_0000;
array[33409] <= 16'b0000_0000_0000_0000;
array[33410] <= 16'b0000_0000_0000_0000;
array[33411] <= 16'b0000_0000_0000_0000;
array[33412] <= 16'b0000_0000_0000_0000;
array[33413] <= 16'b0000_0000_0000_0000;
array[33414] <= 16'b0000_0000_0000_0000;
array[33415] <= 16'b0000_0000_0000_0000;
array[33416] <= 16'b0000_0000_0000_0000;
array[33417] <= 16'b0000_0000_0000_0000;
array[33418] <= 16'b0000_0000_0000_0000;
array[33419] <= 16'b0000_0000_0000_0000;
array[33420] <= 16'b0000_0000_0000_0000;
array[33421] <= 16'b0000_0000_0000_0000;
array[33422] <= 16'b0000_0000_0000_0000;
array[33423] <= 16'b0000_0000_0000_0000;
array[33424] <= 16'b0000_0000_0000_0000;
array[33425] <= 16'b0000_0000_0000_0000;
array[33426] <= 16'b0000_0000_0000_0000;
array[33427] <= 16'b0000_0000_0000_0000;
array[33428] <= 16'b0000_0000_0000_0000;
array[33429] <= 16'b0000_0000_0000_0000;
array[33430] <= 16'b0000_0000_0000_0000;
array[33431] <= 16'b0000_0000_0000_0000;
array[33432] <= 16'b0000_0000_0000_0000;
array[33433] <= 16'b0000_0000_0000_0000;
array[33434] <= 16'b0000_0000_0000_0000;
array[33435] <= 16'b0000_0000_0000_0000;
array[33436] <= 16'b0000_0000_0000_0000;
array[33437] <= 16'b0000_0000_0000_0000;
array[33438] <= 16'b0000_0000_0000_0000;
array[33439] <= 16'b0000_0000_0000_0000;
array[33440] <= 16'b0000_0000_0000_0000;
array[33441] <= 16'b0000_0000_0000_0000;
array[33442] <= 16'b0000_0000_0000_0000;
array[33443] <= 16'b0000_0000_0000_0000;
array[33444] <= 16'b0000_0000_0000_0000;
array[33445] <= 16'b0000_0000_0000_0000;
array[33446] <= 16'b0000_0000_0000_0000;
array[33447] <= 16'b0000_0000_0000_0000;
array[33448] <= 16'b0000_0000_0000_0000;
array[33449] <= 16'b0000_0000_0000_0000;
array[33450] <= 16'b0000_0000_0000_0000;
array[33451] <= 16'b0000_0000_0000_0000;
array[33452] <= 16'b0000_0000_0000_0000;
array[33453] <= 16'b0000_0000_0000_0000;
array[33454] <= 16'b0000_0000_0000_0000;
array[33455] <= 16'b0000_0000_0000_0000;
array[33456] <= 16'b0000_0000_0000_0000;
array[33457] <= 16'b0000_0000_0000_0000;
array[33458] <= 16'b0000_0000_0000_0000;
array[33459] <= 16'b0000_0000_0000_0000;
array[33460] <= 16'b0000_0000_0000_0000;
array[33461] <= 16'b0000_0000_0000_0000;
array[33462] <= 16'b0000_0000_0000_0000;
array[33463] <= 16'b0000_0000_0000_0000;
array[33464] <= 16'b0000_0000_0000_0000;
array[33465] <= 16'b0000_0000_0000_0000;
array[33466] <= 16'b0000_0000_0000_0000;
array[33467] <= 16'b0000_0000_0000_0000;
array[33468] <= 16'b0000_0000_0000_0000;
array[33469] <= 16'b0000_0000_0000_0000;
array[33470] <= 16'b0000_0000_0000_0000;
array[33471] <= 16'b0000_0000_0000_0000;
array[33472] <= 16'b0000_0000_0000_0000;
array[33473] <= 16'b0000_0000_0000_0000;
array[33474] <= 16'b0000_0000_0000_0000;
array[33475] <= 16'b0000_0000_0000_0000;
array[33476] <= 16'b0000_0000_0000_0000;
array[33477] <= 16'b0000_0000_0000_0000;
array[33478] <= 16'b0000_0000_0000_0000;
array[33479] <= 16'b0000_0000_0000_0000;
array[33480] <= 16'b0000_0000_0000_0000;
array[33481] <= 16'b0000_0000_0000_0000;
array[33482] <= 16'b0000_0000_0000_0000;
array[33483] <= 16'b0000_0000_0000_0000;
array[33484] <= 16'b0000_0000_0000_0000;
array[33485] <= 16'b0000_0000_0000_0000;
array[33486] <= 16'b0000_0000_0000_0000;
array[33487] <= 16'b0000_0000_0000_0000;
array[33488] <= 16'b0000_0000_0000_0000;
array[33489] <= 16'b0000_0000_0000_0000;
array[33490] <= 16'b0000_0000_0000_0000;
array[33491] <= 16'b0000_0000_0000_0000;
array[33492] <= 16'b0000_0000_0000_0000;
array[33493] <= 16'b0000_0000_0000_0000;
array[33494] <= 16'b0000_0000_0000_0000;
array[33495] <= 16'b0000_0000_0000_0000;
array[33496] <= 16'b0000_0000_0000_0000;
array[33497] <= 16'b0000_0000_0000_0000;
array[33498] <= 16'b0000_0000_0000_0000;
array[33499] <= 16'b0000_0000_0000_0000;
array[33500] <= 16'b0000_0000_0000_0000;
array[33501] <= 16'b0000_0000_0000_0000;
array[33502] <= 16'b0000_0000_0000_0000;
array[33503] <= 16'b0000_0000_0000_0000;
array[33504] <= 16'b0000_0000_0000_0000;
array[33505] <= 16'b0000_0000_0000_0000;
array[33506] <= 16'b0000_0000_0000_0000;
array[33507] <= 16'b0000_0000_0000_0000;
array[33508] <= 16'b0000_0000_0000_0000;
array[33509] <= 16'b0000_0000_0000_0000;
array[33510] <= 16'b0000_0000_0000_0000;
array[33511] <= 16'b0000_0000_0000_0000;
array[33512] <= 16'b0000_0000_0000_0000;
array[33513] <= 16'b0000_0000_0000_0000;
array[33514] <= 16'b0000_0000_0000_0000;
array[33515] <= 16'b0000_0000_0000_0000;
array[33516] <= 16'b0000_0000_0000_0000;
array[33517] <= 16'b0000_0000_0000_0000;
array[33518] <= 16'b0000_0000_0000_0000;
array[33519] <= 16'b0000_0000_0000_0000;
array[33520] <= 16'b0000_0000_0000_0000;
array[33521] <= 16'b0000_0000_0000_0000;
array[33522] <= 16'b0000_0000_0000_0000;
array[33523] <= 16'b0000_0000_0000_0000;
array[33524] <= 16'b0000_0000_0000_0000;
array[33525] <= 16'b0000_0000_0000_0000;
array[33526] <= 16'b0000_0000_0000_0000;
array[33527] <= 16'b0000_0000_0000_0000;
array[33528] <= 16'b0000_0000_0000_0000;
array[33529] <= 16'b0000_0000_0000_0000;
array[33530] <= 16'b0000_0000_0000_0000;
array[33531] <= 16'b0000_0000_0000_0000;
array[33532] <= 16'b0000_0000_0000_0000;
array[33533] <= 16'b0000_0000_0000_0000;
array[33534] <= 16'b0000_0000_0000_0000;
array[33535] <= 16'b0000_0000_0000_0000;
array[33536] <= 16'b0000_0000_0000_0000;
array[33537] <= 16'b0000_0000_0000_0000;
array[33538] <= 16'b0000_0000_0000_0000;
array[33539] <= 16'b0000_0000_0000_0000;
array[33540] <= 16'b0000_0000_0000_0000;
array[33541] <= 16'b0000_0000_0000_0000;
array[33542] <= 16'b0000_0000_0000_0000;
array[33543] <= 16'b0000_0000_0000_0000;
array[33544] <= 16'b0000_0000_0000_0000;
array[33545] <= 16'b0000_0000_0000_0000;
array[33546] <= 16'b0000_0000_0000_0000;
array[33547] <= 16'b0000_0000_0000_0000;
array[33548] <= 16'b0000_0000_0000_0000;
array[33549] <= 16'b0000_0000_0000_0000;
array[33550] <= 16'b0000_0000_0000_0000;
array[33551] <= 16'b0000_0000_0000_0000;
array[33552] <= 16'b0000_0000_0000_0000;
array[33553] <= 16'b0000_0000_0000_0000;
array[33554] <= 16'b0000_0000_0000_0000;
array[33555] <= 16'b0000_0000_0000_0000;
array[33556] <= 16'b0000_0000_0000_0000;
array[33557] <= 16'b0000_0000_0000_0000;
array[33558] <= 16'b0000_0000_0000_0000;
array[33559] <= 16'b0000_0000_0000_0000;
array[33560] <= 16'b0000_0000_0000_0000;
array[33561] <= 16'b0000_0000_0000_0000;
array[33562] <= 16'b0000_0000_0000_0000;
array[33563] <= 16'b0000_0000_0000_0000;
array[33564] <= 16'b0000_0000_0000_0000;
array[33565] <= 16'b0000_0000_0000_0000;
array[33566] <= 16'b0000_0000_0000_0000;
array[33567] <= 16'b0000_0000_0000_0000;
array[33568] <= 16'b0000_0000_0000_0000;
array[33569] <= 16'b0000_0000_0000_0000;
array[33570] <= 16'b0000_0000_0000_0000;
array[33571] <= 16'b0000_0000_0000_0000;
array[33572] <= 16'b0000_0000_0000_0000;
array[33573] <= 16'b0000_0000_0000_0000;
array[33574] <= 16'b0000_0000_0000_0000;
array[33575] <= 16'b0000_0000_0000_0000;
array[33576] <= 16'b0000_0000_0000_0000;
array[33577] <= 16'b0000_0000_0000_0000;
array[33578] <= 16'b0000_0000_0000_0000;
array[33579] <= 16'b0000_0000_0000_0000;
array[33580] <= 16'b0000_0000_0000_0000;
array[33581] <= 16'b0000_0000_0000_0000;
array[33582] <= 16'b0000_0000_0000_0000;
array[33583] <= 16'b0000_0000_0000_0000;
array[33584] <= 16'b0000_0000_0000_0000;
array[33585] <= 16'b0000_0000_0000_0000;
array[33586] <= 16'b0000_0000_0000_0000;
array[33587] <= 16'b0000_0000_0000_0000;
array[33588] <= 16'b0000_0000_0000_0000;
array[33589] <= 16'b0000_0000_0000_0000;
array[33590] <= 16'b0000_0000_0000_0000;
array[33591] <= 16'b0000_0000_0000_0000;
array[33592] <= 16'b0000_0000_0000_0000;
array[33593] <= 16'b0000_0000_0000_0000;
array[33594] <= 16'b0000_0000_0000_0000;
array[33595] <= 16'b0000_0000_0000_0000;
array[33596] <= 16'b0000_0000_0000_0000;
array[33597] <= 16'b0000_0000_0000_0000;
array[33598] <= 16'b0000_0000_0000_0000;
array[33599] <= 16'b0000_0000_0000_0000;
array[33600] <= 16'b0000_0000_0000_0000;
array[33601] <= 16'b0000_0000_0000_0000;
array[33602] <= 16'b0000_0000_0000_0000;
array[33603] <= 16'b0000_0000_0000_0000;
array[33604] <= 16'b0000_0000_0000_0000;
array[33605] <= 16'b0000_0000_0000_0000;
array[33606] <= 16'b0000_0000_0000_0000;
array[33607] <= 16'b0000_0000_0000_0000;
array[33608] <= 16'b0000_0000_0000_0000;
array[33609] <= 16'b0000_0000_0000_0000;
array[33610] <= 16'b0000_0000_0000_0000;
array[33611] <= 16'b0000_0000_0000_0000;
array[33612] <= 16'b0000_0000_0000_0000;
array[33613] <= 16'b0000_0000_0000_0000;
array[33614] <= 16'b0000_0000_0000_0000;
array[33615] <= 16'b0000_0000_0000_0000;
array[33616] <= 16'b0000_0000_0000_0000;
array[33617] <= 16'b0000_0000_0000_0000;
array[33618] <= 16'b0000_0000_0000_0000;
array[33619] <= 16'b0000_0000_0000_0000;
array[33620] <= 16'b0000_0000_0000_0000;
array[33621] <= 16'b0000_0000_0000_0000;
array[33622] <= 16'b0000_0000_0000_0000;
array[33623] <= 16'b0000_0000_0000_0000;
array[33624] <= 16'b0000_0000_0000_0000;
array[33625] <= 16'b0000_0000_0000_0000;
array[33626] <= 16'b0000_0000_0000_0000;
array[33627] <= 16'b0000_0000_0000_0000;
array[33628] <= 16'b0000_0000_0000_0000;
array[33629] <= 16'b0000_0000_0000_0000;
array[33630] <= 16'b0000_0000_0000_0000;
array[33631] <= 16'b0000_0000_0000_0000;
array[33632] <= 16'b0000_0000_0000_0000;
array[33633] <= 16'b0000_0000_0000_0000;
array[33634] <= 16'b0000_0000_0000_0000;
array[33635] <= 16'b0000_0000_0000_0000;
array[33636] <= 16'b0000_0000_0000_0000;
array[33637] <= 16'b0000_0000_0000_0000;
array[33638] <= 16'b0000_0000_0000_0000;
array[33639] <= 16'b0000_0000_0000_0000;
array[33640] <= 16'b0000_0000_0000_0000;
array[33641] <= 16'b0000_0000_0000_0000;
array[33642] <= 16'b0000_0000_0000_0000;
array[33643] <= 16'b0000_0000_0000_0000;
array[33644] <= 16'b0000_0000_0000_0000;
array[33645] <= 16'b0000_0000_0000_0000;
array[33646] <= 16'b0000_0000_0000_0000;
array[33647] <= 16'b0000_0000_0000_0000;
array[33648] <= 16'b0000_0000_0000_0000;
array[33649] <= 16'b0000_0000_0000_0000;
array[33650] <= 16'b0000_0000_0000_0000;
array[33651] <= 16'b0000_0000_0000_0000;
array[33652] <= 16'b0000_0000_0000_0000;
array[33653] <= 16'b0000_0000_0000_0000;
array[33654] <= 16'b0000_0000_0000_0000;
array[33655] <= 16'b0000_0000_0000_0000;
array[33656] <= 16'b0000_0000_0000_0000;
array[33657] <= 16'b0000_0000_0000_0000;
array[33658] <= 16'b0000_0000_0000_0000;
array[33659] <= 16'b0000_0000_0000_0000;
array[33660] <= 16'b0000_0000_0000_0000;
array[33661] <= 16'b0000_0000_0000_0000;
array[33662] <= 16'b0000_0000_0000_0000;
array[33663] <= 16'b0000_0000_0000_0000;
array[33664] <= 16'b0000_0000_0000_0000;
array[33665] <= 16'b0000_0000_0000_0000;
array[33666] <= 16'b0000_0000_0000_0000;
array[33667] <= 16'b0000_0000_0000_0000;
array[33668] <= 16'b0000_0000_0000_0000;
array[33669] <= 16'b0000_0000_0000_0000;
array[33670] <= 16'b0000_0000_0000_0000;
array[33671] <= 16'b0000_0000_0000_0000;
array[33672] <= 16'b0000_0000_0000_0000;
array[33673] <= 16'b0000_0000_0000_0000;
array[33674] <= 16'b0000_0000_0000_0000;
array[33675] <= 16'b0000_0000_0000_0000;
array[33676] <= 16'b0000_0000_0000_0000;
array[33677] <= 16'b0000_0000_0000_0000;
array[33678] <= 16'b0000_0000_0000_0000;
array[33679] <= 16'b0000_0000_0000_0000;
array[33680] <= 16'b0000_0000_0000_0000;
array[33681] <= 16'b0000_0000_0000_0000;
array[33682] <= 16'b0000_0000_0000_0000;
array[33683] <= 16'b0000_0000_0000_0000;
array[33684] <= 16'b0000_0000_0000_0000;
array[33685] <= 16'b0000_0000_0000_0000;
array[33686] <= 16'b0000_0000_0000_0000;
array[33687] <= 16'b0000_0000_0000_0000;
array[33688] <= 16'b0000_0000_0000_0000;
array[33689] <= 16'b0000_0000_0000_0000;
array[33690] <= 16'b0000_0000_0000_0000;
array[33691] <= 16'b0000_0000_0000_0000;
array[33692] <= 16'b0000_0000_0000_0000;
array[33693] <= 16'b0000_0000_0000_0000;
array[33694] <= 16'b0000_0000_0000_0000;
array[33695] <= 16'b0000_0000_0000_0000;
array[33696] <= 16'b0000_0000_0000_0000;
array[33697] <= 16'b0000_0000_0000_0000;
array[33698] <= 16'b0000_0000_0000_0000;
array[33699] <= 16'b0000_0000_0000_0000;
array[33700] <= 16'b0000_0000_0000_0000;
array[33701] <= 16'b0000_0000_0000_0000;
array[33702] <= 16'b0000_0000_0000_0000;
array[33703] <= 16'b0000_0000_0000_0000;
array[33704] <= 16'b0000_0000_0000_0000;
array[33705] <= 16'b0000_0000_0000_0000;
array[33706] <= 16'b0000_0000_0000_0000;
array[33707] <= 16'b0000_0000_0000_0000;
array[33708] <= 16'b0000_0000_0000_0000;
array[33709] <= 16'b0000_0000_0000_0000;
array[33710] <= 16'b0000_0000_0000_0000;
array[33711] <= 16'b0000_0000_0000_0000;
array[33712] <= 16'b0000_0000_0000_0000;
array[33713] <= 16'b0000_0000_0000_0000;
array[33714] <= 16'b0000_0000_0000_0000;
array[33715] <= 16'b0000_0000_0000_0000;
array[33716] <= 16'b0000_0000_0000_0000;
array[33717] <= 16'b0000_0000_0000_0000;
array[33718] <= 16'b0000_0000_0000_0000;
array[33719] <= 16'b0000_0000_0000_0000;
array[33720] <= 16'b0000_0000_0000_0000;
array[33721] <= 16'b0000_0000_0000_0000;
array[33722] <= 16'b0000_0000_0000_0000;
array[33723] <= 16'b0000_0000_0000_0000;
array[33724] <= 16'b0000_0000_0000_0000;
array[33725] <= 16'b0000_0000_0000_0000;
array[33726] <= 16'b0000_0000_0000_0000;
array[33727] <= 16'b0000_0000_0000_0000;
array[33728] <= 16'b0000_0000_0000_0000;
array[33729] <= 16'b0000_0000_0000_0000;
array[33730] <= 16'b0000_0000_0000_0000;
array[33731] <= 16'b0000_0000_0000_0000;
array[33732] <= 16'b0000_0000_0000_0000;
array[33733] <= 16'b0000_0000_0000_0000;
array[33734] <= 16'b0000_0000_0000_0000;
array[33735] <= 16'b0000_0000_0000_0000;
array[33736] <= 16'b0000_0000_0000_0000;
array[33737] <= 16'b0000_0000_0000_0000;
array[33738] <= 16'b0000_0000_0000_0000;
array[33739] <= 16'b0000_0000_0000_0000;
array[33740] <= 16'b0000_0000_0000_0000;
array[33741] <= 16'b0000_0000_0000_0000;
array[33742] <= 16'b0000_0000_0000_0000;
array[33743] <= 16'b0000_0000_0000_0000;
array[33744] <= 16'b0000_0000_0000_0000;
array[33745] <= 16'b0000_0000_0000_0000;
array[33746] <= 16'b0000_0000_0000_0000;
array[33747] <= 16'b0000_0000_0000_0000;
array[33748] <= 16'b0000_0000_0000_0000;
array[33749] <= 16'b0000_0000_0000_0000;
array[33750] <= 16'b0000_0000_0000_0000;
array[33751] <= 16'b0000_0000_0000_0000;
array[33752] <= 16'b0000_0000_0000_0000;
array[33753] <= 16'b0000_0000_0000_0000;
array[33754] <= 16'b0000_0000_0000_0000;
array[33755] <= 16'b0000_0000_0000_0000;
array[33756] <= 16'b0000_0000_0000_0000;
array[33757] <= 16'b0000_0000_0000_0000;
array[33758] <= 16'b0000_0000_0000_0000;
array[33759] <= 16'b0000_0000_0000_0000;
array[33760] <= 16'b0000_0000_0000_0000;
array[33761] <= 16'b0000_0000_0000_0000;
array[33762] <= 16'b0000_0000_0000_0000;
array[33763] <= 16'b0000_0000_0000_0000;
array[33764] <= 16'b0000_0000_0000_0000;
array[33765] <= 16'b0000_0000_0000_0000;
array[33766] <= 16'b0000_0000_0000_0000;
array[33767] <= 16'b0000_0000_0000_0000;
array[33768] <= 16'b0000_0000_0000_0000;
array[33769] <= 16'b0000_0000_0000_0000;
array[33770] <= 16'b0000_0000_0000_0000;
array[33771] <= 16'b0000_0000_0000_0000;
array[33772] <= 16'b0000_0000_0000_0000;
array[33773] <= 16'b0000_0000_0000_0000;
array[33774] <= 16'b0000_0000_0000_0000;
array[33775] <= 16'b0000_0000_0000_0000;
array[33776] <= 16'b0000_0000_0000_0000;
array[33777] <= 16'b0000_0000_0000_0000;
array[33778] <= 16'b0000_0000_0000_0000;
array[33779] <= 16'b0000_0000_0000_0000;
array[33780] <= 16'b0000_0000_0000_0000;
array[33781] <= 16'b0000_0000_0000_0000;
array[33782] <= 16'b0000_0000_0000_0000;
array[33783] <= 16'b0000_0000_0000_0000;
array[33784] <= 16'b0000_0000_0000_0000;
array[33785] <= 16'b0000_0000_0000_0000;
array[33786] <= 16'b0000_0000_0000_0000;
array[33787] <= 16'b0000_0000_0000_0000;
array[33788] <= 16'b0000_0000_0000_0000;
array[33789] <= 16'b0000_0000_0000_0000;
array[33790] <= 16'b0000_0000_0000_0000;
array[33791] <= 16'b0000_0000_0000_0000;
array[33792] <= 16'b0000_0000_0000_0000;
array[33793] <= 16'b0000_0000_0000_0000;
array[33794] <= 16'b0000_0000_0000_0000;
array[33795] <= 16'b0000_0000_0000_0000;
array[33796] <= 16'b0000_0000_0000_0000;
array[33797] <= 16'b0000_0000_0000_0000;
array[33798] <= 16'b0000_0000_0000_0000;
array[33799] <= 16'b0000_0000_0000_0000;
array[33800] <= 16'b0000_0000_0000_0000;
array[33801] <= 16'b0000_0000_0000_0000;
array[33802] <= 16'b0000_0000_0000_0000;
array[33803] <= 16'b0000_0000_0000_0000;
array[33804] <= 16'b0000_0000_0000_0000;
array[33805] <= 16'b0000_0000_0000_0000;
array[33806] <= 16'b0000_0000_0000_0000;
array[33807] <= 16'b0000_0000_0000_0000;
array[33808] <= 16'b0000_0000_0000_0000;
array[33809] <= 16'b0000_0000_0000_0000;
array[33810] <= 16'b0000_0000_0000_0000;
array[33811] <= 16'b0000_0000_0000_0000;
array[33812] <= 16'b0000_0000_0000_0000;
array[33813] <= 16'b0000_0000_0000_0000;
array[33814] <= 16'b0000_0000_0000_0000;
array[33815] <= 16'b0000_0000_0000_0000;
array[33816] <= 16'b0000_0000_0000_0000;
array[33817] <= 16'b0000_0000_0000_0000;
array[33818] <= 16'b0000_0000_0000_0000;
array[33819] <= 16'b0000_0000_0000_0000;
array[33820] <= 16'b0000_0000_0000_0000;
array[33821] <= 16'b0000_0000_0000_0000;
array[33822] <= 16'b0000_0000_0000_0000;
array[33823] <= 16'b0000_0000_0000_0000;
array[33824] <= 16'b0000_0000_0000_0000;
array[33825] <= 16'b0000_0000_0000_0000;
array[33826] <= 16'b0000_0000_0000_0000;
array[33827] <= 16'b0000_0000_0000_0000;
array[33828] <= 16'b0000_0000_0000_0000;
array[33829] <= 16'b0000_0000_0000_0000;
array[33830] <= 16'b0000_0000_0000_0000;
array[33831] <= 16'b0000_0000_0000_0000;
array[33832] <= 16'b0000_0000_0000_0000;
array[33833] <= 16'b0000_0000_0000_0000;
array[33834] <= 16'b0000_0000_0000_0000;
array[33835] <= 16'b0000_0000_0000_0000;
array[33836] <= 16'b0000_0000_0000_0000;
array[33837] <= 16'b0000_0000_0000_0000;
array[33838] <= 16'b0000_0000_0000_0000;
array[33839] <= 16'b0000_0000_0000_0000;
array[33840] <= 16'b0000_0000_0000_0000;
array[33841] <= 16'b0000_0000_0000_0000;
array[33842] <= 16'b0000_0000_0000_0000;
array[33843] <= 16'b0000_0000_0000_0000;
array[33844] <= 16'b0000_0000_0000_0000;
array[33845] <= 16'b0000_0000_0000_0000;
array[33846] <= 16'b0000_0000_0000_0000;
array[33847] <= 16'b0000_0000_0000_0000;
array[33848] <= 16'b0000_0000_0000_0000;
array[33849] <= 16'b0000_0000_0000_0000;
array[33850] <= 16'b0000_0000_0000_0000;
array[33851] <= 16'b0000_0000_0000_0000;
array[33852] <= 16'b0000_0000_0000_0000;
array[33853] <= 16'b0000_0000_0000_0000;
array[33854] <= 16'b0000_0000_0000_0000;
array[33855] <= 16'b0000_0000_0000_0000;
array[33856] <= 16'b0000_0000_0000_0000;
array[33857] <= 16'b0000_0000_0000_0000;
array[33858] <= 16'b0000_0000_0000_0000;
array[33859] <= 16'b0000_0000_0000_0000;
array[33860] <= 16'b0000_0000_0000_0000;
array[33861] <= 16'b0000_0000_0000_0000;
array[33862] <= 16'b0000_0000_0000_0000;
array[33863] <= 16'b0000_0000_0000_0000;
array[33864] <= 16'b0000_0000_0000_0000;
array[33865] <= 16'b0000_0000_0000_0000;
array[33866] <= 16'b0000_0000_0000_0000;
array[33867] <= 16'b0000_0000_0000_0000;
array[33868] <= 16'b0000_0000_0000_0000;
array[33869] <= 16'b0000_0000_0000_0000;
array[33870] <= 16'b0000_0000_0000_0000;
array[33871] <= 16'b0000_0000_0000_0000;
array[33872] <= 16'b0000_0000_0000_0000;
array[33873] <= 16'b0000_0000_0000_0000;
array[33874] <= 16'b0000_0000_0000_0000;
array[33875] <= 16'b0000_0000_0000_0000;
array[33876] <= 16'b0000_0000_0000_0000;
array[33877] <= 16'b0000_0000_0000_0000;
array[33878] <= 16'b0000_0000_0000_0000;
array[33879] <= 16'b0000_0000_0000_0000;
array[33880] <= 16'b0000_0000_0000_0000;
array[33881] <= 16'b0000_0000_0000_0000;
array[33882] <= 16'b0000_0000_0000_0000;
array[33883] <= 16'b0000_0000_0000_0000;
array[33884] <= 16'b0000_0000_0000_0000;
array[33885] <= 16'b0000_0000_0000_0000;
array[33886] <= 16'b0000_0000_0000_0000;
array[33887] <= 16'b0000_0000_0000_0000;
array[33888] <= 16'b0000_0000_0000_0000;
array[33889] <= 16'b0000_0000_0000_0000;
array[33890] <= 16'b0000_0000_0000_0000;
array[33891] <= 16'b0000_0000_0000_0000;
array[33892] <= 16'b0000_0000_0000_0000;
array[33893] <= 16'b0000_0000_0000_0000;
array[33894] <= 16'b0000_0000_0000_0000;
array[33895] <= 16'b0000_0000_0000_0000;
array[33896] <= 16'b0000_0000_0000_0000;
array[33897] <= 16'b0000_0000_0000_0000;
array[33898] <= 16'b0000_0000_0000_0000;
array[33899] <= 16'b0000_0000_0000_0000;
array[33900] <= 16'b0000_0000_0000_0000;
array[33901] <= 16'b0000_0000_0000_0000;
array[33902] <= 16'b0000_0000_0000_0000;
array[33903] <= 16'b0000_0000_0000_0000;
array[33904] <= 16'b0000_0000_0000_0000;
array[33905] <= 16'b0000_0000_0000_0000;
array[33906] <= 16'b0000_0000_0000_0000;
array[33907] <= 16'b0000_0000_0000_0000;
array[33908] <= 16'b0000_0000_0000_0000;
array[33909] <= 16'b0000_0000_0000_0000;
array[33910] <= 16'b0000_0000_0000_0000;
array[33911] <= 16'b0000_0000_0000_0000;
array[33912] <= 16'b0000_0000_0000_0000;
array[33913] <= 16'b0000_0000_0000_0000;
array[33914] <= 16'b0000_0000_0000_0000;
array[33915] <= 16'b0000_0000_0000_0000;
array[33916] <= 16'b0000_0000_0000_0000;
array[33917] <= 16'b0000_0000_0000_0000;
array[33918] <= 16'b0000_0000_0000_0000;
array[33919] <= 16'b0000_0000_0000_0000;
array[33920] <= 16'b0000_0000_0000_0000;
array[33921] <= 16'b0000_0000_0000_0000;
array[33922] <= 16'b0000_0000_0000_0000;
array[33923] <= 16'b0000_0000_0000_0000;
array[33924] <= 16'b0000_0000_0000_0000;
array[33925] <= 16'b0000_0000_0000_0000;
array[33926] <= 16'b0000_0000_0000_0000;
array[33927] <= 16'b0000_0000_0000_0000;
array[33928] <= 16'b0000_0000_0000_0000;
array[33929] <= 16'b0000_0000_0000_0000;
array[33930] <= 16'b0000_0000_0000_0000;
array[33931] <= 16'b0000_0000_0000_0000;
array[33932] <= 16'b0000_0000_0000_0000;
array[33933] <= 16'b0000_0000_0000_0000;
array[33934] <= 16'b0000_0000_0000_0000;
array[33935] <= 16'b0000_0000_0000_0000;
array[33936] <= 16'b0000_0000_0000_0000;
array[33937] <= 16'b0000_0000_0000_0000;
array[33938] <= 16'b0000_0000_0000_0000;
array[33939] <= 16'b0000_0000_0000_0000;
array[33940] <= 16'b0000_0000_0000_0000;
array[33941] <= 16'b0000_0000_0000_0000;
array[33942] <= 16'b0000_0000_0000_0000;
array[33943] <= 16'b0000_0000_0000_0000;
array[33944] <= 16'b0000_0000_0000_0000;
array[33945] <= 16'b0000_0000_0000_0000;
array[33946] <= 16'b0000_0000_0000_0000;
array[33947] <= 16'b0000_0000_0000_0000;
array[33948] <= 16'b0000_0000_0000_0000;
array[33949] <= 16'b0000_0000_0000_0000;
array[33950] <= 16'b0000_0000_0000_0000;
array[33951] <= 16'b0000_0000_0000_0000;
array[33952] <= 16'b0000_0000_0000_0000;
array[33953] <= 16'b0000_0000_0000_0000;
array[33954] <= 16'b0000_0000_0000_0000;
array[33955] <= 16'b0000_0000_0000_0000;
array[33956] <= 16'b0000_0000_0000_0000;
array[33957] <= 16'b0000_0000_0000_0000;
array[33958] <= 16'b0000_0000_0000_0000;
array[33959] <= 16'b0000_0000_0000_0000;
array[33960] <= 16'b0000_0000_0000_0000;
array[33961] <= 16'b0000_0000_0000_0000;
array[33962] <= 16'b0000_0000_0000_0000;
array[33963] <= 16'b0000_0000_0000_0000;
array[33964] <= 16'b0000_0000_0000_0000;
array[33965] <= 16'b0000_0000_0000_0000;
array[33966] <= 16'b0000_0000_0000_0000;
array[33967] <= 16'b0000_0000_0000_0000;
array[33968] <= 16'b0000_0000_0000_0000;
array[33969] <= 16'b0000_0000_0000_0000;
array[33970] <= 16'b0000_0000_0000_0000;
array[33971] <= 16'b0000_0000_0000_0000;
array[33972] <= 16'b0000_0000_0000_0000;
array[33973] <= 16'b0000_0000_0000_0000;
array[33974] <= 16'b0000_0000_0000_0000;
array[33975] <= 16'b0000_0000_0000_0000;
array[33976] <= 16'b0000_0000_0000_0000;
array[33977] <= 16'b0000_0000_0000_0000;
array[33978] <= 16'b0000_0000_0000_0000;
array[33979] <= 16'b0000_0000_0000_0000;
array[33980] <= 16'b0000_0000_0000_0000;
array[33981] <= 16'b0000_0000_0000_0000;
array[33982] <= 16'b0000_0000_0000_0000;
array[33983] <= 16'b0000_0000_0000_0000;
array[33984] <= 16'b0000_0000_0000_0000;
array[33985] <= 16'b0000_0000_0000_0000;
array[33986] <= 16'b0000_0000_0000_0000;
array[33987] <= 16'b0000_0000_0000_0000;
array[33988] <= 16'b0000_0000_0000_0000;
array[33989] <= 16'b0000_0000_0000_0000;
array[33990] <= 16'b0000_0000_0000_0000;
array[33991] <= 16'b0000_0000_0000_0000;
array[33992] <= 16'b0000_0000_0000_0000;
array[33993] <= 16'b0000_0000_0000_0000;
array[33994] <= 16'b0000_0000_0000_0000;
array[33995] <= 16'b0000_0000_0000_0000;
array[33996] <= 16'b0000_0000_0000_0000;
array[33997] <= 16'b0000_0000_0000_0000;
array[33998] <= 16'b0000_0000_0000_0000;
array[33999] <= 16'b0000_0000_0000_0000;
array[34000] <= 16'b0000_0000_0000_0000;
array[34001] <= 16'b0000_0000_0000_0000;
array[34002] <= 16'b0000_0000_0000_0000;
array[34003] <= 16'b0000_0000_0000_0000;
array[34004] <= 16'b0000_0000_0000_0000;
array[34005] <= 16'b0000_0000_0000_0000;
array[34006] <= 16'b0000_0000_0000_0000;
array[34007] <= 16'b0000_0000_0000_0000;
array[34008] <= 16'b0000_0000_0000_0000;
array[34009] <= 16'b0000_0000_0000_0000;
array[34010] <= 16'b0000_0000_0000_0000;
array[34011] <= 16'b0000_0000_0000_0000;
array[34012] <= 16'b0000_0000_0000_0000;
array[34013] <= 16'b0000_0000_0000_0000;
array[34014] <= 16'b0000_0000_0000_0000;
array[34015] <= 16'b0000_0000_0000_0000;
array[34016] <= 16'b0000_0000_0000_0000;
array[34017] <= 16'b0000_0000_0000_0000;
array[34018] <= 16'b0000_0000_0000_0000;
array[34019] <= 16'b0000_0000_0000_0000;
array[34020] <= 16'b0000_0000_0000_0000;
array[34021] <= 16'b0000_0000_0000_0000;
array[34022] <= 16'b0000_0000_0000_0000;
array[34023] <= 16'b0000_0000_0000_0000;
array[34024] <= 16'b0000_0000_0000_0000;
array[34025] <= 16'b0000_0000_0000_0000;
array[34026] <= 16'b0000_0000_0000_0000;
array[34027] <= 16'b0000_0000_0000_0000;
array[34028] <= 16'b0000_0000_0000_0000;
array[34029] <= 16'b0000_0000_0000_0000;
array[34030] <= 16'b0000_0000_0000_0000;
array[34031] <= 16'b0000_0000_0000_0000;
array[34032] <= 16'b0000_0000_0000_0000;
array[34033] <= 16'b0000_0000_0000_0000;
array[34034] <= 16'b0000_0000_0000_0000;
array[34035] <= 16'b0000_0000_0000_0000;
array[34036] <= 16'b0000_0000_0000_0000;
array[34037] <= 16'b0000_0000_0000_0000;
array[34038] <= 16'b0000_0000_0000_0000;
array[34039] <= 16'b0000_0000_0000_0000;
array[34040] <= 16'b0000_0000_0000_0000;
array[34041] <= 16'b0000_0000_0000_0000;
array[34042] <= 16'b0000_0000_0000_0000;
array[34043] <= 16'b0000_0000_0000_0000;
array[34044] <= 16'b0000_0000_0000_0000;
array[34045] <= 16'b0000_0000_0000_0000;
array[34046] <= 16'b0000_0000_0000_0000;
array[34047] <= 16'b0000_0000_0000_0000;
array[34048] <= 16'b0000_0000_0000_0000;
array[34049] <= 16'b0000_0000_0000_0000;
array[34050] <= 16'b0000_0000_0000_0000;
array[34051] <= 16'b0000_0000_0000_0000;
array[34052] <= 16'b0000_0000_0000_0000;
array[34053] <= 16'b0000_0000_0000_0000;
array[34054] <= 16'b0000_0000_0000_0000;
array[34055] <= 16'b0000_0000_0000_0000;
array[34056] <= 16'b0000_0000_0000_0000;
array[34057] <= 16'b0000_0000_0000_0000;
array[34058] <= 16'b0000_0000_0000_0000;
array[34059] <= 16'b0000_0000_0000_0000;
array[34060] <= 16'b0000_0000_0000_0000;
array[34061] <= 16'b0000_0000_0000_0000;
array[34062] <= 16'b0000_0000_0000_0000;
array[34063] <= 16'b0000_0000_0000_0000;
array[34064] <= 16'b0000_0000_0000_0000;
array[34065] <= 16'b0000_0000_0000_0000;
array[34066] <= 16'b0000_0000_0000_0000;
array[34067] <= 16'b0000_0000_0000_0000;
array[34068] <= 16'b0000_0000_0000_0000;
array[34069] <= 16'b0000_0000_0000_0000;
array[34070] <= 16'b0000_0000_0000_0000;
array[34071] <= 16'b0000_0000_0000_0000;
array[34072] <= 16'b0000_0000_0000_0000;
array[34073] <= 16'b0000_0000_0000_0000;
array[34074] <= 16'b0000_0000_0000_0000;
array[34075] <= 16'b0000_0000_0000_0000;
array[34076] <= 16'b0000_0000_0000_0000;
array[34077] <= 16'b0000_0000_0000_0000;
array[34078] <= 16'b0000_0000_0000_0000;
array[34079] <= 16'b0000_0000_0000_0000;
array[34080] <= 16'b0000_0000_0000_0000;
array[34081] <= 16'b0000_0000_0000_0000;
array[34082] <= 16'b0000_0000_0000_0000;
array[34083] <= 16'b0000_0000_0000_0000;
array[34084] <= 16'b0000_0000_0000_0000;
array[34085] <= 16'b0000_0000_0000_0000;
array[34086] <= 16'b0000_0000_0000_0000;
array[34087] <= 16'b0000_0000_0000_0000;
array[34088] <= 16'b0000_0000_0000_0000;
array[34089] <= 16'b0000_0000_0000_0000;
array[34090] <= 16'b0000_0000_0000_0000;
array[34091] <= 16'b0000_0000_0000_0000;
array[34092] <= 16'b0000_0000_0000_0000;
array[34093] <= 16'b0000_0000_0000_0000;
array[34094] <= 16'b0000_0000_0000_0000;
array[34095] <= 16'b0000_0000_0000_0000;
array[34096] <= 16'b0000_0000_0000_0000;
array[34097] <= 16'b0000_0000_0000_0000;
array[34098] <= 16'b0000_0000_0000_0000;
array[34099] <= 16'b0000_0000_0000_0000;
array[34100] <= 16'b0000_0000_0000_0000;
array[34101] <= 16'b0000_0000_0000_0000;
array[34102] <= 16'b0000_0000_0000_0000;
array[34103] <= 16'b0000_0000_0000_0000;
array[34104] <= 16'b0000_0000_0000_0000;
array[34105] <= 16'b0000_0000_0000_0000;
array[34106] <= 16'b0000_0000_0000_0000;
array[34107] <= 16'b0000_0000_0000_0000;
array[34108] <= 16'b0000_0000_0000_0000;
array[34109] <= 16'b0000_0000_0000_0000;
array[34110] <= 16'b0000_0000_0000_0000;
array[34111] <= 16'b0000_0000_0000_0000;
array[34112] <= 16'b0000_0000_0000_0000;
array[34113] <= 16'b0000_0000_0000_0000;
array[34114] <= 16'b0000_0000_0000_0000;
array[34115] <= 16'b0000_0000_0000_0000;
array[34116] <= 16'b0000_0000_0000_0000;
array[34117] <= 16'b0000_0000_0000_0000;
array[34118] <= 16'b0000_0000_0000_0000;
array[34119] <= 16'b0000_0000_0000_0000;
array[34120] <= 16'b0000_0000_0000_0000;
array[34121] <= 16'b0000_0000_0000_0000;
array[34122] <= 16'b0000_0000_0000_0000;
array[34123] <= 16'b0000_0000_0000_0000;
array[34124] <= 16'b0000_0000_0000_0000;
array[34125] <= 16'b0000_0000_0000_0000;
array[34126] <= 16'b0000_0000_0000_0000;
array[34127] <= 16'b0000_0000_0000_0000;
array[34128] <= 16'b0000_0000_0000_0000;
array[34129] <= 16'b0000_0000_0000_0000;
array[34130] <= 16'b0000_0000_0000_0000;
array[34131] <= 16'b0000_0000_0000_0000;
array[34132] <= 16'b0000_0000_0000_0000;
array[34133] <= 16'b0000_0000_0000_0000;
array[34134] <= 16'b0000_0000_0000_0000;
array[34135] <= 16'b0000_0000_0000_0000;
array[34136] <= 16'b0000_0000_0000_0000;
array[34137] <= 16'b0000_0000_0000_0000;
array[34138] <= 16'b0000_0000_0000_0000;
array[34139] <= 16'b0000_0000_0000_0000;
array[34140] <= 16'b0000_0000_0000_0000;
array[34141] <= 16'b0000_0000_0000_0000;
array[34142] <= 16'b0000_0000_0000_0000;
array[34143] <= 16'b0000_0000_0000_0000;
array[34144] <= 16'b0000_0000_0000_0000;
array[34145] <= 16'b0000_0000_0000_0000;
array[34146] <= 16'b0000_0000_0000_0000;
array[34147] <= 16'b0000_0000_0000_0000;
array[34148] <= 16'b0000_0000_0000_0000;
array[34149] <= 16'b0000_0000_0000_0000;
array[34150] <= 16'b0000_0000_0000_0000;
array[34151] <= 16'b0000_0000_0000_0000;
array[34152] <= 16'b0000_0000_0000_0000;
array[34153] <= 16'b0000_0000_0000_0000;
array[34154] <= 16'b0000_0000_0000_0000;
array[34155] <= 16'b0000_0000_0000_0000;
array[34156] <= 16'b0000_0000_0000_0000;
array[34157] <= 16'b0000_0000_0000_0000;
array[34158] <= 16'b0000_0000_0000_0000;
array[34159] <= 16'b0000_0000_0000_0000;
array[34160] <= 16'b0000_0000_0000_0000;
array[34161] <= 16'b0000_0000_0000_0000;
array[34162] <= 16'b0000_0000_0000_0000;
array[34163] <= 16'b0000_0000_0000_0000;
array[34164] <= 16'b0000_0000_0000_0000;
array[34165] <= 16'b0000_0000_0000_0000;
array[34166] <= 16'b0000_0000_0000_0000;
array[34167] <= 16'b0000_0000_0000_0000;
array[34168] <= 16'b0000_0000_0000_0000;
array[34169] <= 16'b0000_0000_0000_0000;
array[34170] <= 16'b0000_0000_0000_0000;
array[34171] <= 16'b0000_0000_0000_0000;
array[34172] <= 16'b0000_0000_0000_0000;
array[34173] <= 16'b0000_0000_0000_0000;
array[34174] <= 16'b0000_0000_0000_0000;
array[34175] <= 16'b0000_0000_0000_0000;
array[34176] <= 16'b0000_0000_0000_0000;
array[34177] <= 16'b0000_0000_0000_0000;
array[34178] <= 16'b0000_0000_0000_0000;
array[34179] <= 16'b0000_0000_0000_0000;
array[34180] <= 16'b0000_0000_0000_0000;
array[34181] <= 16'b0000_0000_0000_0000;
array[34182] <= 16'b0000_0000_0000_0000;
array[34183] <= 16'b0000_0000_0000_0000;
array[34184] <= 16'b0000_0000_0000_0000;
array[34185] <= 16'b0000_0000_0000_0000;
array[34186] <= 16'b0000_0000_0000_0000;
array[34187] <= 16'b0000_0000_0000_0000;
array[34188] <= 16'b0000_0000_0000_0000;
array[34189] <= 16'b0000_0000_0000_0000;
array[34190] <= 16'b0000_0000_0000_0000;
array[34191] <= 16'b0000_0000_0000_0000;
array[34192] <= 16'b0000_0000_0000_0000;
array[34193] <= 16'b0000_0000_0000_0000;
array[34194] <= 16'b0000_0000_0000_0000;
array[34195] <= 16'b0000_0000_0000_0000;
array[34196] <= 16'b0000_0000_0000_0000;
array[34197] <= 16'b0000_0000_0000_0000;
array[34198] <= 16'b0000_0000_0000_0000;
array[34199] <= 16'b0000_0000_0000_0000;
array[34200] <= 16'b0000_0000_0000_0000;
array[34201] <= 16'b0000_0000_0000_0000;
array[34202] <= 16'b0000_0000_0000_0000;
array[34203] <= 16'b0000_0000_0000_0000;
array[34204] <= 16'b0000_0000_0000_0000;
array[34205] <= 16'b0000_0000_0000_0000;
array[34206] <= 16'b0000_0000_0000_0000;
array[34207] <= 16'b0000_0000_0000_0000;
array[34208] <= 16'b0000_0000_0000_0000;
array[34209] <= 16'b0000_0000_0000_0000;
array[34210] <= 16'b0000_0000_0000_0000;
array[34211] <= 16'b0000_0000_0000_0000;
array[34212] <= 16'b0000_0000_0000_0000;
array[34213] <= 16'b0000_0000_0000_0000;
array[34214] <= 16'b0000_0000_0000_0000;
array[34215] <= 16'b0000_0000_0000_0000;
array[34216] <= 16'b0000_0000_0000_0000;
array[34217] <= 16'b0000_0000_0000_0000;
array[34218] <= 16'b0000_0000_0000_0000;
array[34219] <= 16'b0000_0000_0000_0000;
array[34220] <= 16'b0000_0000_0000_0000;
array[34221] <= 16'b0000_0000_0000_0000;
array[34222] <= 16'b0000_0000_0000_0000;
array[34223] <= 16'b0000_0000_0000_0000;
array[34224] <= 16'b0000_0000_0000_0000;
array[34225] <= 16'b0000_0000_0000_0000;
array[34226] <= 16'b0000_0000_0000_0000;
array[34227] <= 16'b0000_0000_0000_0000;
array[34228] <= 16'b0000_0000_0000_0000;
array[34229] <= 16'b0000_0000_0000_0000;
array[34230] <= 16'b0000_0000_0000_0000;
array[34231] <= 16'b0000_0000_0000_0000;
array[34232] <= 16'b0000_0000_0000_0000;
array[34233] <= 16'b0000_0000_0000_0000;
array[34234] <= 16'b0000_0000_0000_0000;
array[34235] <= 16'b0000_0000_0000_0000;
array[34236] <= 16'b0000_0000_0000_0000;
array[34237] <= 16'b0000_0000_0000_0000;
array[34238] <= 16'b0000_0000_0000_0000;
array[34239] <= 16'b0000_0000_0000_0000;
array[34240] <= 16'b0000_0000_0000_0000;
array[34241] <= 16'b0000_0000_0000_0000;
array[34242] <= 16'b0000_0000_0000_0000;
array[34243] <= 16'b0000_0000_0000_0000;
array[34244] <= 16'b0000_0000_0000_0000;
array[34245] <= 16'b0000_0000_0000_0000;
array[34246] <= 16'b0000_0000_0000_0000;
array[34247] <= 16'b0000_0000_0000_0000;
array[34248] <= 16'b0000_0000_0000_0000;
array[34249] <= 16'b0000_0000_0000_0000;
array[34250] <= 16'b0000_0000_0000_0000;
array[34251] <= 16'b0000_0000_0000_0000;
array[34252] <= 16'b0000_0000_0000_0000;
array[34253] <= 16'b0000_0000_0000_0000;
array[34254] <= 16'b0000_0000_0000_0000;
array[34255] <= 16'b0000_0000_0000_0000;
array[34256] <= 16'b0000_0000_0000_0000;
array[34257] <= 16'b0000_0000_0000_0000;
array[34258] <= 16'b0000_0000_0000_0000;
array[34259] <= 16'b0000_0000_0000_0000;
array[34260] <= 16'b0000_0000_0000_0000;
array[34261] <= 16'b0000_0000_0000_0000;
array[34262] <= 16'b0000_0000_0000_0000;
array[34263] <= 16'b0000_0000_0000_0000;
array[34264] <= 16'b0000_0000_0000_0000;
array[34265] <= 16'b0000_0000_0000_0000;
array[34266] <= 16'b0000_0000_0000_0000;
array[34267] <= 16'b0000_0000_0000_0000;
array[34268] <= 16'b0000_0000_0000_0000;
array[34269] <= 16'b0000_0000_0000_0000;
array[34270] <= 16'b0000_0000_0000_0000;
array[34271] <= 16'b0000_0000_0000_0000;
array[34272] <= 16'b0000_0000_0000_0000;
array[34273] <= 16'b0000_0000_0000_0000;
array[34274] <= 16'b0000_0000_0000_0000;
array[34275] <= 16'b0000_0000_0000_0000;
array[34276] <= 16'b0000_0000_0000_0000;
array[34277] <= 16'b0000_0000_0000_0000;
array[34278] <= 16'b0000_0000_0000_0000;
array[34279] <= 16'b0000_0000_0000_0000;
array[34280] <= 16'b0000_0000_0000_0000;
array[34281] <= 16'b0000_0000_0000_0000;
array[34282] <= 16'b0000_0000_0000_0000;
array[34283] <= 16'b0000_0000_0000_0000;
array[34284] <= 16'b0000_0000_0000_0000;
array[34285] <= 16'b0000_0000_0000_0000;
array[34286] <= 16'b0000_0000_0000_0000;
array[34287] <= 16'b0000_0000_0000_0000;
array[34288] <= 16'b0000_0000_0000_0000;
array[34289] <= 16'b0000_0000_0000_0000;
array[34290] <= 16'b0000_0000_0000_0000;
array[34291] <= 16'b0000_0000_0000_0000;
array[34292] <= 16'b0000_0000_0000_0000;
array[34293] <= 16'b0000_0000_0000_0000;
array[34294] <= 16'b0000_0000_0000_0000;
array[34295] <= 16'b0000_0000_0000_0000;
array[34296] <= 16'b0000_0000_0000_0000;
array[34297] <= 16'b0000_0000_0000_0000;
array[34298] <= 16'b0000_0000_0000_0000;
array[34299] <= 16'b0000_0000_0000_0000;
array[34300] <= 16'b0000_0000_0000_0000;
array[34301] <= 16'b0000_0000_0000_0000;
array[34302] <= 16'b0000_0000_0000_0000;
array[34303] <= 16'b0000_0000_0000_0000;
array[34304] <= 16'b0000_0000_0000_0000;
array[34305] <= 16'b0000_0000_0000_0000;
array[34306] <= 16'b0000_0000_0000_0000;
array[34307] <= 16'b0000_0000_0000_0000;
array[34308] <= 16'b0000_0000_0000_0000;
array[34309] <= 16'b0000_0000_0000_0000;
array[34310] <= 16'b0000_0000_0000_0000;
array[34311] <= 16'b0000_0000_0000_0000;
array[34312] <= 16'b0000_0000_0000_0000;
array[34313] <= 16'b0000_0000_0000_0000;
array[34314] <= 16'b0000_0000_0000_0000;
array[34315] <= 16'b0000_0000_0000_0000;
array[34316] <= 16'b0000_0000_0000_0000;
array[34317] <= 16'b0000_0000_0000_0000;
array[34318] <= 16'b0000_0000_0000_0000;
array[34319] <= 16'b0000_0000_0000_0000;
array[34320] <= 16'b0000_0000_0000_0000;
array[34321] <= 16'b0000_0000_0000_0000;
array[34322] <= 16'b0000_0000_0000_0000;
array[34323] <= 16'b0000_0000_0000_0000;
array[34324] <= 16'b0000_0000_0000_0000;
array[34325] <= 16'b0000_0000_0000_0000;
array[34326] <= 16'b0000_0000_0000_0000;
array[34327] <= 16'b0000_0000_0000_0000;
array[34328] <= 16'b0000_0000_0000_0000;
array[34329] <= 16'b0000_0000_0000_0000;
array[34330] <= 16'b0000_0000_0000_0000;
array[34331] <= 16'b0000_0000_0000_0000;
array[34332] <= 16'b0000_0000_0000_0000;
array[34333] <= 16'b0000_0000_0000_0000;
array[34334] <= 16'b0000_0000_0000_0000;
array[34335] <= 16'b0000_0000_0000_0000;
array[34336] <= 16'b0000_0000_0000_0000;
array[34337] <= 16'b0000_0000_0000_0000;
array[34338] <= 16'b0000_0000_0000_0000;
array[34339] <= 16'b0000_0000_0000_0000;
array[34340] <= 16'b0000_0000_0000_0000;
array[34341] <= 16'b0000_0000_0000_0000;
array[34342] <= 16'b0000_0000_0000_0000;
array[34343] <= 16'b0000_0000_0000_0000;
array[34344] <= 16'b0000_0000_0000_0000;
array[34345] <= 16'b0000_0000_0000_0000;
array[34346] <= 16'b0000_0000_0000_0000;
array[34347] <= 16'b0000_0000_0000_0000;
array[34348] <= 16'b0000_0000_0000_0000;
array[34349] <= 16'b0000_0000_0000_0000;
array[34350] <= 16'b0000_0000_0000_0000;
array[34351] <= 16'b0000_0000_0000_0000;
array[34352] <= 16'b0000_0000_0000_0000;
array[34353] <= 16'b0000_0000_0000_0000;
array[34354] <= 16'b0000_0000_0000_0000;
array[34355] <= 16'b0000_0000_0000_0000;
array[34356] <= 16'b0000_0000_0000_0000;
array[34357] <= 16'b0000_0000_0000_0000;
array[34358] <= 16'b0000_0000_0000_0000;
array[34359] <= 16'b0000_0000_0000_0000;
array[34360] <= 16'b0000_0000_0000_0000;
array[34361] <= 16'b0000_0000_0000_0000;
array[34362] <= 16'b0000_0000_0000_0000;
array[34363] <= 16'b0000_0000_0000_0000;
array[34364] <= 16'b0000_0000_0000_0000;
array[34365] <= 16'b0000_0000_0000_0000;
array[34366] <= 16'b0000_0000_0000_0000;
array[34367] <= 16'b0000_0000_0000_0000;
array[34368] <= 16'b0000_0000_0000_0000;
array[34369] <= 16'b0000_0000_0000_0000;
array[34370] <= 16'b0000_0000_0000_0000;
array[34371] <= 16'b0000_0000_0000_0000;
array[34372] <= 16'b0000_0000_0000_0000;
array[34373] <= 16'b0000_0000_0000_0000;
array[34374] <= 16'b0000_0000_0000_0000;
array[34375] <= 16'b0000_0000_0000_0000;
array[34376] <= 16'b0000_0000_0000_0000;
array[34377] <= 16'b0000_0000_0000_0000;
array[34378] <= 16'b0000_0000_0000_0000;
array[34379] <= 16'b0000_0000_0000_0000;
array[34380] <= 16'b0000_0000_0000_0000;
array[34381] <= 16'b0000_0000_0000_0000;
array[34382] <= 16'b0000_0000_0000_0000;
array[34383] <= 16'b0000_0000_0000_0000;
array[34384] <= 16'b0000_0000_0000_0000;
array[34385] <= 16'b0000_0000_0000_0000;
array[34386] <= 16'b0000_0000_0000_0000;
array[34387] <= 16'b0000_0000_0000_0000;
array[34388] <= 16'b0000_0000_0000_0000;
array[34389] <= 16'b0000_0000_0000_0000;
array[34390] <= 16'b0000_0000_0000_0000;
array[34391] <= 16'b0000_0000_0000_0000;
array[34392] <= 16'b0000_0000_0000_0000;
array[34393] <= 16'b0000_0000_0000_0000;
array[34394] <= 16'b0000_0000_0000_0000;
array[34395] <= 16'b0000_0000_0000_0000;
array[34396] <= 16'b0000_0000_0000_0000;
array[34397] <= 16'b0000_0000_0000_0000;
array[34398] <= 16'b0000_0000_0000_0000;
array[34399] <= 16'b0000_0000_0000_0000;
array[34400] <= 16'b0000_0000_0000_0000;
array[34401] <= 16'b0000_0000_0000_0000;
array[34402] <= 16'b0000_0000_0000_0000;
array[34403] <= 16'b0000_0000_0000_0000;
array[34404] <= 16'b0000_0000_0000_0000;
array[34405] <= 16'b0000_0000_0000_0000;
array[34406] <= 16'b0000_0000_0000_0000;
array[34407] <= 16'b0000_0000_0000_0000;
array[34408] <= 16'b0000_0000_0000_0000;
array[34409] <= 16'b0000_0000_0000_0000;
array[34410] <= 16'b0000_0000_0000_0000;
array[34411] <= 16'b0000_0000_0000_0000;
array[34412] <= 16'b0000_0000_0000_0000;
array[34413] <= 16'b0000_0000_0000_0000;
array[34414] <= 16'b0000_0000_0000_0000;
array[34415] <= 16'b0000_0000_0000_0000;
array[34416] <= 16'b0000_0000_0000_0000;
array[34417] <= 16'b0000_0000_0000_0000;
array[34418] <= 16'b0000_0000_0000_0000;
array[34419] <= 16'b0000_0000_0000_0000;
array[34420] <= 16'b0000_0000_0000_0000;
array[34421] <= 16'b0000_0000_0000_0000;
array[34422] <= 16'b0000_0000_0000_0000;
array[34423] <= 16'b0000_0000_0000_0000;
array[34424] <= 16'b0000_0000_0000_0000;
array[34425] <= 16'b0000_0000_0000_0000;
array[34426] <= 16'b0000_0000_0000_0000;
array[34427] <= 16'b0000_0000_0000_0000;
array[34428] <= 16'b0000_0000_0000_0000;
array[34429] <= 16'b0000_0000_0000_0000;
array[34430] <= 16'b0000_0000_0000_0000;
array[34431] <= 16'b0000_0000_0000_0000;
array[34432] <= 16'b0000_0000_0000_0000;
array[34433] <= 16'b0000_0000_0000_0000;
array[34434] <= 16'b0000_0000_0000_0000;
array[34435] <= 16'b0000_0000_0000_0000;
array[34436] <= 16'b0000_0000_0000_0000;
array[34437] <= 16'b0000_0000_0000_0000;
array[34438] <= 16'b0000_0000_0000_0000;
array[34439] <= 16'b0000_0000_0000_0000;
array[34440] <= 16'b0000_0000_0000_0000;
array[34441] <= 16'b0000_0000_0000_0000;
array[34442] <= 16'b0000_0000_0000_0000;
array[34443] <= 16'b0000_0000_0000_0000;
array[34444] <= 16'b0000_0000_0000_0000;
array[34445] <= 16'b0000_0000_0000_0000;
array[34446] <= 16'b0000_0000_0000_0000;
array[34447] <= 16'b0000_0000_0000_0000;
array[34448] <= 16'b0000_0000_0000_0000;
array[34449] <= 16'b0000_0000_0000_0000;
array[34450] <= 16'b0000_0000_0000_0000;
array[34451] <= 16'b0000_0000_0000_0000;
array[34452] <= 16'b0000_0000_0000_0000;
array[34453] <= 16'b0000_0000_0000_0000;
array[34454] <= 16'b0000_0000_0000_0000;
array[34455] <= 16'b0000_0000_0000_0000;
array[34456] <= 16'b0000_0000_0000_0000;
array[34457] <= 16'b0000_0000_0000_0000;
array[34458] <= 16'b0000_0000_0000_0000;
array[34459] <= 16'b0000_0000_0000_0000;
array[34460] <= 16'b0000_0000_0000_0000;
array[34461] <= 16'b0000_0000_0000_0000;
array[34462] <= 16'b0000_0000_0000_0000;
array[34463] <= 16'b0000_0000_0000_0000;
array[34464] <= 16'b0000_0000_0000_0000;
array[34465] <= 16'b0000_0000_0000_0000;
array[34466] <= 16'b0000_0000_0000_0000;
array[34467] <= 16'b0000_0000_0000_0000;
array[34468] <= 16'b0000_0000_0000_0000;
array[34469] <= 16'b0000_0000_0000_0000;
array[34470] <= 16'b0000_0000_0000_0000;
array[34471] <= 16'b0000_0000_0000_0000;
array[34472] <= 16'b0000_0000_0000_0000;
array[34473] <= 16'b0000_0000_0000_0000;
array[34474] <= 16'b0000_0000_0000_0000;
array[34475] <= 16'b0000_0000_0000_0000;
array[34476] <= 16'b0000_0000_0000_0000;
array[34477] <= 16'b0000_0000_0000_0000;
array[34478] <= 16'b0000_0000_0000_0000;
array[34479] <= 16'b0000_0000_0000_0000;
array[34480] <= 16'b0000_0000_0000_0000;
array[34481] <= 16'b0000_0000_0000_0000;
array[34482] <= 16'b0000_0000_0000_0000;
array[34483] <= 16'b0000_0000_0000_0000;
array[34484] <= 16'b0000_0000_0000_0000;
array[34485] <= 16'b0000_0000_0000_0000;
array[34486] <= 16'b0000_0000_0000_0000;
array[34487] <= 16'b0000_0000_0000_0000;
array[34488] <= 16'b0000_0000_0000_0000;
array[34489] <= 16'b0000_0000_0000_0000;
array[34490] <= 16'b0000_0000_0000_0000;
array[34491] <= 16'b0000_0000_0000_0000;
array[34492] <= 16'b0000_0000_0000_0000;
array[34493] <= 16'b0000_0000_0000_0000;
array[34494] <= 16'b0000_0000_0000_0000;
array[34495] <= 16'b0000_0000_0000_0000;
array[34496] <= 16'b0000_0000_0000_0000;
array[34497] <= 16'b0000_0000_0000_0000;
array[34498] <= 16'b0000_0000_0000_0000;
array[34499] <= 16'b0000_0000_0000_0000;
array[34500] <= 16'b0000_0000_0000_0000;
array[34501] <= 16'b0000_0000_0000_0000;
array[34502] <= 16'b0000_0000_0000_0000;
array[34503] <= 16'b0000_0000_0000_0000;
array[34504] <= 16'b0000_0000_0000_0000;
array[34505] <= 16'b0000_0000_0000_0000;
array[34506] <= 16'b0000_0000_0000_0000;
array[34507] <= 16'b0000_0000_0000_0000;
array[34508] <= 16'b0000_0000_0000_0000;
array[34509] <= 16'b0000_0000_0000_0000;
array[34510] <= 16'b0000_0000_0000_0000;
array[34511] <= 16'b0000_0000_0000_0000;
array[34512] <= 16'b0000_0000_0000_0000;
array[34513] <= 16'b0000_0000_0000_0000;
array[34514] <= 16'b0000_0000_0000_0000;
array[34515] <= 16'b0000_0000_0000_0000;
array[34516] <= 16'b0000_0000_0000_0000;
array[34517] <= 16'b0000_0000_0000_0000;
array[34518] <= 16'b0000_0000_0000_0000;
array[34519] <= 16'b0000_0000_0000_0000;
array[34520] <= 16'b0000_0000_0000_0000;
array[34521] <= 16'b0000_0000_0000_0000;
array[34522] <= 16'b0000_0000_0000_0000;
array[34523] <= 16'b0000_0000_0000_0000;
array[34524] <= 16'b0000_0000_0000_0000;
array[34525] <= 16'b0000_0000_0000_0000;
array[34526] <= 16'b0000_0000_0000_0000;
array[34527] <= 16'b0000_0000_0000_0000;
array[34528] <= 16'b0000_0000_0000_0000;
array[34529] <= 16'b0000_0000_0000_0000;
array[34530] <= 16'b0000_0000_0000_0000;
array[34531] <= 16'b0000_0000_0000_0000;
array[34532] <= 16'b0000_0000_0000_0000;
array[34533] <= 16'b0000_0000_0000_0000;
array[34534] <= 16'b0000_0000_0000_0000;
array[34535] <= 16'b0000_0000_0000_0000;
array[34536] <= 16'b0000_0000_0000_0000;
array[34537] <= 16'b0000_0000_0000_0000;
array[34538] <= 16'b0000_0000_0000_0000;
array[34539] <= 16'b0000_0000_0000_0000;
array[34540] <= 16'b0000_0000_0000_0000;
array[34541] <= 16'b0000_0000_0000_0000;
array[34542] <= 16'b0000_0000_0000_0000;
array[34543] <= 16'b0000_0000_0000_0000;
array[34544] <= 16'b0000_0000_0000_0000;
array[34545] <= 16'b0000_0000_0000_0000;
array[34546] <= 16'b0000_0000_0000_0000;
array[34547] <= 16'b0000_0000_0000_0000;
array[34548] <= 16'b0000_0000_0000_0000;
array[34549] <= 16'b0000_0000_0000_0000;
array[34550] <= 16'b0000_0000_0000_0000;
array[34551] <= 16'b0000_0000_0000_0000;
array[34552] <= 16'b0000_0000_0000_0000;
array[34553] <= 16'b0000_0000_0000_0000;
array[34554] <= 16'b0000_0000_0000_0000;
array[34555] <= 16'b0000_0000_0000_0000;
array[34556] <= 16'b0000_0000_0000_0000;
array[34557] <= 16'b0000_0000_0000_0000;
array[34558] <= 16'b0000_0000_0000_0000;
array[34559] <= 16'b0000_0000_0000_0000;
array[34560] <= 16'b0000_0000_0000_0000;
array[34561] <= 16'b0000_0000_0000_0000;
array[34562] <= 16'b0000_0000_0000_0000;
array[34563] <= 16'b0000_0000_0000_0000;
array[34564] <= 16'b0000_0000_0000_0000;
array[34565] <= 16'b0000_0000_0000_0000;
array[34566] <= 16'b0000_0000_0000_0000;
array[34567] <= 16'b0000_0000_0000_0000;
array[34568] <= 16'b0000_0000_0000_0000;
array[34569] <= 16'b0000_0000_0000_0000;
array[34570] <= 16'b0000_0000_0000_0000;
array[34571] <= 16'b0000_0000_0000_0000;
array[34572] <= 16'b0000_0000_0000_0000;
array[34573] <= 16'b0000_0000_0000_0000;
array[34574] <= 16'b0000_0000_0000_0000;
array[34575] <= 16'b0000_0000_0000_0000;
array[34576] <= 16'b0000_0000_0000_0000;
array[34577] <= 16'b0000_0000_0000_0000;
array[34578] <= 16'b0000_0000_0000_0000;
array[34579] <= 16'b0000_0000_0000_0000;
array[34580] <= 16'b0000_0000_0000_0000;
array[34581] <= 16'b0000_0000_0000_0000;
array[34582] <= 16'b0000_0000_0000_0000;
array[34583] <= 16'b0000_0000_0000_0000;
array[34584] <= 16'b0000_0000_0000_0000;
array[34585] <= 16'b0000_0000_0000_0000;
array[34586] <= 16'b0000_0000_0000_0000;
array[34587] <= 16'b0000_0000_0000_0000;
array[34588] <= 16'b0000_0000_0000_0000;
array[34589] <= 16'b0000_0000_0000_0000;
array[34590] <= 16'b0000_0000_0000_0000;
array[34591] <= 16'b0000_0000_0000_0000;
array[34592] <= 16'b0000_0000_0000_0000;
array[34593] <= 16'b0000_0000_0000_0000;
array[34594] <= 16'b0000_0000_0000_0000;
array[34595] <= 16'b0000_0000_0000_0000;
array[34596] <= 16'b0000_0000_0000_0000;
array[34597] <= 16'b0000_0000_0000_0000;
array[34598] <= 16'b0000_0000_0000_0000;
array[34599] <= 16'b0000_0000_0000_0000;
array[34600] <= 16'b0000_0000_0000_0000;
array[34601] <= 16'b0000_0000_0000_0000;
array[34602] <= 16'b0000_0000_0000_0000;
array[34603] <= 16'b0000_0000_0000_0000;
array[34604] <= 16'b0000_0000_0000_0000;
array[34605] <= 16'b0000_0000_0000_0000;
array[34606] <= 16'b0000_0000_0000_0000;
array[34607] <= 16'b0000_0000_0000_0000;
array[34608] <= 16'b0000_0000_0000_0000;
array[34609] <= 16'b0000_0000_0000_0000;
array[34610] <= 16'b0000_0000_0000_0000;
array[34611] <= 16'b0000_0000_0000_0000;
array[34612] <= 16'b0000_0000_0000_0000;
array[34613] <= 16'b0000_0000_0000_0000;
array[34614] <= 16'b0000_0000_0000_0000;
array[34615] <= 16'b0000_0000_0000_0000;
array[34616] <= 16'b0000_0000_0000_0000;
array[34617] <= 16'b0000_0000_0000_0000;
array[34618] <= 16'b0000_0000_0000_0000;
array[34619] <= 16'b0000_0000_0000_0000;
array[34620] <= 16'b0000_0000_0000_0000;
array[34621] <= 16'b0000_0000_0000_0000;
array[34622] <= 16'b0000_0000_0000_0000;
array[34623] <= 16'b0000_0000_0000_0000;
array[34624] <= 16'b0000_0000_0000_0000;
array[34625] <= 16'b0000_0000_0000_0000;
array[34626] <= 16'b0000_0000_0000_0000;
array[34627] <= 16'b0000_0000_0000_0000;
array[34628] <= 16'b0000_0000_0000_0000;
array[34629] <= 16'b0000_0000_0000_0000;
array[34630] <= 16'b0000_0000_0000_0000;
array[34631] <= 16'b0000_0000_0000_0000;
array[34632] <= 16'b0000_0000_0000_0000;
array[34633] <= 16'b0000_0000_0000_0000;
array[34634] <= 16'b0000_0000_0000_0000;
array[34635] <= 16'b0000_0000_0000_0000;
array[34636] <= 16'b0000_0000_0000_0000;
array[34637] <= 16'b0000_0000_0000_0000;
array[34638] <= 16'b0000_0000_0000_0000;
array[34639] <= 16'b0000_0000_0000_0000;
array[34640] <= 16'b0000_0000_0000_0000;
array[34641] <= 16'b0000_0000_0000_0000;
array[34642] <= 16'b0000_0000_0000_0000;
array[34643] <= 16'b0000_0000_0000_0000;
array[34644] <= 16'b0000_0000_0000_0000;
array[34645] <= 16'b0000_0000_0000_0000;
array[34646] <= 16'b0000_0000_0000_0000;
array[34647] <= 16'b0000_0000_0000_0000;
array[34648] <= 16'b0000_0000_0000_0000;
array[34649] <= 16'b0000_0000_0000_0000;
array[34650] <= 16'b0000_0000_0000_0000;
array[34651] <= 16'b0000_0000_0000_0000;
array[34652] <= 16'b0000_0000_0000_0000;
array[34653] <= 16'b0000_0000_0000_0000;
array[34654] <= 16'b0000_0000_0000_0000;
array[34655] <= 16'b0000_0000_0000_0000;
array[34656] <= 16'b0000_0000_0000_0000;
array[34657] <= 16'b0000_0000_0000_0000;
array[34658] <= 16'b0000_0000_0000_0000;
array[34659] <= 16'b0000_0000_0000_0000;
array[34660] <= 16'b0000_0000_0000_0000;
array[34661] <= 16'b0000_0000_0000_0000;
array[34662] <= 16'b0000_0000_0000_0000;
array[34663] <= 16'b0000_0000_0000_0000;
array[34664] <= 16'b0000_0000_0000_0000;
array[34665] <= 16'b0000_0000_0000_0000;
array[34666] <= 16'b0000_0000_0000_0000;
array[34667] <= 16'b0000_0000_0000_0000;
array[34668] <= 16'b0000_0000_0000_0000;
array[34669] <= 16'b0000_0000_0000_0000;
array[34670] <= 16'b0000_0000_0000_0000;
array[34671] <= 16'b0000_0000_0000_0000;
array[34672] <= 16'b0000_0000_0000_0000;
array[34673] <= 16'b0000_0000_0000_0000;
array[34674] <= 16'b0000_0000_0000_0000;
array[34675] <= 16'b0000_0000_0000_0000;
array[34676] <= 16'b0000_0000_0000_0000;
array[34677] <= 16'b0000_0000_0000_0000;
array[34678] <= 16'b0000_0000_0000_0000;
array[34679] <= 16'b0000_0000_0000_0000;
array[34680] <= 16'b0000_0000_0000_0000;
array[34681] <= 16'b0000_0000_0000_0000;
array[34682] <= 16'b0000_0000_0000_0000;
array[34683] <= 16'b0000_0000_0000_0000;
array[34684] <= 16'b0000_0000_0000_0000;
array[34685] <= 16'b0000_0000_0000_0000;
array[34686] <= 16'b0000_0000_0000_0000;
array[34687] <= 16'b0000_0000_0000_0000;
array[34688] <= 16'b0000_0000_0000_0000;
array[34689] <= 16'b0000_0000_0000_0000;
array[34690] <= 16'b0000_0000_0000_0000;
array[34691] <= 16'b0000_0000_0000_0000;
array[34692] <= 16'b0000_0000_0000_0000;
array[34693] <= 16'b0000_0000_0000_0000;
array[34694] <= 16'b0000_0000_0000_0000;
array[34695] <= 16'b0000_0000_0000_0000;
array[34696] <= 16'b0000_0000_0000_0000;
array[34697] <= 16'b0000_0000_0000_0000;
array[34698] <= 16'b0000_0000_0000_0000;
array[34699] <= 16'b0000_0000_0000_0000;
array[34700] <= 16'b0000_0000_0000_0000;
array[34701] <= 16'b0000_0000_0000_0000;
array[34702] <= 16'b0000_0000_0000_0000;
array[34703] <= 16'b0000_0000_0000_0000;
array[34704] <= 16'b0000_0000_0000_0000;
array[34705] <= 16'b0000_0000_0000_0000;
array[34706] <= 16'b0000_0000_0000_0000;
array[34707] <= 16'b0000_0000_0000_0000;
array[34708] <= 16'b0000_0000_0000_0000;
array[34709] <= 16'b0000_0000_0000_0000;
array[34710] <= 16'b0000_0000_0000_0000;
array[34711] <= 16'b0000_0000_0000_0000;
array[34712] <= 16'b0000_0000_0000_0000;
array[34713] <= 16'b0000_0000_0000_0000;
array[34714] <= 16'b0000_0000_0000_0000;
array[34715] <= 16'b0000_0000_0000_0000;
array[34716] <= 16'b0000_0000_0000_0000;
array[34717] <= 16'b0000_0000_0000_0000;
array[34718] <= 16'b0000_0000_0000_0000;
array[34719] <= 16'b0000_0000_0000_0000;
array[34720] <= 16'b0000_0000_0000_0000;
array[34721] <= 16'b0000_0000_0000_0000;
array[34722] <= 16'b0000_0000_0000_0000;
array[34723] <= 16'b0000_0000_0000_0000;
array[34724] <= 16'b0000_0000_0000_0000;
array[34725] <= 16'b0000_0000_0000_0000;
array[34726] <= 16'b0000_0000_0000_0000;
array[34727] <= 16'b0000_0000_0000_0000;
array[34728] <= 16'b0000_0000_0000_0000;
array[34729] <= 16'b0000_0000_0000_0000;
array[34730] <= 16'b0000_0000_0000_0000;
array[34731] <= 16'b0000_0000_0000_0000;
array[34732] <= 16'b0000_0000_0000_0000;
array[34733] <= 16'b0000_0000_0000_0000;
array[34734] <= 16'b0000_0000_0000_0000;
array[34735] <= 16'b0000_0000_0000_0000;
array[34736] <= 16'b0000_0000_0000_0000;
array[34737] <= 16'b0000_0000_0000_0000;
array[34738] <= 16'b0000_0000_0000_0000;
array[34739] <= 16'b0000_0000_0000_0000;
array[34740] <= 16'b0000_0000_0000_0000;
array[34741] <= 16'b0000_0000_0000_0000;
array[34742] <= 16'b0000_0000_0000_0000;
array[34743] <= 16'b0000_0000_0000_0000;
array[34744] <= 16'b0000_0000_0000_0000;
array[34745] <= 16'b0000_0000_0000_0000;
array[34746] <= 16'b0000_0000_0000_0000;
array[34747] <= 16'b0000_0000_0000_0000;
array[34748] <= 16'b0000_0000_0000_0000;
array[34749] <= 16'b0000_0000_0000_0000;
array[34750] <= 16'b0000_0000_0000_0000;
array[34751] <= 16'b0000_0000_0000_0000;
array[34752] <= 16'b0000_0000_0000_0000;
array[34753] <= 16'b0000_0000_0000_0000;
array[34754] <= 16'b0000_0000_0000_0000;
array[34755] <= 16'b0000_0000_0000_0000;
array[34756] <= 16'b0000_0000_0000_0000;
array[34757] <= 16'b0000_0000_0000_0000;
array[34758] <= 16'b0000_0000_0000_0000;
array[34759] <= 16'b0000_0000_0000_0000;
array[34760] <= 16'b0000_0000_0000_0000;
array[34761] <= 16'b0000_0000_0000_0000;
array[34762] <= 16'b0000_0000_0000_0000;
array[34763] <= 16'b0000_0000_0000_0000;
array[34764] <= 16'b0000_0000_0000_0000;
array[34765] <= 16'b0000_0000_0000_0000;
array[34766] <= 16'b0000_0000_0000_0000;
array[34767] <= 16'b0000_0000_0000_0000;
array[34768] <= 16'b0000_0000_0000_0000;
array[34769] <= 16'b0000_0000_0000_0000;
array[34770] <= 16'b0000_0000_0000_0000;
array[34771] <= 16'b0000_0000_0000_0000;
array[34772] <= 16'b0000_0000_0000_0000;
array[34773] <= 16'b0000_0000_0000_0000;
array[34774] <= 16'b0000_0000_0000_0000;
array[34775] <= 16'b0000_0000_0000_0000;
array[34776] <= 16'b0000_0000_0000_0000;
array[34777] <= 16'b0000_0000_0000_0000;
array[34778] <= 16'b0000_0000_0000_0000;
array[34779] <= 16'b0000_0000_0000_0000;
array[34780] <= 16'b0000_0000_0000_0000;
array[34781] <= 16'b0000_0000_0000_0000;
array[34782] <= 16'b0000_0000_0000_0000;
array[34783] <= 16'b0000_0000_0000_0000;
array[34784] <= 16'b0000_0000_0000_0000;
array[34785] <= 16'b0000_0000_0000_0000;
array[34786] <= 16'b0000_0000_0000_0000;
array[34787] <= 16'b0000_0000_0000_0000;
array[34788] <= 16'b0000_0000_0000_0000;
array[34789] <= 16'b0000_0000_0000_0000;
array[34790] <= 16'b0000_0000_0000_0000;
array[34791] <= 16'b0000_0000_0000_0000;
array[34792] <= 16'b0000_0000_0000_0000;
array[34793] <= 16'b0000_0000_0000_0000;
array[34794] <= 16'b0000_0000_0000_0000;
array[34795] <= 16'b0000_0000_0000_0000;
array[34796] <= 16'b0000_0000_0000_0000;
array[34797] <= 16'b0000_0000_0000_0000;
array[34798] <= 16'b0000_0000_0000_0000;
array[34799] <= 16'b0000_0000_0000_0000;
array[34800] <= 16'b0000_0000_0000_0000;
array[34801] <= 16'b0000_0000_0000_0000;
array[34802] <= 16'b0000_0000_0000_0000;
array[34803] <= 16'b0000_0000_0000_0000;
array[34804] <= 16'b0000_0000_0000_0000;
array[34805] <= 16'b0000_0000_0000_0000;
array[34806] <= 16'b0000_0000_0000_0000;
array[34807] <= 16'b0000_0000_0000_0000;
array[34808] <= 16'b0000_0000_0000_0000;
array[34809] <= 16'b0000_0000_0000_0000;
array[34810] <= 16'b0000_0000_0000_0000;
array[34811] <= 16'b0000_0000_0000_0000;
array[34812] <= 16'b0000_0000_0000_0000;
array[34813] <= 16'b0000_0000_0000_0000;
array[34814] <= 16'b0000_0000_0000_0000;
array[34815] <= 16'b0000_0000_0000_0000;
array[34816] <= 16'b0000_0000_0000_0000;
array[34817] <= 16'b0000_0000_0000_0000;
array[34818] <= 16'b0000_0000_0000_0000;
array[34819] <= 16'b0000_0000_0000_0000;
array[34820] <= 16'b0000_0000_0000_0000;
array[34821] <= 16'b0000_0000_0000_0000;
array[34822] <= 16'b0000_0000_0000_0000;
array[34823] <= 16'b0000_0000_0000_0000;
array[34824] <= 16'b0000_0000_0000_0000;
array[34825] <= 16'b0000_0000_0000_0000;
array[34826] <= 16'b0000_0000_0000_0000;
array[34827] <= 16'b0000_0000_0000_0000;
array[34828] <= 16'b0000_0000_0000_0000;
array[34829] <= 16'b0000_0000_0000_0000;
array[34830] <= 16'b0000_0000_0000_0000;
array[34831] <= 16'b0000_0000_0000_0000;
array[34832] <= 16'b0000_0000_0000_0000;
array[34833] <= 16'b0000_0000_0000_0000;
array[34834] <= 16'b0000_0000_0000_0000;
array[34835] <= 16'b0000_0000_0000_0000;
array[34836] <= 16'b0000_0000_0000_0000;
array[34837] <= 16'b0000_0000_0000_0000;
array[34838] <= 16'b0000_0000_0000_0000;
array[34839] <= 16'b0000_0000_0000_0000;
array[34840] <= 16'b0000_0000_0000_0000;
array[34841] <= 16'b0000_0000_0000_0000;
array[34842] <= 16'b0000_0000_0000_0000;
array[34843] <= 16'b0000_0000_0000_0000;
array[34844] <= 16'b0000_0000_0000_0000;
array[34845] <= 16'b0000_0000_0000_0000;
array[34846] <= 16'b0000_0000_0000_0000;
array[34847] <= 16'b0000_0000_0000_0000;
array[34848] <= 16'b0000_0000_0000_0000;
array[34849] <= 16'b0000_0000_0000_0000;
array[34850] <= 16'b0000_0000_0000_0000;
array[34851] <= 16'b0000_0000_0000_0000;
array[34852] <= 16'b0000_0000_0000_0000;
array[34853] <= 16'b0000_0000_0000_0000;
array[34854] <= 16'b0000_0000_0000_0000;
array[34855] <= 16'b0000_0000_0000_0000;
array[34856] <= 16'b0000_0000_0000_0000;
array[34857] <= 16'b0000_0000_0000_0000;
array[34858] <= 16'b0000_0000_0000_0000;
array[34859] <= 16'b0000_0000_0000_0000;
array[34860] <= 16'b0000_0000_0000_0000;
array[34861] <= 16'b0000_0000_0000_0000;
array[34862] <= 16'b0000_0000_0000_0000;
array[34863] <= 16'b0000_0000_0000_0000;
array[34864] <= 16'b0000_0000_0000_0000;
array[34865] <= 16'b0000_0000_0000_0000;
array[34866] <= 16'b0000_0000_0000_0000;
array[34867] <= 16'b0000_0000_0000_0000;
array[34868] <= 16'b0000_0000_0000_0000;
array[34869] <= 16'b0000_0000_0000_0000;
array[34870] <= 16'b0000_0000_0000_0000;
array[34871] <= 16'b0000_0000_0000_0000;
array[34872] <= 16'b0000_0000_0000_0000;
array[34873] <= 16'b0000_0000_0000_0000;
array[34874] <= 16'b0000_0000_0000_0000;
array[34875] <= 16'b0000_0000_0000_0000;
array[34876] <= 16'b0000_0000_0000_0000;
array[34877] <= 16'b0000_0000_0000_0000;
array[34878] <= 16'b0000_0000_0000_0000;
array[34879] <= 16'b0000_0000_0000_0000;
array[34880] <= 16'b0000_0000_0000_0000;
array[34881] <= 16'b0000_0000_0000_0000;
array[34882] <= 16'b0000_0000_0000_0000;
array[34883] <= 16'b0000_0000_0000_0000;
array[34884] <= 16'b0000_0000_0000_0000;
array[34885] <= 16'b0000_0000_0000_0000;
array[34886] <= 16'b0000_0000_0000_0000;
array[34887] <= 16'b0000_0000_0000_0000;
array[34888] <= 16'b0000_0000_0000_0000;
array[34889] <= 16'b0000_0000_0000_0000;
array[34890] <= 16'b0000_0000_0000_0000;
array[34891] <= 16'b0000_0000_0000_0000;
array[34892] <= 16'b0000_0000_0000_0000;
array[34893] <= 16'b0000_0000_0000_0000;
array[34894] <= 16'b0000_0000_0000_0000;
array[34895] <= 16'b0000_0000_0000_0000;
array[34896] <= 16'b0000_0000_0000_0000;
array[34897] <= 16'b0000_0000_0000_0000;
array[34898] <= 16'b0000_0000_0000_0000;
array[34899] <= 16'b0000_0000_0000_0000;
array[34900] <= 16'b0000_0000_0000_0000;
array[34901] <= 16'b0000_0000_0000_0000;
array[34902] <= 16'b0000_0000_0000_0000;
array[34903] <= 16'b0000_0000_0000_0000;
array[34904] <= 16'b0000_0000_0000_0000;
array[34905] <= 16'b0000_0000_0000_0000;
array[34906] <= 16'b0000_0000_0000_0000;
array[34907] <= 16'b0000_0000_0000_0000;
array[34908] <= 16'b0000_0000_0000_0000;
array[34909] <= 16'b0000_0000_0000_0000;
array[34910] <= 16'b0000_0000_0000_0000;
array[34911] <= 16'b0000_0000_0000_0000;
array[34912] <= 16'b0000_0000_0000_0000;
array[34913] <= 16'b0000_0000_0000_0000;
array[34914] <= 16'b0000_0000_0000_0000;
array[34915] <= 16'b0000_0000_0000_0000;
array[34916] <= 16'b0000_0000_0000_0000;
array[34917] <= 16'b0000_0000_0000_0000;
array[34918] <= 16'b0000_0000_0000_0000;
array[34919] <= 16'b0000_0000_0000_0000;
array[34920] <= 16'b0000_0000_0000_0000;
array[34921] <= 16'b0000_0000_0000_0000;
array[34922] <= 16'b0000_0000_0000_0000;
array[34923] <= 16'b0000_0000_0000_0000;
array[34924] <= 16'b0000_0000_0000_0000;
array[34925] <= 16'b0000_0000_0000_0000;
array[34926] <= 16'b0000_0000_0000_0000;
array[34927] <= 16'b0000_0000_0000_0000;
array[34928] <= 16'b0000_0000_0000_0000;
array[34929] <= 16'b0000_0000_0000_0000;
array[34930] <= 16'b0000_0000_0000_0000;
array[34931] <= 16'b0000_0000_0000_0000;
array[34932] <= 16'b0000_0000_0000_0000;
array[34933] <= 16'b0000_0000_0000_0000;
array[34934] <= 16'b0000_0000_0000_0000;
array[34935] <= 16'b0000_0000_0000_0000;
array[34936] <= 16'b0000_0000_0000_0000;
array[34937] <= 16'b0000_0000_0000_0000;
array[34938] <= 16'b0000_0000_0000_0000;
array[34939] <= 16'b0000_0000_0000_0000;
array[34940] <= 16'b0000_0000_0000_0000;
array[34941] <= 16'b0000_0000_0000_0000;
array[34942] <= 16'b0000_0000_0000_0000;
array[34943] <= 16'b0000_0000_0000_0000;
array[34944] <= 16'b0000_0000_0000_0000;
array[34945] <= 16'b0000_0000_0000_0000;
array[34946] <= 16'b0000_0000_0000_0000;
array[34947] <= 16'b0000_0000_0000_0000;
array[34948] <= 16'b0000_0000_0000_0000;
array[34949] <= 16'b0000_0000_0000_0000;
array[34950] <= 16'b0000_0000_0000_0000;
array[34951] <= 16'b0000_0000_0000_0000;
array[34952] <= 16'b0000_0000_0000_0000;
array[34953] <= 16'b0000_0000_0000_0000;
array[34954] <= 16'b0000_0000_0000_0000;
array[34955] <= 16'b0000_0000_0000_0000;
array[34956] <= 16'b0000_0000_0000_0000;
array[34957] <= 16'b0000_0000_0000_0000;
array[34958] <= 16'b0000_0000_0000_0000;
array[34959] <= 16'b0000_0000_0000_0000;
array[34960] <= 16'b0000_0000_0000_0000;
array[34961] <= 16'b0000_0000_0000_0000;
array[34962] <= 16'b0000_0000_0000_0000;
array[34963] <= 16'b0000_0000_0000_0000;
array[34964] <= 16'b0000_0000_0000_0000;
array[34965] <= 16'b0000_0000_0000_0000;
array[34966] <= 16'b0000_0000_0000_0000;
array[34967] <= 16'b0000_0000_0000_0000;
array[34968] <= 16'b0000_0000_0000_0000;
array[34969] <= 16'b0000_0000_0000_0000;
array[34970] <= 16'b0000_0000_0000_0000;
array[34971] <= 16'b0000_0000_0000_0000;
array[34972] <= 16'b0000_0000_0000_0000;
array[34973] <= 16'b0000_0000_0000_0000;
array[34974] <= 16'b0000_0000_0000_0000;
array[34975] <= 16'b0000_0000_0000_0000;
array[34976] <= 16'b0000_0000_0000_0000;
array[34977] <= 16'b0000_0000_0000_0000;
array[34978] <= 16'b0000_0000_0000_0000;
array[34979] <= 16'b0000_0000_0000_0000;
array[34980] <= 16'b0000_0000_0000_0000;
array[34981] <= 16'b0000_0000_0000_0000;
array[34982] <= 16'b0000_0000_0000_0000;
array[34983] <= 16'b0000_0000_0000_0000;
array[34984] <= 16'b0000_0000_0000_0000;
array[34985] <= 16'b0000_0000_0000_0000;
array[34986] <= 16'b0000_0000_0000_0000;
array[34987] <= 16'b0000_0000_0000_0000;
array[34988] <= 16'b0000_0000_0000_0000;
array[34989] <= 16'b0000_0000_0000_0000;
array[34990] <= 16'b0000_0000_0000_0000;
array[34991] <= 16'b0000_0000_0000_0000;
array[34992] <= 16'b0000_0000_0000_0000;
array[34993] <= 16'b0000_0000_0000_0000;
array[34994] <= 16'b0000_0000_0000_0000;
array[34995] <= 16'b0000_0000_0000_0000;
array[34996] <= 16'b0000_0000_0000_0000;
array[34997] <= 16'b0000_0000_0000_0000;
array[34998] <= 16'b0000_0000_0000_0000;
array[34999] <= 16'b0000_0000_0000_0000;
array[35000] <= 16'b0000_0000_0000_0000;
array[35001] <= 16'b0000_0000_0000_0000;
array[35002] <= 16'b0000_0000_0000_0000;
array[35003] <= 16'b0000_0000_0000_0000;
array[35004] <= 16'b0000_0000_0000_0000;
array[35005] <= 16'b0000_0000_0000_0000;
array[35006] <= 16'b0000_0000_0000_0000;
array[35007] <= 16'b0000_0000_0000_0000;
array[35008] <= 16'b0000_0000_0000_0000;
array[35009] <= 16'b0000_0000_0000_0000;
array[35010] <= 16'b0000_0000_0000_0000;
array[35011] <= 16'b0000_0000_0000_0000;
array[35012] <= 16'b0000_0000_0000_0000;
array[35013] <= 16'b0000_0000_0000_0000;
array[35014] <= 16'b0000_0000_0000_0000;
array[35015] <= 16'b0000_0000_0000_0000;
array[35016] <= 16'b0000_0000_0000_0000;
array[35017] <= 16'b0000_0000_0000_0000;
array[35018] <= 16'b0000_0000_0000_0000;
array[35019] <= 16'b0000_0000_0000_0000;
array[35020] <= 16'b0000_0000_0000_0000;
array[35021] <= 16'b0000_0000_0000_0000;
array[35022] <= 16'b0000_0000_0000_0000;
array[35023] <= 16'b0000_0000_0000_0000;
array[35024] <= 16'b0000_0000_0000_0000;
array[35025] <= 16'b0000_0000_0000_0000;
array[35026] <= 16'b0000_0000_0000_0000;
array[35027] <= 16'b0000_0000_0000_0000;
array[35028] <= 16'b0000_0000_0000_0000;
array[35029] <= 16'b0000_0000_0000_0000;
array[35030] <= 16'b0000_0000_0000_0000;
array[35031] <= 16'b0000_0000_0000_0000;
array[35032] <= 16'b0000_0000_0000_0000;
array[35033] <= 16'b0000_0000_0000_0000;
array[35034] <= 16'b0000_0000_0000_0000;
array[35035] <= 16'b0000_0000_0000_0000;
array[35036] <= 16'b0000_0000_0000_0000;
array[35037] <= 16'b0000_0000_0000_0000;
array[35038] <= 16'b0000_0000_0000_0000;
array[35039] <= 16'b0000_0000_0000_0000;
array[35040] <= 16'b0000_0000_0000_0000;
array[35041] <= 16'b0000_0000_0000_0000;
array[35042] <= 16'b0000_0000_0000_0000;
array[35043] <= 16'b0000_0000_0000_0000;
array[35044] <= 16'b0000_0000_0000_0000;
array[35045] <= 16'b0000_0000_0000_0000;
array[35046] <= 16'b0000_0000_0000_0000;
array[35047] <= 16'b0000_0000_0000_0000;
array[35048] <= 16'b0000_0000_0000_0000;
array[35049] <= 16'b0000_0000_0000_0000;
array[35050] <= 16'b0000_0000_0000_0000;
array[35051] <= 16'b0000_0000_0000_0000;
array[35052] <= 16'b0000_0000_0000_0000;
array[35053] <= 16'b0000_0000_0000_0000;
array[35054] <= 16'b0000_0000_0000_0000;
array[35055] <= 16'b0000_0000_0000_0000;
array[35056] <= 16'b0000_0000_0000_0000;
array[35057] <= 16'b0000_0000_0000_0000;
array[35058] <= 16'b0000_0000_0000_0000;
array[35059] <= 16'b0000_0000_0000_0000;
array[35060] <= 16'b0000_0000_0000_0000;
array[35061] <= 16'b0000_0000_0000_0000;
array[35062] <= 16'b0000_0000_0000_0000;
array[35063] <= 16'b0000_0000_0000_0000;
array[35064] <= 16'b0000_0000_0000_0000;
array[35065] <= 16'b0000_0000_0000_0000;
array[35066] <= 16'b0000_0000_0000_0000;
array[35067] <= 16'b0000_0000_0000_0000;
array[35068] <= 16'b0000_0000_0000_0000;
array[35069] <= 16'b0000_0000_0000_0000;
array[35070] <= 16'b0000_0000_0000_0000;
array[35071] <= 16'b0000_0000_0000_0000;
array[35072] <= 16'b0000_0000_0000_0000;
array[35073] <= 16'b0000_0000_0000_0000;
array[35074] <= 16'b0000_0000_0000_0000;
array[35075] <= 16'b0000_0000_0000_0000;
array[35076] <= 16'b0000_0000_0000_0000;
array[35077] <= 16'b0000_0000_0000_0000;
array[35078] <= 16'b0000_0000_0000_0000;
array[35079] <= 16'b0000_0000_0000_0000;
array[35080] <= 16'b0000_0000_0000_0000;
array[35081] <= 16'b0000_0000_0000_0000;
array[35082] <= 16'b0000_0000_0000_0000;
array[35083] <= 16'b0000_0000_0000_0000;
array[35084] <= 16'b0000_0000_0000_0000;
array[35085] <= 16'b0000_0000_0000_0000;
array[35086] <= 16'b0000_0000_0000_0000;
array[35087] <= 16'b0000_0000_0000_0000;
array[35088] <= 16'b0000_0000_0000_0000;
array[35089] <= 16'b0000_0000_0000_0000;
array[35090] <= 16'b0000_0000_0000_0000;
array[35091] <= 16'b0000_0000_0000_0000;
array[35092] <= 16'b0000_0000_0000_0000;
array[35093] <= 16'b0000_0000_0000_0000;
array[35094] <= 16'b0000_0000_0000_0000;
array[35095] <= 16'b0000_0000_0000_0000;
array[35096] <= 16'b0000_0000_0000_0000;
array[35097] <= 16'b0000_0000_0000_0000;
array[35098] <= 16'b0000_0000_0000_0000;
array[35099] <= 16'b0000_0000_0000_0000;
array[35100] <= 16'b0000_0000_0000_0000;
array[35101] <= 16'b0000_0000_0000_0000;
array[35102] <= 16'b0000_0000_0000_0000;
array[35103] <= 16'b0000_0000_0000_0000;
array[35104] <= 16'b0000_0000_0000_0000;
array[35105] <= 16'b0000_0000_0000_0000;
array[35106] <= 16'b0000_0000_0000_0000;
array[35107] <= 16'b0000_0000_0000_0000;
array[35108] <= 16'b0000_0000_0000_0000;
array[35109] <= 16'b0000_0000_0000_0000;
array[35110] <= 16'b0000_0000_0000_0000;
array[35111] <= 16'b0000_0000_0000_0000;
array[35112] <= 16'b0000_0000_0000_0000;
array[35113] <= 16'b0000_0000_0000_0000;
array[35114] <= 16'b0000_0000_0000_0000;
array[35115] <= 16'b0000_0000_0000_0000;
array[35116] <= 16'b0000_0000_0000_0000;
array[35117] <= 16'b0000_0000_0000_0000;
array[35118] <= 16'b0000_0000_0000_0000;
array[35119] <= 16'b0000_0000_0000_0000;
array[35120] <= 16'b0000_0000_0000_0000;
array[35121] <= 16'b0000_0000_0000_0000;
array[35122] <= 16'b0000_0000_0000_0000;
array[35123] <= 16'b0000_0000_0000_0000;
array[35124] <= 16'b0000_0000_0000_0000;
array[35125] <= 16'b0000_0000_0000_0000;
array[35126] <= 16'b0000_0000_0000_0000;
array[35127] <= 16'b0000_0000_0000_0000;
array[35128] <= 16'b0000_0000_0000_0000;
array[35129] <= 16'b0000_0000_0000_0000;
array[35130] <= 16'b0000_0000_0000_0000;
array[35131] <= 16'b0000_0000_0000_0000;
array[35132] <= 16'b0000_0000_0000_0000;
array[35133] <= 16'b0000_0000_0000_0000;
array[35134] <= 16'b0000_0000_0000_0000;
array[35135] <= 16'b0000_0000_0000_0000;
array[35136] <= 16'b0000_0000_0000_0000;
array[35137] <= 16'b0000_0000_0000_0000;
array[35138] <= 16'b0000_0000_0000_0000;
array[35139] <= 16'b0000_0000_0000_0000;
array[35140] <= 16'b0000_0000_0000_0000;
array[35141] <= 16'b0000_0000_0000_0000;
array[35142] <= 16'b0000_0000_0000_0000;
array[35143] <= 16'b0000_0000_0000_0000;
array[35144] <= 16'b0000_0000_0000_0000;
array[35145] <= 16'b0000_0000_0000_0000;
array[35146] <= 16'b0000_0000_0000_0000;
array[35147] <= 16'b0000_0000_0000_0000;
array[35148] <= 16'b0000_0000_0000_0000;
array[35149] <= 16'b0000_0000_0000_0000;
array[35150] <= 16'b0000_0000_0000_0000;
array[35151] <= 16'b0000_0000_0000_0000;
array[35152] <= 16'b0000_0000_0000_0000;
array[35153] <= 16'b0000_0000_0000_0000;
array[35154] <= 16'b0000_0000_0000_0000;
array[35155] <= 16'b0000_0000_0000_0000;
array[35156] <= 16'b0000_0000_0000_0000;
array[35157] <= 16'b0000_0000_0000_0000;
array[35158] <= 16'b0000_0000_0000_0000;
array[35159] <= 16'b0000_0000_0000_0000;
array[35160] <= 16'b0000_0000_0000_0000;
array[35161] <= 16'b0000_0000_0000_0000;
array[35162] <= 16'b0000_0000_0000_0000;
array[35163] <= 16'b0000_0000_0000_0000;
array[35164] <= 16'b0000_0000_0000_0000;
array[35165] <= 16'b0000_0000_0000_0000;
array[35166] <= 16'b0000_0000_0000_0000;
array[35167] <= 16'b0000_0000_0000_0000;
array[35168] <= 16'b0000_0000_0000_0000;
array[35169] <= 16'b0000_0000_0000_0000;
array[35170] <= 16'b0000_0000_0000_0000;
array[35171] <= 16'b0000_0000_0000_0000;
array[35172] <= 16'b0000_0000_0000_0000;
array[35173] <= 16'b0000_0000_0000_0000;
array[35174] <= 16'b0000_0000_0000_0000;
array[35175] <= 16'b0000_0000_0000_0000;
array[35176] <= 16'b0000_0000_0000_0000;
array[35177] <= 16'b0000_0000_0000_0000;
array[35178] <= 16'b0000_0000_0000_0000;
array[35179] <= 16'b0000_0000_0000_0000;
array[35180] <= 16'b0000_0000_0000_0000;
array[35181] <= 16'b0000_0000_0000_0000;
array[35182] <= 16'b0000_0000_0000_0000;
array[35183] <= 16'b0000_0000_0000_0000;
array[35184] <= 16'b0000_0000_0000_0000;
array[35185] <= 16'b0000_0000_0000_0000;
array[35186] <= 16'b0000_0000_0000_0000;
array[35187] <= 16'b0000_0000_0000_0000;
array[35188] <= 16'b0000_0000_0000_0000;
array[35189] <= 16'b0000_0000_0000_0000;
array[35190] <= 16'b0000_0000_0000_0000;
array[35191] <= 16'b0000_0000_0000_0000;
array[35192] <= 16'b0000_0000_0000_0000;
array[35193] <= 16'b0000_0000_0000_0000;
array[35194] <= 16'b0000_0000_0000_0000;
array[35195] <= 16'b0000_0000_0000_0000;
array[35196] <= 16'b0000_0000_0000_0000;
array[35197] <= 16'b0000_0000_0000_0000;
array[35198] <= 16'b0000_0000_0000_0000;
array[35199] <= 16'b0000_0000_0000_0000;
array[35200] <= 16'b0000_0000_0000_0000;
array[35201] <= 16'b0000_0000_0000_0000;
array[35202] <= 16'b0000_0000_0000_0000;
array[35203] <= 16'b0000_0000_0000_0000;
array[35204] <= 16'b0000_0000_0000_0000;
array[35205] <= 16'b0000_0000_0000_0000;
array[35206] <= 16'b0000_0000_0000_0000;
array[35207] <= 16'b0000_0000_0000_0000;
array[35208] <= 16'b0000_0000_0000_0000;
array[35209] <= 16'b0000_0000_0000_0000;
array[35210] <= 16'b0000_0000_0000_0000;
array[35211] <= 16'b0000_0000_0000_0000;
array[35212] <= 16'b0000_0000_0000_0000;
array[35213] <= 16'b0000_0000_0000_0000;
array[35214] <= 16'b0000_0000_0000_0000;
array[35215] <= 16'b0000_0000_0000_0000;
array[35216] <= 16'b0000_0000_0000_0000;
array[35217] <= 16'b0000_0000_0000_0000;
array[35218] <= 16'b0000_0000_0000_0000;
array[35219] <= 16'b0000_0000_0000_0000;
array[35220] <= 16'b0000_0000_0000_0000;
array[35221] <= 16'b0000_0000_0000_0000;
array[35222] <= 16'b0000_0000_0000_0000;
array[35223] <= 16'b0000_0000_0000_0000;
array[35224] <= 16'b0000_0000_0000_0000;
array[35225] <= 16'b0000_0000_0000_0000;
array[35226] <= 16'b0000_0000_0000_0000;
array[35227] <= 16'b0000_0000_0000_0000;
array[35228] <= 16'b0000_0000_0000_0000;
array[35229] <= 16'b0000_0000_0000_0000;
array[35230] <= 16'b0000_0000_0000_0000;
array[35231] <= 16'b0000_0000_0000_0000;
array[35232] <= 16'b0000_0000_0000_0000;
array[35233] <= 16'b0000_0000_0000_0000;
array[35234] <= 16'b0000_0000_0000_0000;
array[35235] <= 16'b0000_0000_0000_0000;
array[35236] <= 16'b0000_0000_0000_0000;
array[35237] <= 16'b0000_0000_0000_0000;
array[35238] <= 16'b0000_0000_0000_0000;
array[35239] <= 16'b0000_0000_0000_0000;
array[35240] <= 16'b0000_0000_0000_0000;
array[35241] <= 16'b0000_0000_0000_0000;
array[35242] <= 16'b0000_0000_0000_0000;
array[35243] <= 16'b0000_0000_0000_0000;
array[35244] <= 16'b0000_0000_0000_0000;
array[35245] <= 16'b0000_0000_0000_0000;
array[35246] <= 16'b0000_0000_0000_0000;
array[35247] <= 16'b0000_0000_0000_0000;
array[35248] <= 16'b0000_0000_0000_0000;
array[35249] <= 16'b0000_0000_0000_0000;
array[35250] <= 16'b0000_0000_0000_0000;
array[35251] <= 16'b0000_0000_0000_0000;
array[35252] <= 16'b0000_0000_0000_0000;
array[35253] <= 16'b0000_0000_0000_0000;
array[35254] <= 16'b0000_0000_0000_0000;
array[35255] <= 16'b0000_0000_0000_0000;
array[35256] <= 16'b0000_0000_0000_0000;
array[35257] <= 16'b0000_0000_0000_0000;
array[35258] <= 16'b0000_0000_0000_0000;
array[35259] <= 16'b0000_0000_0000_0000;
array[35260] <= 16'b0000_0000_0000_0000;
array[35261] <= 16'b0000_0000_0000_0000;
array[35262] <= 16'b0000_0000_0000_0000;
array[35263] <= 16'b0000_0000_0000_0000;
array[35264] <= 16'b0000_0000_0000_0000;
array[35265] <= 16'b0000_0000_0000_0000;
array[35266] <= 16'b0000_0000_0000_0000;
array[35267] <= 16'b0000_0000_0000_0000;
array[35268] <= 16'b0000_0000_0000_0000;
array[35269] <= 16'b0000_0000_0000_0000;
array[35270] <= 16'b0000_0000_0000_0000;
array[35271] <= 16'b0000_0000_0000_0000;
array[35272] <= 16'b0000_0000_0000_0000;
array[35273] <= 16'b0000_0000_0000_0000;
array[35274] <= 16'b0000_0000_0000_0000;
array[35275] <= 16'b0000_0000_0000_0000;
array[35276] <= 16'b0000_0000_0000_0000;
array[35277] <= 16'b0000_0000_0000_0000;
array[35278] <= 16'b0000_0000_0000_0000;
array[35279] <= 16'b0000_0000_0000_0000;
array[35280] <= 16'b0000_0000_0000_0000;
array[35281] <= 16'b0000_0000_0000_0000;
array[35282] <= 16'b0000_0000_0000_0000;
array[35283] <= 16'b0000_0000_0000_0000;
array[35284] <= 16'b0000_0000_0000_0000;
array[35285] <= 16'b0000_0000_0000_0000;
array[35286] <= 16'b0000_0000_0000_0000;
array[35287] <= 16'b0000_0000_0000_0000;
array[35288] <= 16'b0000_0000_0000_0000;
array[35289] <= 16'b0000_0000_0000_0000;
array[35290] <= 16'b0000_0000_0000_0000;
array[35291] <= 16'b0000_0000_0000_0000;
array[35292] <= 16'b0000_0000_0000_0000;
array[35293] <= 16'b0000_0000_0000_0000;
array[35294] <= 16'b0000_0000_0000_0000;
array[35295] <= 16'b0000_0000_0000_0000;
array[35296] <= 16'b0000_0000_0000_0000;
array[35297] <= 16'b0000_0000_0000_0000;
array[35298] <= 16'b0000_0000_0000_0000;
array[35299] <= 16'b0000_0000_0000_0000;
array[35300] <= 16'b0000_0000_0000_0000;
array[35301] <= 16'b0000_0000_0000_0000;
array[35302] <= 16'b0000_0000_0000_0000;
array[35303] <= 16'b0000_0000_0000_0000;
array[35304] <= 16'b0000_0000_0000_0000;
array[35305] <= 16'b0000_0000_0000_0000;
array[35306] <= 16'b0000_0000_0000_0000;
array[35307] <= 16'b0000_0000_0000_0000;
array[35308] <= 16'b0000_0000_0000_0000;
array[35309] <= 16'b0000_0000_0000_0000;
array[35310] <= 16'b0000_0000_0000_0000;
array[35311] <= 16'b0000_0000_0000_0000;
array[35312] <= 16'b0000_0000_0000_0000;
array[35313] <= 16'b0000_0000_0000_0000;
array[35314] <= 16'b0000_0000_0000_0000;
array[35315] <= 16'b0000_0000_0000_0000;
array[35316] <= 16'b0000_0000_0000_0000;
array[35317] <= 16'b0000_0000_0000_0000;
array[35318] <= 16'b0000_0000_0000_0000;
array[35319] <= 16'b0000_0000_0000_0000;
array[35320] <= 16'b0000_0000_0000_0000;
array[35321] <= 16'b0000_0000_0000_0000;
array[35322] <= 16'b0000_0000_0000_0000;
array[35323] <= 16'b0000_0000_0000_0000;
array[35324] <= 16'b0000_0000_0000_0000;
array[35325] <= 16'b0000_0000_0000_0000;
array[35326] <= 16'b0000_0000_0000_0000;
array[35327] <= 16'b0000_0000_0000_0000;
array[35328] <= 16'b0000_0000_0000_0000;
array[35329] <= 16'b0000_0000_0000_0000;
array[35330] <= 16'b0000_0000_0000_0000;
array[35331] <= 16'b0000_0000_0000_0000;
array[35332] <= 16'b0000_0000_0000_0000;
array[35333] <= 16'b0000_0000_0000_0000;
array[35334] <= 16'b0000_0000_0000_0000;
array[35335] <= 16'b0000_0000_0000_0000;
array[35336] <= 16'b0000_0000_0000_0000;
array[35337] <= 16'b0000_0000_0000_0000;
array[35338] <= 16'b0000_0000_0000_0000;
array[35339] <= 16'b0000_0000_0000_0000;
array[35340] <= 16'b0000_0000_0000_0000;
array[35341] <= 16'b0000_0000_0000_0000;
array[35342] <= 16'b0000_0000_0000_0000;
array[35343] <= 16'b0000_0000_0000_0000;
array[35344] <= 16'b0000_0000_0000_0000;
array[35345] <= 16'b0000_0000_0000_0000;
array[35346] <= 16'b0000_0000_0000_0000;
array[35347] <= 16'b0000_0000_0000_0000;
array[35348] <= 16'b0000_0000_0000_0000;
array[35349] <= 16'b0000_0000_0000_0000;
array[35350] <= 16'b0000_0000_0000_0000;
array[35351] <= 16'b0000_0000_0000_0000;
array[35352] <= 16'b0000_0000_0000_0000;
array[35353] <= 16'b0000_0000_0000_0000;
array[35354] <= 16'b0000_0000_0000_0000;
array[35355] <= 16'b0000_0000_0000_0000;
array[35356] <= 16'b0000_0000_0000_0000;
array[35357] <= 16'b0000_0000_0000_0000;
array[35358] <= 16'b0000_0000_0000_0000;
array[35359] <= 16'b0000_0000_0000_0000;
array[35360] <= 16'b0000_0000_0000_0000;
array[35361] <= 16'b0000_0000_0000_0000;
array[35362] <= 16'b0000_0000_0000_0000;
array[35363] <= 16'b0000_0000_0000_0000;
array[35364] <= 16'b0000_0000_0000_0000;
array[35365] <= 16'b0000_0000_0000_0000;
array[35366] <= 16'b0000_0000_0000_0000;
array[35367] <= 16'b0000_0000_0000_0000;
array[35368] <= 16'b0000_0000_0000_0000;
array[35369] <= 16'b0000_0000_0000_0000;
array[35370] <= 16'b0000_0000_0000_0000;
array[35371] <= 16'b0000_0000_0000_0000;
array[35372] <= 16'b0000_0000_0000_0000;
array[35373] <= 16'b0000_0000_0000_0000;
array[35374] <= 16'b0000_0000_0000_0000;
array[35375] <= 16'b0000_0000_0000_0000;
array[35376] <= 16'b0000_0000_0000_0000;
array[35377] <= 16'b0000_0000_0000_0000;
array[35378] <= 16'b0000_0000_0000_0000;
array[35379] <= 16'b0000_0000_0000_0000;
array[35380] <= 16'b0000_0000_0000_0000;
array[35381] <= 16'b0000_0000_0000_0000;
array[35382] <= 16'b0000_0000_0000_0000;
array[35383] <= 16'b0000_0000_0000_0000;
array[35384] <= 16'b0000_0000_0000_0000;
array[35385] <= 16'b0000_0000_0000_0000;
array[35386] <= 16'b0000_0000_0000_0000;
array[35387] <= 16'b0000_0000_0000_0000;
array[35388] <= 16'b0000_0000_0000_0000;
array[35389] <= 16'b0000_0000_0000_0000;
array[35390] <= 16'b0000_0000_0000_0000;
array[35391] <= 16'b0000_0000_0000_0000;
array[35392] <= 16'b0000_0000_0000_0000;
array[35393] <= 16'b0000_0000_0000_0000;
array[35394] <= 16'b0000_0000_0000_0000;
array[35395] <= 16'b0000_0000_0000_0000;
array[35396] <= 16'b0000_0000_0000_0000;
array[35397] <= 16'b0000_0000_0000_0000;
array[35398] <= 16'b0000_0000_0000_0000;
array[35399] <= 16'b0000_0000_0000_0000;
array[35400] <= 16'b0000_0000_0000_0000;
array[35401] <= 16'b0000_0000_0000_0000;
array[35402] <= 16'b0000_0000_0000_0000;
array[35403] <= 16'b0000_0000_0000_0000;
array[35404] <= 16'b0000_0000_0000_0000;
array[35405] <= 16'b0000_0000_0000_0000;
array[35406] <= 16'b0000_0000_0000_0000;
array[35407] <= 16'b0000_0000_0000_0000;
array[35408] <= 16'b0000_0000_0000_0000;
array[35409] <= 16'b0000_0000_0000_0000;
array[35410] <= 16'b0000_0000_0000_0000;
array[35411] <= 16'b0000_0000_0000_0000;
array[35412] <= 16'b0000_0000_0000_0000;
array[35413] <= 16'b0000_0000_0000_0000;
array[35414] <= 16'b0000_0000_0000_0000;
array[35415] <= 16'b0000_0000_0000_0000;
array[35416] <= 16'b0000_0000_0000_0000;
array[35417] <= 16'b0000_0000_0000_0000;
array[35418] <= 16'b0000_0000_0000_0000;
array[35419] <= 16'b0000_0000_0000_0000;
array[35420] <= 16'b0000_0000_0000_0000;
array[35421] <= 16'b0000_0000_0000_0000;
array[35422] <= 16'b0000_0000_0000_0000;
array[35423] <= 16'b0000_0000_0000_0000;
array[35424] <= 16'b0000_0000_0000_0000;
array[35425] <= 16'b0000_0000_0000_0000;
array[35426] <= 16'b0000_0000_0000_0000;
array[35427] <= 16'b0000_0000_0000_0000;
array[35428] <= 16'b0000_0000_0000_0000;
array[35429] <= 16'b0000_0000_0000_0000;
array[35430] <= 16'b0000_0000_0000_0000;
array[35431] <= 16'b0000_0000_0000_0000;
array[35432] <= 16'b0000_0000_0000_0000;
array[35433] <= 16'b0000_0000_0000_0000;
array[35434] <= 16'b0000_0000_0000_0000;
array[35435] <= 16'b0000_0000_0000_0000;
array[35436] <= 16'b0000_0000_0000_0000;
array[35437] <= 16'b0000_0000_0000_0000;
array[35438] <= 16'b0000_0000_0000_0000;
array[35439] <= 16'b0000_0000_0000_0000;
array[35440] <= 16'b0000_0000_0000_0000;
array[35441] <= 16'b0000_0000_0000_0000;
array[35442] <= 16'b0000_0000_0000_0000;
array[35443] <= 16'b0000_0000_0000_0000;
array[35444] <= 16'b0000_0000_0000_0000;
array[35445] <= 16'b0000_0000_0000_0000;
array[35446] <= 16'b0000_0000_0000_0000;
array[35447] <= 16'b0000_0000_0000_0000;
array[35448] <= 16'b0000_0000_0000_0000;
array[35449] <= 16'b0000_0000_0000_0000;
array[35450] <= 16'b0000_0000_0000_0000;
array[35451] <= 16'b0000_0000_0000_0000;
array[35452] <= 16'b0000_0000_0000_0000;
array[35453] <= 16'b0000_0000_0000_0000;
array[35454] <= 16'b0000_0000_0000_0000;
array[35455] <= 16'b0000_0000_0000_0000;
array[35456] <= 16'b0000_0000_0000_0000;
array[35457] <= 16'b0000_0000_0000_0000;
array[35458] <= 16'b0000_0000_0000_0000;
array[35459] <= 16'b0000_0000_0000_0000;
array[35460] <= 16'b0000_0000_0000_0000;
array[35461] <= 16'b0000_0000_0000_0000;
array[35462] <= 16'b0000_0000_0000_0000;
array[35463] <= 16'b0000_0000_0000_0000;
array[35464] <= 16'b0000_0000_0000_0000;
array[35465] <= 16'b0000_0000_0000_0000;
array[35466] <= 16'b0000_0000_0000_0000;
array[35467] <= 16'b0000_0000_0000_0000;
array[35468] <= 16'b0000_0000_0000_0000;
array[35469] <= 16'b0000_0000_0000_0000;
array[35470] <= 16'b0000_0000_0000_0000;
array[35471] <= 16'b0000_0000_0000_0000;
array[35472] <= 16'b0000_0000_0000_0000;
array[35473] <= 16'b0000_0000_0000_0000;
array[35474] <= 16'b0000_0000_0000_0000;
array[35475] <= 16'b0000_0000_0000_0000;
array[35476] <= 16'b0000_0000_0000_0000;
array[35477] <= 16'b0000_0000_0000_0000;
array[35478] <= 16'b0000_0000_0000_0000;
array[35479] <= 16'b0000_0000_0000_0000;
array[35480] <= 16'b0000_0000_0000_0000;
array[35481] <= 16'b0000_0000_0000_0000;
array[35482] <= 16'b0000_0000_0000_0000;
array[35483] <= 16'b0000_0000_0000_0000;
array[35484] <= 16'b0000_0000_0000_0000;
array[35485] <= 16'b0000_0000_0000_0000;
array[35486] <= 16'b0000_0000_0000_0000;
array[35487] <= 16'b0000_0000_0000_0000;
array[35488] <= 16'b0000_0000_0000_0000;
array[35489] <= 16'b0000_0000_0000_0000;
array[35490] <= 16'b0000_0000_0000_0000;
array[35491] <= 16'b0000_0000_0000_0000;
array[35492] <= 16'b0000_0000_0000_0000;
array[35493] <= 16'b0000_0000_0000_0000;
array[35494] <= 16'b0000_0000_0000_0000;
array[35495] <= 16'b0000_0000_0000_0000;
array[35496] <= 16'b0000_0000_0000_0000;
array[35497] <= 16'b0000_0000_0000_0000;
array[35498] <= 16'b0000_0000_0000_0000;
array[35499] <= 16'b0000_0000_0000_0000;
array[35500] <= 16'b0000_0000_0000_0000;
array[35501] <= 16'b0000_0000_0000_0000;
array[35502] <= 16'b0000_0000_0000_0000;
array[35503] <= 16'b0000_0000_0000_0000;
array[35504] <= 16'b0000_0000_0000_0000;
array[35505] <= 16'b0000_0000_0000_0000;
array[35506] <= 16'b0000_0000_0000_0000;
array[35507] <= 16'b0000_0000_0000_0000;
array[35508] <= 16'b0000_0000_0000_0000;
array[35509] <= 16'b0000_0000_0000_0000;
array[35510] <= 16'b0000_0000_0000_0000;
array[35511] <= 16'b0000_0000_0000_0000;
array[35512] <= 16'b0000_0000_0000_0000;
array[35513] <= 16'b0000_0000_0000_0000;
array[35514] <= 16'b0000_0000_0000_0000;
array[35515] <= 16'b0000_0000_0000_0000;
array[35516] <= 16'b0000_0000_0000_0000;
array[35517] <= 16'b0000_0000_0000_0000;
array[35518] <= 16'b0000_0000_0000_0000;
array[35519] <= 16'b0000_0000_0000_0000;
array[35520] <= 16'b0000_0000_0000_0000;
array[35521] <= 16'b0000_0000_0000_0000;
array[35522] <= 16'b0000_0000_0000_0000;
array[35523] <= 16'b0000_0000_0000_0000;
array[35524] <= 16'b0000_0000_0000_0000;
array[35525] <= 16'b0000_0000_0000_0000;
array[35526] <= 16'b0000_0000_0000_0000;
array[35527] <= 16'b0000_0000_0000_0000;
array[35528] <= 16'b0000_0000_0000_0000;
array[35529] <= 16'b0000_0000_0000_0000;
array[35530] <= 16'b0000_0000_0000_0000;
array[35531] <= 16'b0000_0000_0000_0000;
array[35532] <= 16'b0000_0000_0000_0000;
array[35533] <= 16'b0000_0000_0000_0000;
array[35534] <= 16'b0000_0000_0000_0000;
array[35535] <= 16'b0000_0000_0000_0000;
array[35536] <= 16'b0000_0000_0000_0000;
array[35537] <= 16'b0000_0000_0000_0000;
array[35538] <= 16'b0000_0000_0000_0000;
array[35539] <= 16'b0000_0000_0000_0000;
array[35540] <= 16'b0000_0000_0000_0000;
array[35541] <= 16'b0000_0000_0000_0000;
array[35542] <= 16'b0000_0000_0000_0000;
array[35543] <= 16'b0000_0000_0000_0000;
array[35544] <= 16'b0000_0000_0000_0000;
array[35545] <= 16'b0000_0000_0000_0000;
array[35546] <= 16'b0000_0000_0000_0000;
array[35547] <= 16'b0000_0000_0000_0000;
array[35548] <= 16'b0000_0000_0000_0000;
array[35549] <= 16'b0000_0000_0000_0000;
array[35550] <= 16'b0000_0000_0000_0000;
array[35551] <= 16'b0000_0000_0000_0000;
array[35552] <= 16'b0000_0000_0000_0000;
array[35553] <= 16'b0000_0000_0000_0000;
array[35554] <= 16'b0000_0000_0000_0000;
array[35555] <= 16'b0000_0000_0000_0000;
array[35556] <= 16'b0000_0000_0000_0000;
array[35557] <= 16'b0000_0000_0000_0000;
array[35558] <= 16'b0000_0000_0000_0000;
array[35559] <= 16'b0000_0000_0000_0000;
array[35560] <= 16'b0000_0000_0000_0000;
array[35561] <= 16'b0000_0000_0000_0000;
array[35562] <= 16'b0000_0000_0000_0000;
array[35563] <= 16'b0000_0000_0000_0000;
array[35564] <= 16'b0000_0000_0000_0000;
array[35565] <= 16'b0000_0000_0000_0000;
array[35566] <= 16'b0000_0000_0000_0000;
array[35567] <= 16'b0000_0000_0000_0000;
array[35568] <= 16'b0000_0000_0000_0000;
array[35569] <= 16'b0000_0000_0000_0000;
array[35570] <= 16'b0000_0000_0000_0000;
array[35571] <= 16'b0000_0000_0000_0000;
array[35572] <= 16'b0000_0000_0000_0000;
array[35573] <= 16'b0000_0000_0000_0000;
array[35574] <= 16'b0000_0000_0000_0000;
array[35575] <= 16'b0000_0000_0000_0000;
array[35576] <= 16'b0000_0000_0000_0000;
array[35577] <= 16'b0000_0000_0000_0000;
array[35578] <= 16'b0000_0000_0000_0000;
array[35579] <= 16'b0000_0000_0000_0000;
array[35580] <= 16'b0000_0000_0000_0000;
array[35581] <= 16'b0000_0000_0000_0000;
array[35582] <= 16'b0000_0000_0000_0000;
array[35583] <= 16'b0000_0000_0000_0000;
array[35584] <= 16'b0000_0000_0000_0000;
array[35585] <= 16'b0000_0000_0000_0000;
array[35586] <= 16'b0000_0000_0000_0000;
array[35587] <= 16'b0000_0000_0000_0000;
array[35588] <= 16'b0000_0000_0000_0000;
array[35589] <= 16'b0000_0000_0000_0000;
array[35590] <= 16'b0000_0000_0000_0000;
array[35591] <= 16'b0000_0000_0000_0000;
array[35592] <= 16'b0000_0000_0000_0000;
array[35593] <= 16'b0000_0000_0000_0000;
array[35594] <= 16'b0000_0000_0000_0000;
array[35595] <= 16'b0000_0000_0000_0000;
array[35596] <= 16'b0000_0000_0000_0000;
array[35597] <= 16'b0000_0000_0000_0000;
array[35598] <= 16'b0000_0000_0000_0000;
array[35599] <= 16'b0000_0000_0000_0000;
array[35600] <= 16'b0000_0000_0000_0000;
array[35601] <= 16'b0000_0000_0000_0000;
array[35602] <= 16'b0000_0000_0000_0000;
array[35603] <= 16'b0000_0000_0000_0000;
array[35604] <= 16'b0000_0000_0000_0000;
array[35605] <= 16'b0000_0000_0000_0000;
array[35606] <= 16'b0000_0000_0000_0000;
array[35607] <= 16'b0000_0000_0000_0000;
array[35608] <= 16'b0000_0000_0000_0000;
array[35609] <= 16'b0000_0000_0000_0000;
array[35610] <= 16'b0000_0000_0000_0000;
array[35611] <= 16'b0000_0000_0000_0000;
array[35612] <= 16'b0000_0000_0000_0000;
array[35613] <= 16'b0000_0000_0000_0000;
array[35614] <= 16'b0000_0000_0000_0000;
array[35615] <= 16'b0000_0000_0000_0000;
array[35616] <= 16'b0000_0000_0000_0000;
array[35617] <= 16'b0000_0000_0000_0000;
array[35618] <= 16'b0000_0000_0000_0000;
array[35619] <= 16'b0000_0000_0000_0000;
array[35620] <= 16'b0000_0000_0000_0000;
array[35621] <= 16'b0000_0000_0000_0000;
array[35622] <= 16'b0000_0000_0000_0000;
array[35623] <= 16'b0000_0000_0000_0000;
array[35624] <= 16'b0000_0000_0000_0000;
array[35625] <= 16'b0000_0000_0000_0000;
array[35626] <= 16'b0000_0000_0000_0000;
array[35627] <= 16'b0000_0000_0000_0000;
array[35628] <= 16'b0000_0000_0000_0000;
array[35629] <= 16'b0000_0000_0000_0000;
array[35630] <= 16'b0000_0000_0000_0000;
array[35631] <= 16'b0000_0000_0000_0000;
array[35632] <= 16'b0000_0000_0000_0000;
array[35633] <= 16'b0000_0000_0000_0000;
array[35634] <= 16'b0000_0000_0000_0000;
array[35635] <= 16'b0000_0000_0000_0000;
array[35636] <= 16'b0000_0000_0000_0000;
array[35637] <= 16'b0000_0000_0000_0000;
array[35638] <= 16'b0000_0000_0000_0000;
array[35639] <= 16'b0000_0000_0000_0000;
array[35640] <= 16'b0000_0000_0000_0000;
array[35641] <= 16'b0000_0000_0000_0000;
array[35642] <= 16'b0000_0000_0000_0000;
array[35643] <= 16'b0000_0000_0000_0000;
array[35644] <= 16'b0000_0000_0000_0000;
array[35645] <= 16'b0000_0000_0000_0000;
array[35646] <= 16'b0000_0000_0000_0000;
array[35647] <= 16'b0000_0000_0000_0000;
array[35648] <= 16'b0000_0000_0000_0000;
array[35649] <= 16'b0000_0000_0000_0000;
array[35650] <= 16'b0000_0000_0000_0000;
array[35651] <= 16'b0000_0000_0000_0000;
array[35652] <= 16'b0000_0000_0000_0000;
array[35653] <= 16'b0000_0000_0000_0000;
array[35654] <= 16'b0000_0000_0000_0000;
array[35655] <= 16'b0000_0000_0000_0000;
array[35656] <= 16'b0000_0000_0000_0000;
array[35657] <= 16'b0000_0000_0000_0000;
array[35658] <= 16'b0000_0000_0000_0000;
array[35659] <= 16'b0000_0000_0000_0000;
array[35660] <= 16'b0000_0000_0000_0000;
array[35661] <= 16'b0000_0000_0000_0000;
array[35662] <= 16'b0000_0000_0000_0000;
array[35663] <= 16'b0000_0000_0000_0000;
array[35664] <= 16'b0000_0000_0000_0000;
array[35665] <= 16'b0000_0000_0000_0000;
array[35666] <= 16'b0000_0000_0000_0000;
array[35667] <= 16'b0000_0000_0000_0000;
array[35668] <= 16'b0000_0000_0000_0000;
array[35669] <= 16'b0000_0000_0000_0000;
array[35670] <= 16'b0000_0000_0000_0000;
array[35671] <= 16'b0000_0000_0000_0000;
array[35672] <= 16'b0000_0000_0000_0000;
array[35673] <= 16'b0000_0000_0000_0000;
array[35674] <= 16'b0000_0000_0000_0000;
array[35675] <= 16'b0000_0000_0000_0000;
array[35676] <= 16'b0000_0000_0000_0000;
array[35677] <= 16'b0000_0000_0000_0000;
array[35678] <= 16'b0000_0000_0000_0000;
array[35679] <= 16'b0000_0000_0000_0000;
array[35680] <= 16'b0000_0000_0000_0000;
array[35681] <= 16'b0000_0000_0000_0000;
array[35682] <= 16'b0000_0000_0000_0000;
array[35683] <= 16'b0000_0000_0000_0000;
array[35684] <= 16'b0000_0000_0000_0000;
array[35685] <= 16'b0000_0000_0000_0000;
array[35686] <= 16'b0000_0000_0000_0000;
array[35687] <= 16'b0000_0000_0000_0000;
array[35688] <= 16'b0000_0000_0000_0000;
array[35689] <= 16'b0000_0000_0000_0000;
array[35690] <= 16'b0000_0000_0000_0000;
array[35691] <= 16'b0000_0000_0000_0000;
array[35692] <= 16'b0000_0000_0000_0000;
array[35693] <= 16'b0000_0000_0000_0000;
array[35694] <= 16'b0000_0000_0000_0000;
array[35695] <= 16'b0000_0000_0000_0000;
array[35696] <= 16'b0000_0000_0000_0000;
array[35697] <= 16'b0000_0000_0000_0000;
array[35698] <= 16'b0000_0000_0000_0000;
array[35699] <= 16'b0000_0000_0000_0000;
array[35700] <= 16'b0000_0000_0000_0000;
array[35701] <= 16'b0000_0000_0000_0000;
array[35702] <= 16'b0000_0000_0000_0000;
array[35703] <= 16'b0000_0000_0000_0000;
array[35704] <= 16'b0000_0000_0000_0000;
array[35705] <= 16'b0000_0000_0000_0000;
array[35706] <= 16'b0000_0000_0000_0000;
array[35707] <= 16'b0000_0000_0000_0000;
array[35708] <= 16'b0000_0000_0000_0000;
array[35709] <= 16'b0000_0000_0000_0000;
array[35710] <= 16'b0000_0000_0000_0000;
array[35711] <= 16'b0000_0000_0000_0000;
array[35712] <= 16'b0000_0000_0000_0000;
array[35713] <= 16'b0000_0000_0000_0000;
array[35714] <= 16'b0000_0000_0000_0000;
array[35715] <= 16'b0000_0000_0000_0000;
array[35716] <= 16'b0000_0000_0000_0000;
array[35717] <= 16'b0000_0000_0000_0000;
array[35718] <= 16'b0000_0000_0000_0000;
array[35719] <= 16'b0000_0000_0000_0000;
array[35720] <= 16'b0000_0000_0000_0000;
array[35721] <= 16'b0000_0000_0000_0000;
array[35722] <= 16'b0000_0000_0000_0000;
array[35723] <= 16'b0000_0000_0000_0000;
array[35724] <= 16'b0000_0000_0000_0000;
array[35725] <= 16'b0000_0000_0000_0000;
array[35726] <= 16'b0000_0000_0000_0000;
array[35727] <= 16'b0000_0000_0000_0000;
array[35728] <= 16'b0000_0000_0000_0000;
array[35729] <= 16'b0000_0000_0000_0000;
array[35730] <= 16'b0000_0000_0000_0000;
array[35731] <= 16'b0000_0000_0000_0000;
array[35732] <= 16'b0000_0000_0000_0000;
array[35733] <= 16'b0000_0000_0000_0000;
array[35734] <= 16'b0000_0000_0000_0000;
array[35735] <= 16'b0000_0000_0000_0000;
array[35736] <= 16'b0000_0000_0000_0000;
array[35737] <= 16'b0000_0000_0000_0000;
array[35738] <= 16'b0000_0000_0000_0000;
array[35739] <= 16'b0000_0000_0000_0000;
array[35740] <= 16'b0000_0000_0000_0000;
array[35741] <= 16'b0000_0000_0000_0000;
array[35742] <= 16'b0000_0000_0000_0000;
array[35743] <= 16'b0000_0000_0000_0000;
array[35744] <= 16'b0000_0000_0000_0000;
array[35745] <= 16'b0000_0000_0000_0000;
array[35746] <= 16'b0000_0000_0000_0000;
array[35747] <= 16'b0000_0000_0000_0000;
array[35748] <= 16'b0000_0000_0000_0000;
array[35749] <= 16'b0000_0000_0000_0000;
array[35750] <= 16'b0000_0000_0000_0000;
array[35751] <= 16'b0000_0000_0000_0000;
array[35752] <= 16'b0000_0000_0000_0000;
array[35753] <= 16'b0000_0000_0000_0000;
array[35754] <= 16'b0000_0000_0000_0000;
array[35755] <= 16'b0000_0000_0000_0000;
array[35756] <= 16'b0000_0000_0000_0000;
array[35757] <= 16'b0000_0000_0000_0000;
array[35758] <= 16'b0000_0000_0000_0000;
array[35759] <= 16'b0000_0000_0000_0000;
array[35760] <= 16'b0000_0000_0000_0000;
array[35761] <= 16'b0000_0000_0000_0000;
array[35762] <= 16'b0000_0000_0000_0000;
array[35763] <= 16'b0000_0000_0000_0000;
array[35764] <= 16'b0000_0000_0000_0000;
array[35765] <= 16'b0000_0000_0000_0000;
array[35766] <= 16'b0000_0000_0000_0000;
array[35767] <= 16'b0000_0000_0000_0000;
array[35768] <= 16'b0000_0000_0000_0000;
array[35769] <= 16'b0000_0000_0000_0000;
array[35770] <= 16'b0000_0000_0000_0000;
array[35771] <= 16'b0000_0000_0000_0000;
array[35772] <= 16'b0000_0000_0000_0000;
array[35773] <= 16'b0000_0000_0000_0000;
array[35774] <= 16'b0000_0000_0000_0000;
array[35775] <= 16'b0000_0000_0000_0000;
array[35776] <= 16'b0000_0000_0000_0000;
array[35777] <= 16'b0000_0000_0000_0000;
array[35778] <= 16'b0000_0000_0000_0000;
array[35779] <= 16'b0000_0000_0000_0000;
array[35780] <= 16'b0000_0000_0000_0000;
array[35781] <= 16'b0000_0000_0000_0000;
array[35782] <= 16'b0000_0000_0000_0000;
array[35783] <= 16'b0000_0000_0000_0000;
array[35784] <= 16'b0000_0000_0000_0000;
array[35785] <= 16'b0000_0000_0000_0000;
array[35786] <= 16'b0000_0000_0000_0000;
array[35787] <= 16'b0000_0000_0000_0000;
array[35788] <= 16'b0000_0000_0000_0000;
array[35789] <= 16'b0000_0000_0000_0000;
array[35790] <= 16'b0000_0000_0000_0000;
array[35791] <= 16'b0000_0000_0000_0000;
array[35792] <= 16'b0000_0000_0000_0000;
array[35793] <= 16'b0000_0000_0000_0000;
array[35794] <= 16'b0000_0000_0000_0000;
array[35795] <= 16'b0000_0000_0000_0000;
array[35796] <= 16'b0000_0000_0000_0000;
array[35797] <= 16'b0000_0000_0000_0000;
array[35798] <= 16'b0000_0000_0000_0000;
array[35799] <= 16'b0000_0000_0000_0000;
array[35800] <= 16'b0000_0000_0000_0000;
array[35801] <= 16'b0000_0000_0000_0000;
array[35802] <= 16'b0000_0000_0000_0000;
array[35803] <= 16'b0000_0000_0000_0000;
array[35804] <= 16'b0000_0000_0000_0000;
array[35805] <= 16'b0000_0000_0000_0000;
array[35806] <= 16'b0000_0000_0000_0000;
array[35807] <= 16'b0000_0000_0000_0000;
array[35808] <= 16'b0000_0000_0000_0000;
array[35809] <= 16'b0000_0000_0000_0000;
array[35810] <= 16'b0000_0000_0000_0000;
array[35811] <= 16'b0000_0000_0000_0000;
array[35812] <= 16'b0000_0000_0000_0000;
array[35813] <= 16'b0000_0000_0000_0000;
array[35814] <= 16'b0000_0000_0000_0000;
array[35815] <= 16'b0000_0000_0000_0000;
array[35816] <= 16'b0000_0000_0000_0000;
array[35817] <= 16'b0000_0000_0000_0000;
array[35818] <= 16'b0000_0000_0000_0000;
array[35819] <= 16'b0000_0000_0000_0000;
array[35820] <= 16'b0000_0000_0000_0000;
array[35821] <= 16'b0000_0000_0000_0000;
array[35822] <= 16'b0000_0000_0000_0000;
array[35823] <= 16'b0000_0000_0000_0000;
array[35824] <= 16'b0000_0000_0000_0000;
array[35825] <= 16'b0000_0000_0000_0000;
array[35826] <= 16'b0000_0000_0000_0000;
array[35827] <= 16'b0000_0000_0000_0000;
array[35828] <= 16'b0000_0000_0000_0000;
array[35829] <= 16'b0000_0000_0000_0000;
array[35830] <= 16'b0000_0000_0000_0000;
array[35831] <= 16'b0000_0000_0000_0000;
array[35832] <= 16'b0000_0000_0000_0000;
array[35833] <= 16'b0000_0000_0000_0000;
array[35834] <= 16'b0000_0000_0000_0000;
array[35835] <= 16'b0000_0000_0000_0000;
array[35836] <= 16'b0000_0000_0000_0000;
array[35837] <= 16'b0000_0000_0000_0000;
array[35838] <= 16'b0000_0000_0000_0000;
array[35839] <= 16'b0000_0000_0000_0000;
array[35840] <= 16'b0000_0000_0000_0000;
array[35841] <= 16'b0000_0000_0000_0000;
array[35842] <= 16'b0000_0000_0000_0000;
array[35843] <= 16'b0000_0000_0000_0000;
array[35844] <= 16'b0000_0000_0000_0000;
array[35845] <= 16'b0000_0000_0000_0000;
array[35846] <= 16'b0000_0000_0000_0000;
array[35847] <= 16'b0000_0000_0000_0000;
array[35848] <= 16'b0000_0000_0000_0000;
array[35849] <= 16'b0000_0000_0000_0000;
array[35850] <= 16'b0000_0000_0000_0000;
array[35851] <= 16'b0000_0000_0000_0000;
array[35852] <= 16'b0000_0000_0000_0000;
array[35853] <= 16'b0000_0000_0000_0000;
array[35854] <= 16'b0000_0000_0000_0000;
array[35855] <= 16'b0000_0000_0000_0000;
array[35856] <= 16'b0000_0000_0000_0000;
array[35857] <= 16'b0000_0000_0000_0000;
array[35858] <= 16'b0000_0000_0000_0000;
array[35859] <= 16'b0000_0000_0000_0000;
array[35860] <= 16'b0000_0000_0000_0000;
array[35861] <= 16'b0000_0000_0000_0000;
array[35862] <= 16'b0000_0000_0000_0000;
array[35863] <= 16'b0000_0000_0000_0000;
array[35864] <= 16'b0000_0000_0000_0000;
array[35865] <= 16'b0000_0000_0000_0000;
array[35866] <= 16'b0000_0000_0000_0000;
array[35867] <= 16'b0000_0000_0000_0000;
array[35868] <= 16'b0000_0000_0000_0000;
array[35869] <= 16'b0000_0000_0000_0000;
array[35870] <= 16'b0000_0000_0000_0000;
array[35871] <= 16'b0000_0000_0000_0000;
array[35872] <= 16'b0000_0000_0000_0000;
array[35873] <= 16'b0000_0000_0000_0000;
array[35874] <= 16'b0000_0000_0000_0000;
array[35875] <= 16'b0000_0000_0000_0000;
array[35876] <= 16'b0000_0000_0000_0000;
array[35877] <= 16'b0000_0000_0000_0000;
array[35878] <= 16'b0000_0000_0000_0000;
array[35879] <= 16'b0000_0000_0000_0000;
array[35880] <= 16'b0000_0000_0000_0000;
array[35881] <= 16'b0000_0000_0000_0000;
array[35882] <= 16'b0000_0000_0000_0000;
array[35883] <= 16'b0000_0000_0000_0000;
array[35884] <= 16'b0000_0000_0000_0000;
array[35885] <= 16'b0000_0000_0000_0000;
array[35886] <= 16'b0000_0000_0000_0000;
array[35887] <= 16'b0000_0000_0000_0000;
array[35888] <= 16'b0000_0000_0000_0000;
array[35889] <= 16'b0000_0000_0000_0000;
array[35890] <= 16'b0000_0000_0000_0000;
array[35891] <= 16'b0000_0000_0000_0000;
array[35892] <= 16'b0000_0000_0000_0000;
array[35893] <= 16'b0000_0000_0000_0000;
array[35894] <= 16'b0000_0000_0000_0000;
array[35895] <= 16'b0000_0000_0000_0000;
array[35896] <= 16'b0000_0000_0000_0000;
array[35897] <= 16'b0000_0000_0000_0000;
array[35898] <= 16'b0000_0000_0000_0000;
array[35899] <= 16'b0000_0000_0000_0000;
array[35900] <= 16'b0000_0000_0000_0000;
array[35901] <= 16'b0000_0000_0000_0000;
array[35902] <= 16'b0000_0000_0000_0000;
array[35903] <= 16'b0000_0000_0000_0000;
array[35904] <= 16'b0000_0000_0000_0000;
array[35905] <= 16'b0000_0000_0000_0000;
array[35906] <= 16'b0000_0000_0000_0000;
array[35907] <= 16'b0000_0000_0000_0000;
array[35908] <= 16'b0000_0000_0000_0000;
array[35909] <= 16'b0000_0000_0000_0000;
array[35910] <= 16'b0000_0000_0000_0000;
array[35911] <= 16'b0000_0000_0000_0000;
array[35912] <= 16'b0000_0000_0000_0000;
array[35913] <= 16'b0000_0000_0000_0000;
array[35914] <= 16'b0000_0000_0000_0000;
array[35915] <= 16'b0000_0000_0000_0000;
array[35916] <= 16'b0000_0000_0000_0000;
array[35917] <= 16'b0000_0000_0000_0000;
array[35918] <= 16'b0000_0000_0000_0000;
array[35919] <= 16'b0000_0000_0000_0000;
array[35920] <= 16'b0000_0000_0000_0000;
array[35921] <= 16'b0000_0000_0000_0000;
array[35922] <= 16'b0000_0000_0000_0000;
array[35923] <= 16'b0000_0000_0000_0000;
array[35924] <= 16'b0000_0000_0000_0000;
array[35925] <= 16'b0000_0000_0000_0000;
array[35926] <= 16'b0000_0000_0000_0000;
array[35927] <= 16'b0000_0000_0000_0000;
array[35928] <= 16'b0000_0000_0000_0000;
array[35929] <= 16'b0000_0000_0000_0000;
array[35930] <= 16'b0000_0000_0000_0000;
array[35931] <= 16'b0000_0000_0000_0000;
array[35932] <= 16'b0000_0000_0000_0000;
array[35933] <= 16'b0000_0000_0000_0000;
array[35934] <= 16'b0000_0000_0000_0000;
array[35935] <= 16'b0000_0000_0000_0000;
array[35936] <= 16'b0000_0000_0000_0000;
array[35937] <= 16'b0000_0000_0000_0000;
array[35938] <= 16'b0000_0000_0000_0000;
array[35939] <= 16'b0000_0000_0000_0000;
array[35940] <= 16'b0000_0000_0000_0000;
array[35941] <= 16'b0000_0000_0000_0000;
array[35942] <= 16'b0000_0000_0000_0000;
array[35943] <= 16'b0000_0000_0000_0000;
array[35944] <= 16'b0000_0000_0000_0000;
array[35945] <= 16'b0000_0000_0000_0000;
array[35946] <= 16'b0000_0000_0000_0000;
array[35947] <= 16'b0000_0000_0000_0000;
array[35948] <= 16'b0000_0000_0000_0000;
array[35949] <= 16'b0000_0000_0000_0000;
array[35950] <= 16'b0000_0000_0000_0000;
array[35951] <= 16'b0000_0000_0000_0000;
array[35952] <= 16'b0000_0000_0000_0000;
array[35953] <= 16'b0000_0000_0000_0000;
array[35954] <= 16'b0000_0000_0000_0000;
array[35955] <= 16'b0000_0000_0000_0000;
array[35956] <= 16'b0000_0000_0000_0000;
array[35957] <= 16'b0000_0000_0000_0000;
array[35958] <= 16'b0000_0000_0000_0000;
array[35959] <= 16'b0000_0000_0000_0000;
array[35960] <= 16'b0000_0000_0000_0000;
array[35961] <= 16'b0000_0000_0000_0000;
array[35962] <= 16'b0000_0000_0000_0000;
array[35963] <= 16'b0000_0000_0000_0000;
array[35964] <= 16'b0000_0000_0000_0000;
array[35965] <= 16'b0000_0000_0000_0000;
array[35966] <= 16'b0000_0000_0000_0000;
array[35967] <= 16'b0000_0000_0000_0000;
array[35968] <= 16'b0000_0000_0000_0000;
array[35969] <= 16'b0000_0000_0000_0000;
array[35970] <= 16'b0000_0000_0000_0000;
array[35971] <= 16'b0000_0000_0000_0000;
array[35972] <= 16'b0000_0000_0000_0000;
array[35973] <= 16'b0000_0000_0000_0000;
array[35974] <= 16'b0000_0000_0000_0000;
array[35975] <= 16'b0000_0000_0000_0000;
array[35976] <= 16'b0000_0000_0000_0000;
array[35977] <= 16'b0000_0000_0000_0000;
array[35978] <= 16'b0000_0000_0000_0000;
array[35979] <= 16'b0000_0000_0000_0000;
array[35980] <= 16'b0000_0000_0000_0000;
array[35981] <= 16'b0000_0000_0000_0000;
array[35982] <= 16'b0000_0000_0000_0000;
array[35983] <= 16'b0000_0000_0000_0000;
array[35984] <= 16'b0000_0000_0000_0000;
array[35985] <= 16'b0000_0000_0000_0000;
array[35986] <= 16'b0000_0000_0000_0000;
array[35987] <= 16'b0000_0000_0000_0000;
array[35988] <= 16'b0000_0000_0000_0000;
array[35989] <= 16'b0000_0000_0000_0000;
array[35990] <= 16'b0000_0000_0000_0000;
array[35991] <= 16'b0000_0000_0000_0000;
array[35992] <= 16'b0000_0000_0000_0000;
array[35993] <= 16'b0000_0000_0000_0000;
array[35994] <= 16'b0000_0000_0000_0000;
array[35995] <= 16'b0000_0000_0000_0000;
array[35996] <= 16'b0000_0000_0000_0000;
array[35997] <= 16'b0000_0000_0000_0000;
array[35998] <= 16'b0000_0000_0000_0000;
array[35999] <= 16'b0000_0000_0000_0000;
array[36000] <= 16'b0000_0000_0000_0000;
array[36001] <= 16'b0000_0000_0000_0000;
array[36002] <= 16'b0000_0000_0000_0000;
array[36003] <= 16'b0000_0000_0000_0000;
array[36004] <= 16'b0000_0000_0000_0000;
array[36005] <= 16'b0000_0000_0000_0000;
array[36006] <= 16'b0000_0000_0000_0000;
array[36007] <= 16'b0000_0000_0000_0000;
array[36008] <= 16'b0000_0000_0000_0000;
array[36009] <= 16'b0000_0000_0000_0000;
array[36010] <= 16'b0000_0000_0000_0000;
array[36011] <= 16'b0000_0000_0000_0000;
array[36012] <= 16'b0000_0000_0000_0000;
array[36013] <= 16'b0000_0000_0000_0000;
array[36014] <= 16'b0000_0000_0000_0000;
array[36015] <= 16'b0000_0000_0000_0000;
array[36016] <= 16'b0000_0000_0000_0000;
array[36017] <= 16'b0000_0000_0000_0000;
array[36018] <= 16'b0000_0000_0000_0000;
array[36019] <= 16'b0000_0000_0000_0000;
array[36020] <= 16'b0000_0000_0000_0000;
array[36021] <= 16'b0000_0000_0000_0000;
array[36022] <= 16'b0000_0000_0000_0000;
array[36023] <= 16'b0000_0000_0000_0000;
array[36024] <= 16'b0000_0000_0000_0000;
array[36025] <= 16'b0000_0000_0000_0000;
array[36026] <= 16'b0000_0000_0000_0000;
array[36027] <= 16'b0000_0000_0000_0000;
array[36028] <= 16'b0000_0000_0000_0000;
array[36029] <= 16'b0000_0000_0000_0000;
array[36030] <= 16'b0000_0000_0000_0000;
array[36031] <= 16'b0000_0000_0000_0000;
array[36032] <= 16'b0000_0000_0000_0000;
array[36033] <= 16'b0000_0000_0000_0000;
array[36034] <= 16'b0000_0000_0000_0000;
array[36035] <= 16'b0000_0000_0000_0000;
array[36036] <= 16'b0000_0000_0000_0000;
array[36037] <= 16'b0000_0000_0000_0000;
array[36038] <= 16'b0000_0000_0000_0000;
array[36039] <= 16'b0000_0000_0000_0000;
array[36040] <= 16'b0000_0000_0000_0000;
array[36041] <= 16'b0000_0000_0000_0000;
array[36042] <= 16'b0000_0000_0000_0000;
array[36043] <= 16'b0000_0000_0000_0000;
array[36044] <= 16'b0000_0000_0000_0000;
array[36045] <= 16'b0000_0000_0000_0000;
array[36046] <= 16'b0000_0000_0000_0000;
array[36047] <= 16'b0000_0000_0000_0000;
array[36048] <= 16'b0000_0000_0000_0000;
array[36049] <= 16'b0000_0000_0000_0000;
array[36050] <= 16'b0000_0000_0000_0000;
array[36051] <= 16'b0000_0000_0000_0000;
array[36052] <= 16'b0000_0000_0000_0000;
array[36053] <= 16'b0000_0000_0000_0000;
array[36054] <= 16'b0000_0000_0000_0000;
array[36055] <= 16'b0000_0000_0000_0000;
array[36056] <= 16'b0000_0000_0000_0000;
array[36057] <= 16'b0000_0000_0000_0000;
array[36058] <= 16'b0000_0000_0000_0000;
array[36059] <= 16'b0000_0000_0000_0000;
array[36060] <= 16'b0000_0000_0000_0000;
array[36061] <= 16'b0000_0000_0000_0000;
array[36062] <= 16'b0000_0000_0000_0000;
array[36063] <= 16'b0000_0000_0000_0000;
array[36064] <= 16'b0000_0000_0000_0000;
array[36065] <= 16'b0000_0000_0000_0000;
array[36066] <= 16'b0000_0000_0000_0000;
array[36067] <= 16'b0000_0000_0000_0000;
array[36068] <= 16'b0000_0000_0000_0000;
array[36069] <= 16'b0000_0000_0000_0000;
array[36070] <= 16'b0000_0000_0000_0000;
array[36071] <= 16'b0000_0000_0000_0000;
array[36072] <= 16'b0000_0000_0000_0000;
array[36073] <= 16'b0000_0000_0000_0000;
array[36074] <= 16'b0000_0000_0000_0000;
array[36075] <= 16'b0000_0000_0000_0000;
array[36076] <= 16'b0000_0000_0000_0000;
array[36077] <= 16'b0000_0000_0000_0000;
array[36078] <= 16'b0000_0000_0000_0000;
array[36079] <= 16'b0000_0000_0000_0000;
array[36080] <= 16'b0000_0000_0000_0000;
array[36081] <= 16'b0000_0000_0000_0000;
array[36082] <= 16'b0000_0000_0000_0000;
array[36083] <= 16'b0000_0000_0000_0000;
array[36084] <= 16'b0000_0000_0000_0000;
array[36085] <= 16'b0000_0000_0000_0000;
array[36086] <= 16'b0000_0000_0000_0000;
array[36087] <= 16'b0000_0000_0000_0000;
array[36088] <= 16'b0000_0000_0000_0000;
array[36089] <= 16'b0000_0000_0000_0000;
array[36090] <= 16'b0000_0000_0000_0000;
array[36091] <= 16'b0000_0000_0000_0000;
array[36092] <= 16'b0000_0000_0000_0000;
array[36093] <= 16'b0000_0000_0000_0000;
array[36094] <= 16'b0000_0000_0000_0000;
array[36095] <= 16'b0000_0000_0000_0000;
array[36096] <= 16'b0000_0000_0000_0000;
array[36097] <= 16'b0000_0000_0000_0000;
array[36098] <= 16'b0000_0000_0000_0000;
array[36099] <= 16'b0000_0000_0000_0000;
array[36100] <= 16'b0000_0000_0000_0000;
array[36101] <= 16'b0000_0000_0000_0000;
array[36102] <= 16'b0000_0000_0000_0000;
array[36103] <= 16'b0000_0000_0000_0000;
array[36104] <= 16'b0000_0000_0000_0000;
array[36105] <= 16'b0000_0000_0000_0000;
array[36106] <= 16'b0000_0000_0000_0000;
array[36107] <= 16'b0000_0000_0000_0000;
array[36108] <= 16'b0000_0000_0000_0000;
array[36109] <= 16'b0000_0000_0000_0000;
array[36110] <= 16'b0000_0000_0000_0000;
array[36111] <= 16'b0000_0000_0000_0000;
array[36112] <= 16'b0000_0000_0000_0000;
array[36113] <= 16'b0000_0000_0000_0000;
array[36114] <= 16'b0000_0000_0000_0000;
array[36115] <= 16'b0000_0000_0000_0000;
array[36116] <= 16'b0000_0000_0000_0000;
array[36117] <= 16'b0000_0000_0000_0000;
array[36118] <= 16'b0000_0000_0000_0000;
array[36119] <= 16'b0000_0000_0000_0000;
array[36120] <= 16'b0000_0000_0000_0000;
array[36121] <= 16'b0000_0000_0000_0000;
array[36122] <= 16'b0000_0000_0000_0000;
array[36123] <= 16'b0000_0000_0000_0000;
array[36124] <= 16'b0000_0000_0000_0000;
array[36125] <= 16'b0000_0000_0000_0000;
array[36126] <= 16'b0000_0000_0000_0000;
array[36127] <= 16'b0000_0000_0000_0000;
array[36128] <= 16'b0000_0000_0000_0000;
array[36129] <= 16'b0000_0000_0000_0000;
array[36130] <= 16'b0000_0000_0000_0000;
array[36131] <= 16'b0000_0000_0000_0000;
array[36132] <= 16'b0000_0000_0000_0000;
array[36133] <= 16'b0000_0000_0000_0000;
array[36134] <= 16'b0000_0000_0000_0000;
array[36135] <= 16'b0000_0000_0000_0000;
array[36136] <= 16'b0000_0000_0000_0000;
array[36137] <= 16'b0000_0000_0000_0000;
array[36138] <= 16'b0000_0000_0000_0000;
array[36139] <= 16'b0000_0000_0000_0000;
array[36140] <= 16'b0000_0000_0000_0000;
array[36141] <= 16'b0000_0000_0000_0000;
array[36142] <= 16'b0000_0000_0000_0000;
array[36143] <= 16'b0000_0000_0000_0000;
array[36144] <= 16'b0000_0000_0000_0000;
array[36145] <= 16'b0000_0000_0000_0000;
array[36146] <= 16'b0000_0000_0000_0000;
array[36147] <= 16'b0000_0000_0000_0000;
array[36148] <= 16'b0000_0000_0000_0000;
array[36149] <= 16'b0000_0000_0000_0000;
array[36150] <= 16'b0000_0000_0000_0000;
array[36151] <= 16'b0000_0000_0000_0000;
array[36152] <= 16'b0000_0000_0000_0000;
array[36153] <= 16'b0000_0000_0000_0000;
array[36154] <= 16'b0000_0000_0000_0000;
array[36155] <= 16'b0000_0000_0000_0000;
array[36156] <= 16'b0000_0000_0000_0000;
array[36157] <= 16'b0000_0000_0000_0000;
array[36158] <= 16'b0000_0000_0000_0000;
array[36159] <= 16'b0000_0000_0000_0000;
array[36160] <= 16'b0000_0000_0000_0000;
array[36161] <= 16'b0000_0000_0000_0000;
array[36162] <= 16'b0000_0000_0000_0000;
array[36163] <= 16'b0000_0000_0000_0000;
array[36164] <= 16'b0000_0000_0000_0000;
array[36165] <= 16'b0000_0000_0000_0000;
array[36166] <= 16'b0000_0000_0000_0000;
array[36167] <= 16'b0000_0000_0000_0000;
array[36168] <= 16'b0000_0000_0000_0000;
array[36169] <= 16'b0000_0000_0000_0000;
array[36170] <= 16'b0000_0000_0000_0000;
array[36171] <= 16'b0000_0000_0000_0000;
array[36172] <= 16'b0000_0000_0000_0000;
array[36173] <= 16'b0000_0000_0000_0000;
array[36174] <= 16'b0000_0000_0000_0000;
array[36175] <= 16'b0000_0000_0000_0000;
array[36176] <= 16'b0000_0000_0000_0000;
array[36177] <= 16'b0000_0000_0000_0000;
array[36178] <= 16'b0000_0000_0000_0000;
array[36179] <= 16'b0000_0000_0000_0000;
array[36180] <= 16'b0000_0000_0000_0000;
array[36181] <= 16'b0000_0000_0000_0000;
array[36182] <= 16'b0000_0000_0000_0000;
array[36183] <= 16'b0000_0000_0000_0000;
array[36184] <= 16'b0000_0000_0000_0000;
array[36185] <= 16'b0000_0000_0000_0000;
array[36186] <= 16'b0000_0000_0000_0000;
array[36187] <= 16'b0000_0000_0000_0000;
array[36188] <= 16'b0000_0000_0000_0000;
array[36189] <= 16'b0000_0000_0000_0000;
array[36190] <= 16'b0000_0000_0000_0000;
array[36191] <= 16'b0000_0000_0000_0000;
array[36192] <= 16'b0000_0000_0000_0000;
array[36193] <= 16'b0000_0000_0000_0000;
array[36194] <= 16'b0000_0000_0000_0000;
array[36195] <= 16'b0000_0000_0000_0000;
array[36196] <= 16'b0000_0000_0000_0000;
array[36197] <= 16'b0000_0000_0000_0000;
array[36198] <= 16'b0000_0000_0000_0000;
array[36199] <= 16'b0000_0000_0000_0000;
array[36200] <= 16'b0000_0000_0000_0000;
array[36201] <= 16'b0000_0000_0000_0000;
array[36202] <= 16'b0000_0000_0000_0000;
array[36203] <= 16'b0000_0000_0000_0000;
array[36204] <= 16'b0000_0000_0000_0000;
array[36205] <= 16'b0000_0000_0000_0000;
array[36206] <= 16'b0000_0000_0000_0000;
array[36207] <= 16'b0000_0000_0000_0000;
array[36208] <= 16'b0000_0000_0000_0000;
array[36209] <= 16'b0000_0000_0000_0000;
array[36210] <= 16'b0000_0000_0000_0000;
array[36211] <= 16'b0000_0000_0000_0000;
array[36212] <= 16'b0000_0000_0000_0000;
array[36213] <= 16'b0000_0000_0000_0000;
array[36214] <= 16'b0000_0000_0000_0000;
array[36215] <= 16'b0000_0000_0000_0000;
array[36216] <= 16'b0000_0000_0000_0000;
array[36217] <= 16'b0000_0000_0000_0000;
array[36218] <= 16'b0000_0000_0000_0000;
array[36219] <= 16'b0000_0000_0000_0000;
array[36220] <= 16'b0000_0000_0000_0000;
array[36221] <= 16'b0000_0000_0000_0000;
array[36222] <= 16'b0000_0000_0000_0000;
array[36223] <= 16'b0000_0000_0000_0000;
array[36224] <= 16'b0000_0000_0000_0000;
array[36225] <= 16'b0000_0000_0000_0000;
array[36226] <= 16'b0000_0000_0000_0000;
array[36227] <= 16'b0000_0000_0000_0000;
array[36228] <= 16'b0000_0000_0000_0000;
array[36229] <= 16'b0000_0000_0000_0000;
array[36230] <= 16'b0000_0000_0000_0000;
array[36231] <= 16'b0000_0000_0000_0000;
array[36232] <= 16'b0000_0000_0000_0000;
array[36233] <= 16'b0000_0000_0000_0000;
array[36234] <= 16'b0000_0000_0000_0000;
array[36235] <= 16'b0000_0000_0000_0000;
array[36236] <= 16'b0000_0000_0000_0000;
array[36237] <= 16'b0000_0000_0000_0000;
array[36238] <= 16'b0000_0000_0000_0000;
array[36239] <= 16'b0000_0000_0000_0000;
array[36240] <= 16'b0000_0000_0000_0000;
array[36241] <= 16'b0000_0000_0000_0000;
array[36242] <= 16'b0000_0000_0000_0000;
array[36243] <= 16'b0000_0000_0000_0000;
array[36244] <= 16'b0000_0000_0000_0000;
array[36245] <= 16'b0000_0000_0000_0000;
array[36246] <= 16'b0000_0000_0000_0000;
array[36247] <= 16'b0000_0000_0000_0000;
array[36248] <= 16'b0000_0000_0000_0000;
array[36249] <= 16'b0000_0000_0000_0000;
array[36250] <= 16'b0000_0000_0000_0000;
array[36251] <= 16'b0000_0000_0000_0000;
array[36252] <= 16'b0000_0000_0000_0000;
array[36253] <= 16'b0000_0000_0000_0000;
array[36254] <= 16'b0000_0000_0000_0000;
array[36255] <= 16'b0000_0000_0000_0000;
array[36256] <= 16'b0000_0000_0000_0000;
array[36257] <= 16'b0000_0000_0000_0000;
array[36258] <= 16'b0000_0000_0000_0000;
array[36259] <= 16'b0000_0000_0000_0000;
array[36260] <= 16'b0000_0000_0000_0000;
array[36261] <= 16'b0000_0000_0000_0000;
array[36262] <= 16'b0000_0000_0000_0000;
array[36263] <= 16'b0000_0000_0000_0000;
array[36264] <= 16'b0000_0000_0000_0000;
array[36265] <= 16'b0000_0000_0000_0000;
array[36266] <= 16'b0000_0000_0000_0000;
array[36267] <= 16'b0000_0000_0000_0000;
array[36268] <= 16'b0000_0000_0000_0000;
array[36269] <= 16'b0000_0000_0000_0000;
array[36270] <= 16'b0000_0000_0000_0000;
array[36271] <= 16'b0000_0000_0000_0000;
array[36272] <= 16'b0000_0000_0000_0000;
array[36273] <= 16'b0000_0000_0000_0000;
array[36274] <= 16'b0000_0000_0000_0000;
array[36275] <= 16'b0000_0000_0000_0000;
array[36276] <= 16'b0000_0000_0000_0000;
array[36277] <= 16'b0000_0000_0000_0000;
array[36278] <= 16'b0000_0000_0000_0000;
array[36279] <= 16'b0000_0000_0000_0000;
array[36280] <= 16'b0000_0000_0000_0000;
array[36281] <= 16'b0000_0000_0000_0000;
array[36282] <= 16'b0000_0000_0000_0000;
array[36283] <= 16'b0000_0000_0000_0000;
array[36284] <= 16'b0000_0000_0000_0000;
array[36285] <= 16'b0000_0000_0000_0000;
array[36286] <= 16'b0000_0000_0000_0000;
array[36287] <= 16'b0000_0000_0000_0000;
array[36288] <= 16'b0000_0000_0000_0000;
array[36289] <= 16'b0000_0000_0000_0000;
array[36290] <= 16'b0000_0000_0000_0000;
array[36291] <= 16'b0000_0000_0000_0000;
array[36292] <= 16'b0000_0000_0000_0000;
array[36293] <= 16'b0000_0000_0000_0000;
array[36294] <= 16'b0000_0000_0000_0000;
array[36295] <= 16'b0000_0000_0000_0000;
array[36296] <= 16'b0000_0000_0000_0000;
array[36297] <= 16'b0000_0000_0000_0000;
array[36298] <= 16'b0000_0000_0000_0000;
array[36299] <= 16'b0000_0000_0000_0000;
array[36300] <= 16'b0000_0000_0000_0000;
array[36301] <= 16'b0000_0000_0000_0000;
array[36302] <= 16'b0000_0000_0000_0000;
array[36303] <= 16'b0000_0000_0000_0000;
array[36304] <= 16'b0000_0000_0000_0000;
array[36305] <= 16'b0000_0000_0000_0000;
array[36306] <= 16'b0000_0000_0000_0000;
array[36307] <= 16'b0000_0000_0000_0000;
array[36308] <= 16'b0000_0000_0000_0000;
array[36309] <= 16'b0000_0000_0000_0000;
array[36310] <= 16'b0000_0000_0000_0000;
array[36311] <= 16'b0000_0000_0000_0000;
array[36312] <= 16'b0000_0000_0000_0000;
array[36313] <= 16'b0000_0000_0000_0000;
array[36314] <= 16'b0000_0000_0000_0000;
array[36315] <= 16'b0000_0000_0000_0000;
array[36316] <= 16'b0000_0000_0000_0000;
array[36317] <= 16'b0000_0000_0000_0000;
array[36318] <= 16'b0000_0000_0000_0000;
array[36319] <= 16'b0000_0000_0000_0000;
array[36320] <= 16'b0000_0000_0000_0000;
array[36321] <= 16'b0000_0000_0000_0000;
array[36322] <= 16'b0000_0000_0000_0000;
array[36323] <= 16'b0000_0000_0000_0000;
array[36324] <= 16'b0000_0000_0000_0000;
array[36325] <= 16'b0000_0000_0000_0000;
array[36326] <= 16'b0000_0000_0000_0000;
array[36327] <= 16'b0000_0000_0000_0000;
array[36328] <= 16'b0000_0000_0000_0000;
array[36329] <= 16'b0000_0000_0000_0000;
array[36330] <= 16'b0000_0000_0000_0000;
array[36331] <= 16'b0000_0000_0000_0000;
array[36332] <= 16'b0000_0000_0000_0000;
array[36333] <= 16'b0000_0000_0000_0000;
array[36334] <= 16'b0000_0000_0000_0000;
array[36335] <= 16'b0000_0000_0000_0000;
array[36336] <= 16'b0000_0000_0000_0000;
array[36337] <= 16'b0000_0000_0000_0000;
array[36338] <= 16'b0000_0000_0000_0000;
array[36339] <= 16'b0000_0000_0000_0000;
array[36340] <= 16'b0000_0000_0000_0000;
array[36341] <= 16'b0000_0000_0000_0000;
array[36342] <= 16'b0000_0000_0000_0000;
array[36343] <= 16'b0000_0000_0000_0000;
array[36344] <= 16'b0000_0000_0000_0000;
array[36345] <= 16'b0000_0000_0000_0000;
array[36346] <= 16'b0000_0000_0000_0000;
array[36347] <= 16'b0000_0000_0000_0000;
array[36348] <= 16'b0000_0000_0000_0000;
array[36349] <= 16'b0000_0000_0000_0000;
array[36350] <= 16'b0000_0000_0000_0000;
array[36351] <= 16'b0000_0000_0000_0000;
array[36352] <= 16'b0000_0000_0000_0000;
array[36353] <= 16'b0000_0000_0000_0000;
array[36354] <= 16'b0000_0000_0000_0000;
array[36355] <= 16'b0000_0000_0000_0000;
array[36356] <= 16'b0000_0000_0000_0000;
array[36357] <= 16'b0000_0000_0000_0000;
array[36358] <= 16'b0000_0000_0000_0000;
array[36359] <= 16'b0000_0000_0000_0000;
array[36360] <= 16'b0000_0000_0000_0000;
array[36361] <= 16'b0000_0000_0000_0000;
array[36362] <= 16'b0000_0000_0000_0000;
array[36363] <= 16'b0000_0000_0000_0000;
array[36364] <= 16'b0000_0000_0000_0000;
array[36365] <= 16'b0000_0000_0000_0000;
array[36366] <= 16'b0000_0000_0000_0000;
array[36367] <= 16'b0000_0000_0000_0000;
array[36368] <= 16'b0000_0000_0000_0000;
array[36369] <= 16'b0000_0000_0000_0000;
array[36370] <= 16'b0000_0000_0000_0000;
array[36371] <= 16'b0000_0000_0000_0000;
array[36372] <= 16'b0000_0000_0000_0000;
array[36373] <= 16'b0000_0000_0000_0000;
array[36374] <= 16'b0000_0000_0000_0000;
array[36375] <= 16'b0000_0000_0000_0000;
array[36376] <= 16'b0000_0000_0000_0000;
array[36377] <= 16'b0000_0000_0000_0000;
array[36378] <= 16'b0000_0000_0000_0000;
array[36379] <= 16'b0000_0000_0000_0000;
array[36380] <= 16'b0000_0000_0000_0000;
array[36381] <= 16'b0000_0000_0000_0000;
array[36382] <= 16'b0000_0000_0000_0000;
array[36383] <= 16'b0000_0000_0000_0000;
array[36384] <= 16'b0000_0000_0000_0000;
array[36385] <= 16'b0000_0000_0000_0000;
array[36386] <= 16'b0000_0000_0000_0000;
array[36387] <= 16'b0000_0000_0000_0000;
array[36388] <= 16'b0000_0000_0000_0000;
array[36389] <= 16'b0000_0000_0000_0000;
array[36390] <= 16'b0000_0000_0000_0000;
array[36391] <= 16'b0000_0000_0000_0000;
array[36392] <= 16'b0000_0000_0000_0000;
array[36393] <= 16'b0000_0000_0000_0000;
array[36394] <= 16'b0000_0000_0000_0000;
array[36395] <= 16'b0000_0000_0000_0000;
array[36396] <= 16'b0000_0000_0000_0000;
array[36397] <= 16'b0000_0000_0000_0000;
array[36398] <= 16'b0000_0000_0000_0000;
array[36399] <= 16'b0000_0000_0000_0000;
array[36400] <= 16'b0000_0000_0000_0000;
array[36401] <= 16'b0000_0000_0000_0000;
array[36402] <= 16'b0000_0000_0000_0000;
array[36403] <= 16'b0000_0000_0000_0000;
array[36404] <= 16'b0000_0000_0000_0000;
array[36405] <= 16'b0000_0000_0000_0000;
array[36406] <= 16'b0000_0000_0000_0000;
array[36407] <= 16'b0000_0000_0000_0000;
array[36408] <= 16'b0000_0000_0000_0000;
array[36409] <= 16'b0000_0000_0000_0000;
array[36410] <= 16'b0000_0000_0000_0000;
array[36411] <= 16'b0000_0000_0000_0000;
array[36412] <= 16'b0000_0000_0000_0000;
array[36413] <= 16'b0000_0000_0000_0000;
array[36414] <= 16'b0000_0000_0000_0000;
array[36415] <= 16'b0000_0000_0000_0000;
array[36416] <= 16'b0000_0000_0000_0000;
array[36417] <= 16'b0000_0000_0000_0000;
array[36418] <= 16'b0000_0000_0000_0000;
array[36419] <= 16'b0000_0000_0000_0000;
array[36420] <= 16'b0000_0000_0000_0000;
array[36421] <= 16'b0000_0000_0000_0000;
array[36422] <= 16'b0000_0000_0000_0000;
array[36423] <= 16'b0000_0000_0000_0000;
array[36424] <= 16'b0000_0000_0000_0000;
array[36425] <= 16'b0000_0000_0000_0000;
array[36426] <= 16'b0000_0000_0000_0000;
array[36427] <= 16'b0000_0000_0000_0000;
array[36428] <= 16'b0000_0000_0000_0000;
array[36429] <= 16'b0000_0000_0000_0000;
array[36430] <= 16'b0000_0000_0000_0000;
array[36431] <= 16'b0000_0000_0000_0000;
array[36432] <= 16'b0000_0000_0000_0000;
array[36433] <= 16'b0000_0000_0000_0000;
array[36434] <= 16'b0000_0000_0000_0000;
array[36435] <= 16'b0000_0000_0000_0000;
array[36436] <= 16'b0000_0000_0000_0000;
array[36437] <= 16'b0000_0000_0000_0000;
array[36438] <= 16'b0000_0000_0000_0000;
array[36439] <= 16'b0000_0000_0000_0000;
array[36440] <= 16'b0000_0000_0000_0000;
array[36441] <= 16'b0000_0000_0000_0000;
array[36442] <= 16'b0000_0000_0000_0000;
array[36443] <= 16'b0000_0000_0000_0000;
array[36444] <= 16'b0000_0000_0000_0000;
array[36445] <= 16'b0000_0000_0000_0000;
array[36446] <= 16'b0000_0000_0000_0000;
array[36447] <= 16'b0000_0000_0000_0000;
array[36448] <= 16'b0000_0000_0000_0000;
array[36449] <= 16'b0000_0000_0000_0000;
array[36450] <= 16'b0000_0000_0000_0000;
array[36451] <= 16'b0000_0000_0000_0000;
array[36452] <= 16'b0000_0000_0000_0000;
array[36453] <= 16'b0000_0000_0000_0000;
array[36454] <= 16'b0000_0000_0000_0000;
array[36455] <= 16'b0000_0000_0000_0000;
array[36456] <= 16'b0000_0000_0000_0000;
array[36457] <= 16'b0000_0000_0000_0000;
array[36458] <= 16'b0000_0000_0000_0000;
array[36459] <= 16'b0000_0000_0000_0000;
array[36460] <= 16'b0000_0000_0000_0000;
array[36461] <= 16'b0000_0000_0000_0000;
array[36462] <= 16'b0000_0000_0000_0000;
array[36463] <= 16'b0000_0000_0000_0000;
array[36464] <= 16'b0000_0000_0000_0000;
array[36465] <= 16'b0000_0000_0000_0000;
array[36466] <= 16'b0000_0000_0000_0000;
array[36467] <= 16'b0000_0000_0000_0000;
array[36468] <= 16'b0000_0000_0000_0000;
array[36469] <= 16'b0000_0000_0000_0000;
array[36470] <= 16'b0000_0000_0000_0000;
array[36471] <= 16'b0000_0000_0000_0000;
array[36472] <= 16'b0000_0000_0000_0000;
array[36473] <= 16'b0000_0000_0000_0000;
array[36474] <= 16'b0000_0000_0000_0000;
array[36475] <= 16'b0000_0000_0000_0000;
array[36476] <= 16'b0000_0000_0000_0000;
array[36477] <= 16'b0000_0000_0000_0000;
array[36478] <= 16'b0000_0000_0000_0000;
array[36479] <= 16'b0000_0000_0000_0000;
array[36480] <= 16'b0000_0000_0000_0000;
array[36481] <= 16'b0000_0000_0000_0000;
array[36482] <= 16'b0000_0000_0000_0000;
array[36483] <= 16'b0000_0000_0000_0000;
array[36484] <= 16'b0000_0000_0000_0000;
array[36485] <= 16'b0000_0000_0000_0000;
array[36486] <= 16'b0000_0000_0000_0000;
array[36487] <= 16'b0000_0000_0000_0000;
array[36488] <= 16'b0000_0000_0000_0000;
array[36489] <= 16'b0000_0000_0000_0000;
array[36490] <= 16'b0000_0000_0000_0000;
array[36491] <= 16'b0000_0000_0000_0000;
array[36492] <= 16'b0000_0000_0000_0000;
array[36493] <= 16'b0000_0000_0000_0000;
array[36494] <= 16'b0000_0000_0000_0000;
array[36495] <= 16'b0000_0000_0000_0000;
array[36496] <= 16'b0000_0000_0000_0000;
array[36497] <= 16'b0000_0000_0000_0000;
array[36498] <= 16'b0000_0000_0000_0000;
array[36499] <= 16'b0000_0000_0000_0000;
array[36500] <= 16'b0000_0000_0000_0000;
array[36501] <= 16'b0000_0000_0000_0000;
array[36502] <= 16'b0000_0000_0000_0000;
array[36503] <= 16'b0000_0000_0000_0000;
array[36504] <= 16'b0000_0000_0000_0000;
array[36505] <= 16'b0000_0000_0000_0000;
array[36506] <= 16'b0000_0000_0000_0000;
array[36507] <= 16'b0000_0000_0000_0000;
array[36508] <= 16'b0000_0000_0000_0000;
array[36509] <= 16'b0000_0000_0000_0000;
array[36510] <= 16'b0000_0000_0000_0000;
array[36511] <= 16'b0000_0000_0000_0000;
array[36512] <= 16'b0000_0000_0000_0000;
array[36513] <= 16'b0000_0000_0000_0000;
array[36514] <= 16'b0000_0000_0000_0000;
array[36515] <= 16'b0000_0000_0000_0000;
array[36516] <= 16'b0000_0000_0000_0000;
array[36517] <= 16'b0000_0000_0000_0000;
array[36518] <= 16'b0000_0000_0000_0000;
array[36519] <= 16'b0000_0000_0000_0000;
array[36520] <= 16'b0000_0000_0000_0000;
array[36521] <= 16'b0000_0000_0000_0000;
array[36522] <= 16'b0000_0000_0000_0000;
array[36523] <= 16'b0000_0000_0000_0000;
array[36524] <= 16'b0000_0000_0000_0000;
array[36525] <= 16'b0000_0000_0000_0000;
array[36526] <= 16'b0000_0000_0000_0000;
array[36527] <= 16'b0000_0000_0000_0000;
array[36528] <= 16'b0000_0000_0000_0000;
array[36529] <= 16'b0000_0000_0000_0000;
array[36530] <= 16'b0000_0000_0000_0000;
array[36531] <= 16'b0000_0000_0000_0000;
array[36532] <= 16'b0000_0000_0000_0000;
array[36533] <= 16'b0000_0000_0000_0000;
array[36534] <= 16'b0000_0000_0000_0000;
array[36535] <= 16'b0000_0000_0000_0000;
array[36536] <= 16'b0000_0000_0000_0000;
array[36537] <= 16'b0000_0000_0000_0000;
array[36538] <= 16'b0000_0000_0000_0000;
array[36539] <= 16'b0000_0000_0000_0000;
array[36540] <= 16'b0000_0000_0000_0000;
array[36541] <= 16'b0000_0000_0000_0000;
array[36542] <= 16'b0000_0000_0000_0000;
array[36543] <= 16'b0000_0000_0000_0000;
array[36544] <= 16'b0000_0000_0000_0000;
array[36545] <= 16'b0000_0000_0000_0000;
array[36546] <= 16'b0000_0000_0000_0000;
array[36547] <= 16'b0000_0000_0000_0000;
array[36548] <= 16'b0000_0000_0000_0000;
array[36549] <= 16'b0000_0000_0000_0000;
array[36550] <= 16'b0000_0000_0000_0000;
array[36551] <= 16'b0000_0000_0000_0000;
array[36552] <= 16'b0000_0000_0000_0000;
array[36553] <= 16'b0000_0000_0000_0000;
array[36554] <= 16'b0000_0000_0000_0000;
array[36555] <= 16'b0000_0000_0000_0000;
array[36556] <= 16'b0000_0000_0000_0000;
array[36557] <= 16'b0000_0000_0000_0000;
array[36558] <= 16'b0000_0000_0000_0000;
array[36559] <= 16'b0000_0000_0000_0000;
array[36560] <= 16'b0000_0000_0000_0000;
array[36561] <= 16'b0000_0000_0000_0000;
array[36562] <= 16'b0000_0000_0000_0000;
array[36563] <= 16'b0000_0000_0000_0000;
array[36564] <= 16'b0000_0000_0000_0000;
array[36565] <= 16'b0000_0000_0000_0000;
array[36566] <= 16'b0000_0000_0000_0000;
array[36567] <= 16'b0000_0000_0000_0000;
array[36568] <= 16'b0000_0000_0000_0000;
array[36569] <= 16'b0000_0000_0000_0000;
array[36570] <= 16'b0000_0000_0000_0000;
array[36571] <= 16'b0000_0000_0000_0000;
array[36572] <= 16'b0000_0000_0000_0000;
array[36573] <= 16'b0000_0000_0000_0000;
array[36574] <= 16'b0000_0000_0000_0000;
array[36575] <= 16'b0000_0000_0000_0000;
array[36576] <= 16'b0000_0000_0000_0000;
array[36577] <= 16'b0000_0000_0000_0000;
array[36578] <= 16'b0000_0000_0000_0000;
array[36579] <= 16'b0000_0000_0000_0000;
array[36580] <= 16'b0000_0000_0000_0000;
array[36581] <= 16'b0000_0000_0000_0000;
array[36582] <= 16'b0000_0000_0000_0000;
array[36583] <= 16'b0000_0000_0000_0000;
array[36584] <= 16'b0000_0000_0000_0000;
array[36585] <= 16'b0000_0000_0000_0000;
array[36586] <= 16'b0000_0000_0000_0000;
array[36587] <= 16'b0000_0000_0000_0000;
array[36588] <= 16'b0000_0000_0000_0000;
array[36589] <= 16'b0000_0000_0000_0000;
array[36590] <= 16'b0000_0000_0000_0000;
array[36591] <= 16'b0000_0000_0000_0000;
array[36592] <= 16'b0000_0000_0000_0000;
array[36593] <= 16'b0000_0000_0000_0000;
array[36594] <= 16'b0000_0000_0000_0000;
array[36595] <= 16'b0000_0000_0000_0000;
array[36596] <= 16'b0000_0000_0000_0000;
array[36597] <= 16'b0000_0000_0000_0000;
array[36598] <= 16'b0000_0000_0000_0000;
array[36599] <= 16'b0000_0000_0000_0000;
array[36600] <= 16'b0000_0000_0000_0000;
array[36601] <= 16'b0000_0000_0000_0000;
array[36602] <= 16'b0000_0000_0000_0000;
array[36603] <= 16'b0000_0000_0000_0000;
array[36604] <= 16'b0000_0000_0000_0000;
array[36605] <= 16'b0000_0000_0000_0000;
array[36606] <= 16'b0000_0000_0000_0000;
array[36607] <= 16'b0000_0000_0000_0000;
array[36608] <= 16'b0000_0000_0000_0000;
array[36609] <= 16'b0000_0000_0000_0000;
array[36610] <= 16'b0000_0000_0000_0000;
array[36611] <= 16'b0000_0000_0000_0000;
array[36612] <= 16'b0000_0000_0000_0000;
array[36613] <= 16'b0000_0000_0000_0000;
array[36614] <= 16'b0000_0000_0000_0000;
array[36615] <= 16'b0000_0000_0000_0000;
array[36616] <= 16'b0000_0000_0000_0000;
array[36617] <= 16'b0000_0000_0000_0000;
array[36618] <= 16'b0000_0000_0000_0000;
array[36619] <= 16'b0000_0000_0000_0000;
array[36620] <= 16'b0000_0000_0000_0000;
array[36621] <= 16'b0000_0000_0000_0000;
array[36622] <= 16'b0000_0000_0000_0000;
array[36623] <= 16'b0000_0000_0000_0000;
array[36624] <= 16'b0000_0000_0000_0000;
array[36625] <= 16'b0000_0000_0000_0000;
array[36626] <= 16'b0000_0000_0000_0000;
array[36627] <= 16'b0000_0000_0000_0000;
array[36628] <= 16'b0000_0000_0000_0000;
array[36629] <= 16'b0000_0000_0000_0000;
array[36630] <= 16'b0000_0000_0000_0000;
array[36631] <= 16'b0000_0000_0000_0000;
array[36632] <= 16'b0000_0000_0000_0000;
array[36633] <= 16'b0000_0000_0000_0000;
array[36634] <= 16'b0000_0000_0000_0000;
array[36635] <= 16'b0000_0000_0000_0000;
array[36636] <= 16'b0000_0000_0000_0000;
array[36637] <= 16'b0000_0000_0000_0000;
array[36638] <= 16'b0000_0000_0000_0000;
array[36639] <= 16'b0000_0000_0000_0000;
array[36640] <= 16'b0000_0000_0000_0000;
array[36641] <= 16'b0000_0000_0000_0000;
array[36642] <= 16'b0000_0000_0000_0000;
array[36643] <= 16'b0000_0000_0000_0000;
array[36644] <= 16'b0000_0000_0000_0000;
array[36645] <= 16'b0000_0000_0000_0000;
array[36646] <= 16'b0000_0000_0000_0000;
array[36647] <= 16'b0000_0000_0000_0000;
array[36648] <= 16'b0000_0000_0000_0000;
array[36649] <= 16'b0000_0000_0000_0000;
array[36650] <= 16'b0000_0000_0000_0000;
array[36651] <= 16'b0000_0000_0000_0000;
array[36652] <= 16'b0000_0000_0000_0000;
array[36653] <= 16'b0000_0000_0000_0000;
array[36654] <= 16'b0000_0000_0000_0000;
array[36655] <= 16'b0000_0000_0000_0000;
array[36656] <= 16'b0000_0000_0000_0000;
array[36657] <= 16'b0000_0000_0000_0000;
array[36658] <= 16'b0000_0000_0000_0000;
array[36659] <= 16'b0000_0000_0000_0000;
array[36660] <= 16'b0000_0000_0000_0000;
array[36661] <= 16'b0000_0000_0000_0000;
array[36662] <= 16'b0000_0000_0000_0000;
array[36663] <= 16'b0000_0000_0000_0000;
array[36664] <= 16'b0000_0000_0000_0000;
array[36665] <= 16'b0000_0000_0000_0000;
array[36666] <= 16'b0000_0000_0000_0000;
array[36667] <= 16'b0000_0000_0000_0000;
array[36668] <= 16'b0000_0000_0000_0000;
array[36669] <= 16'b0000_0000_0000_0000;
array[36670] <= 16'b0000_0000_0000_0000;
array[36671] <= 16'b0000_0000_0000_0000;
array[36672] <= 16'b0000_0000_0000_0000;
array[36673] <= 16'b0000_0000_0000_0000;
array[36674] <= 16'b0000_0000_0000_0000;
array[36675] <= 16'b0000_0000_0000_0000;
array[36676] <= 16'b0000_0000_0000_0000;
array[36677] <= 16'b0000_0000_0000_0000;
array[36678] <= 16'b0000_0000_0000_0000;
array[36679] <= 16'b0000_0000_0000_0000;
array[36680] <= 16'b0000_0000_0000_0000;
array[36681] <= 16'b0000_0000_0000_0000;
array[36682] <= 16'b0000_0000_0000_0000;
array[36683] <= 16'b0000_0000_0000_0000;
array[36684] <= 16'b0000_0000_0000_0000;
array[36685] <= 16'b0000_0000_0000_0000;
array[36686] <= 16'b0000_0000_0000_0000;
array[36687] <= 16'b0000_0000_0000_0000;
array[36688] <= 16'b0000_0000_0000_0000;
array[36689] <= 16'b0000_0000_0000_0000;
array[36690] <= 16'b0000_0000_0000_0000;
array[36691] <= 16'b0000_0000_0000_0000;
array[36692] <= 16'b0000_0000_0000_0000;
array[36693] <= 16'b0000_0000_0000_0000;
array[36694] <= 16'b0000_0000_0000_0000;
array[36695] <= 16'b0000_0000_0000_0000;
array[36696] <= 16'b0000_0000_0000_0000;
array[36697] <= 16'b0000_0000_0000_0000;
array[36698] <= 16'b0000_0000_0000_0000;
array[36699] <= 16'b0000_0000_0000_0000;
array[36700] <= 16'b0000_0000_0000_0000;
array[36701] <= 16'b0000_0000_0000_0000;
array[36702] <= 16'b0000_0000_0000_0000;
array[36703] <= 16'b0000_0000_0000_0000;
array[36704] <= 16'b0000_0000_0000_0000;
array[36705] <= 16'b0000_0000_0000_0000;
array[36706] <= 16'b0000_0000_0000_0000;
array[36707] <= 16'b0000_0000_0000_0000;
array[36708] <= 16'b0000_0000_0000_0000;
array[36709] <= 16'b0000_0000_0000_0000;
array[36710] <= 16'b0000_0000_0000_0000;
array[36711] <= 16'b0000_0000_0000_0000;
array[36712] <= 16'b0000_0000_0000_0000;
array[36713] <= 16'b0000_0000_0000_0000;
array[36714] <= 16'b0000_0000_0000_0000;
array[36715] <= 16'b0000_0000_0000_0000;
array[36716] <= 16'b0000_0000_0000_0000;
array[36717] <= 16'b0000_0000_0000_0000;
array[36718] <= 16'b0000_0000_0000_0000;
array[36719] <= 16'b0000_0000_0000_0000;
array[36720] <= 16'b0000_0000_0000_0000;
array[36721] <= 16'b0000_0000_0000_0000;
array[36722] <= 16'b0000_0000_0000_0000;
array[36723] <= 16'b0000_0000_0000_0000;
array[36724] <= 16'b0000_0000_0000_0000;
array[36725] <= 16'b0000_0000_0000_0000;
array[36726] <= 16'b0000_0000_0000_0000;
array[36727] <= 16'b0000_0000_0000_0000;
array[36728] <= 16'b0000_0000_0000_0000;
array[36729] <= 16'b0000_0000_0000_0000;
array[36730] <= 16'b0000_0000_0000_0000;
array[36731] <= 16'b0000_0000_0000_0000;
array[36732] <= 16'b0000_0000_0000_0000;
array[36733] <= 16'b0000_0000_0000_0000;
array[36734] <= 16'b0000_0000_0000_0000;
array[36735] <= 16'b0000_0000_0000_0000;
array[36736] <= 16'b0000_0000_0000_0000;
array[36737] <= 16'b0000_0000_0000_0000;
array[36738] <= 16'b0000_0000_0000_0000;
array[36739] <= 16'b0000_0000_0000_0000;
array[36740] <= 16'b0000_0000_0000_0000;
array[36741] <= 16'b0000_0000_0000_0000;
array[36742] <= 16'b0000_0000_0000_0000;
array[36743] <= 16'b0000_0000_0000_0000;
array[36744] <= 16'b0000_0000_0000_0000;
array[36745] <= 16'b0000_0000_0000_0000;
array[36746] <= 16'b0000_0000_0000_0000;
array[36747] <= 16'b0000_0000_0000_0000;
array[36748] <= 16'b0000_0000_0000_0000;
array[36749] <= 16'b0000_0000_0000_0000;
array[36750] <= 16'b0000_0000_0000_0000;
array[36751] <= 16'b0000_0000_0000_0000;
array[36752] <= 16'b0000_0000_0000_0000;
array[36753] <= 16'b0000_0000_0000_0000;
array[36754] <= 16'b0000_0000_0000_0000;
array[36755] <= 16'b0000_0000_0000_0000;
array[36756] <= 16'b0000_0000_0000_0000;
array[36757] <= 16'b0000_0000_0000_0000;
array[36758] <= 16'b0000_0000_0000_0000;
array[36759] <= 16'b0000_0000_0000_0000;
array[36760] <= 16'b0000_0000_0000_0000;
array[36761] <= 16'b0000_0000_0000_0000;
array[36762] <= 16'b0000_0000_0000_0000;
array[36763] <= 16'b0000_0000_0000_0000;
array[36764] <= 16'b0000_0000_0000_0000;
array[36765] <= 16'b0000_0000_0000_0000;
array[36766] <= 16'b0000_0000_0000_0000;
array[36767] <= 16'b0000_0000_0000_0000;
array[36768] <= 16'b0000_0000_0000_0000;
array[36769] <= 16'b0000_0000_0000_0000;
array[36770] <= 16'b0000_0000_0000_0000;
array[36771] <= 16'b0000_0000_0000_0000;
array[36772] <= 16'b0000_0000_0000_0000;
array[36773] <= 16'b0000_0000_0000_0000;
array[36774] <= 16'b0000_0000_0000_0000;
array[36775] <= 16'b0000_0000_0000_0000;
array[36776] <= 16'b0000_0000_0000_0000;
array[36777] <= 16'b0000_0000_0000_0000;
array[36778] <= 16'b0000_0000_0000_0000;
array[36779] <= 16'b0000_0000_0000_0000;
array[36780] <= 16'b0000_0000_0000_0000;
array[36781] <= 16'b0000_0000_0000_0000;
array[36782] <= 16'b0000_0000_0000_0000;
array[36783] <= 16'b0000_0000_0000_0000;
array[36784] <= 16'b0000_0000_0000_0000;
array[36785] <= 16'b0000_0000_0000_0000;
array[36786] <= 16'b0000_0000_0000_0000;
array[36787] <= 16'b0000_0000_0000_0000;
array[36788] <= 16'b0000_0000_0000_0000;
array[36789] <= 16'b0000_0000_0000_0000;
array[36790] <= 16'b0000_0000_0000_0000;
array[36791] <= 16'b0000_0000_0000_0000;
array[36792] <= 16'b0000_0000_0000_0000;
array[36793] <= 16'b0000_0000_0000_0000;
array[36794] <= 16'b0000_0000_0000_0000;
array[36795] <= 16'b0000_0000_0000_0000;
array[36796] <= 16'b0000_0000_0000_0000;
array[36797] <= 16'b0000_0000_0000_0000;
array[36798] <= 16'b0000_0000_0000_0000;
array[36799] <= 16'b0000_0000_0000_0000;
array[36800] <= 16'b0000_0000_0000_0000;
array[36801] <= 16'b0000_0000_0000_0000;
array[36802] <= 16'b0000_0000_0000_0000;
array[36803] <= 16'b0000_0000_0000_0000;
array[36804] <= 16'b0000_0000_0000_0000;
array[36805] <= 16'b0000_0000_0000_0000;
array[36806] <= 16'b0000_0000_0000_0000;
array[36807] <= 16'b0000_0000_0000_0000;
array[36808] <= 16'b0000_0000_0000_0000;
array[36809] <= 16'b0000_0000_0000_0000;
array[36810] <= 16'b0000_0000_0000_0000;
array[36811] <= 16'b0000_0000_0000_0000;
array[36812] <= 16'b0000_0000_0000_0000;
array[36813] <= 16'b0000_0000_0000_0000;
array[36814] <= 16'b0000_0000_0000_0000;
array[36815] <= 16'b0000_0000_0000_0000;
array[36816] <= 16'b0000_0000_0000_0000;
array[36817] <= 16'b0000_0000_0000_0000;
array[36818] <= 16'b0000_0000_0000_0000;
array[36819] <= 16'b0000_0000_0000_0000;
array[36820] <= 16'b0000_0000_0000_0000;
array[36821] <= 16'b0000_0000_0000_0000;
array[36822] <= 16'b0000_0000_0000_0000;
array[36823] <= 16'b0000_0000_0000_0000;
array[36824] <= 16'b0000_0000_0000_0000;
array[36825] <= 16'b0000_0000_0000_0000;
array[36826] <= 16'b0000_0000_0000_0000;
array[36827] <= 16'b0000_0000_0000_0000;
array[36828] <= 16'b0000_0000_0000_0000;
array[36829] <= 16'b0000_0000_0000_0000;
array[36830] <= 16'b0000_0000_0000_0000;
array[36831] <= 16'b0000_0000_0000_0000;
array[36832] <= 16'b0000_0000_0000_0000;
array[36833] <= 16'b0000_0000_0000_0000;
array[36834] <= 16'b0000_0000_0000_0000;
array[36835] <= 16'b0000_0000_0000_0000;
array[36836] <= 16'b0000_0000_0000_0000;
array[36837] <= 16'b0000_0000_0000_0000;
array[36838] <= 16'b0000_0000_0000_0000;
array[36839] <= 16'b0000_0000_0000_0000;
array[36840] <= 16'b0000_0000_0000_0000;
array[36841] <= 16'b0000_0000_0000_0000;
array[36842] <= 16'b0000_0000_0000_0000;
array[36843] <= 16'b0000_0000_0000_0000;
array[36844] <= 16'b0000_0000_0000_0000;
array[36845] <= 16'b0000_0000_0000_0000;
array[36846] <= 16'b0000_0000_0000_0000;
array[36847] <= 16'b0000_0000_0000_0000;
array[36848] <= 16'b0000_0000_0000_0000;
array[36849] <= 16'b0000_0000_0000_0000;
array[36850] <= 16'b0000_0000_0000_0000;
array[36851] <= 16'b0000_0000_0000_0000;
array[36852] <= 16'b0000_0000_0000_0000;
array[36853] <= 16'b0000_0000_0000_0000;
array[36854] <= 16'b0000_0000_0000_0000;
array[36855] <= 16'b0000_0000_0000_0000;
array[36856] <= 16'b0000_0000_0000_0000;
array[36857] <= 16'b0000_0000_0000_0000;
array[36858] <= 16'b0000_0000_0000_0000;
array[36859] <= 16'b0000_0000_0000_0000;
array[36860] <= 16'b0000_0000_0000_0000;
array[36861] <= 16'b0000_0000_0000_0000;
array[36862] <= 16'b0000_0000_0000_0000;
array[36863] <= 16'b0000_0000_0000_0000;
array[36864] <= 16'b0000_0000_0000_0000;
array[36865] <= 16'b0000_0000_0000_0000;
array[36866] <= 16'b0000_0000_0000_0000;
array[36867] <= 16'b0000_0000_0000_0000;
array[36868] <= 16'b0000_0000_0000_0000;
array[36869] <= 16'b0000_0000_0000_0000;
array[36870] <= 16'b0000_0000_0000_0000;
array[36871] <= 16'b0000_0000_0000_0000;
array[36872] <= 16'b0000_0000_0000_0000;
array[36873] <= 16'b0000_0000_0000_0000;
array[36874] <= 16'b0000_0000_0000_0000;
array[36875] <= 16'b0000_0000_0000_0000;
array[36876] <= 16'b0000_0000_0000_0000;
array[36877] <= 16'b0000_0000_0000_0000;
array[36878] <= 16'b0000_0000_0000_0000;
array[36879] <= 16'b0000_0000_0000_0000;
array[36880] <= 16'b0000_0000_0000_0000;
array[36881] <= 16'b0000_0000_0000_0000;
array[36882] <= 16'b0000_0000_0000_0000;
array[36883] <= 16'b0000_0000_0000_0000;
array[36884] <= 16'b0000_0000_0000_0000;
array[36885] <= 16'b0000_0000_0000_0000;
array[36886] <= 16'b0000_0000_0000_0000;
array[36887] <= 16'b0000_0000_0000_0000;
array[36888] <= 16'b0000_0000_0000_0000;
array[36889] <= 16'b0000_0000_0000_0000;
array[36890] <= 16'b0000_0000_0000_0000;
array[36891] <= 16'b0000_0000_0000_0000;
array[36892] <= 16'b0000_0000_0000_0000;
array[36893] <= 16'b0000_0000_0000_0000;
array[36894] <= 16'b0000_0000_0000_0000;
array[36895] <= 16'b0000_0000_0000_0000;
array[36896] <= 16'b0000_0000_0000_0000;
array[36897] <= 16'b0000_0000_0000_0000;
array[36898] <= 16'b0000_0000_0000_0000;
array[36899] <= 16'b0000_0000_0000_0000;
array[36900] <= 16'b0000_0000_0000_0000;
array[36901] <= 16'b0000_0000_0000_0000;
array[36902] <= 16'b0000_0000_0000_0000;
array[36903] <= 16'b0000_0000_0000_0000;
array[36904] <= 16'b0000_0000_0000_0000;
array[36905] <= 16'b0000_0000_0000_0000;
array[36906] <= 16'b0000_0000_0000_0000;
array[36907] <= 16'b0000_0000_0000_0000;
array[36908] <= 16'b0000_0000_0000_0000;
array[36909] <= 16'b0000_0000_0000_0000;
array[36910] <= 16'b0000_0000_0000_0000;
array[36911] <= 16'b0000_0000_0000_0000;
array[36912] <= 16'b0000_0000_0000_0000;
array[36913] <= 16'b0000_0000_0000_0000;
array[36914] <= 16'b0000_0000_0000_0000;
array[36915] <= 16'b0000_0000_0000_0000;
array[36916] <= 16'b0000_0000_0000_0000;
array[36917] <= 16'b0000_0000_0000_0000;
array[36918] <= 16'b0000_0000_0000_0000;
array[36919] <= 16'b0000_0000_0000_0000;
array[36920] <= 16'b0000_0000_0000_0000;
array[36921] <= 16'b0000_0000_0000_0000;
array[36922] <= 16'b0000_0000_0000_0000;
array[36923] <= 16'b0000_0000_0000_0000;
array[36924] <= 16'b0000_0000_0000_0000;
array[36925] <= 16'b0000_0000_0000_0000;
array[36926] <= 16'b0000_0000_0000_0000;
array[36927] <= 16'b0000_0000_0000_0000;
array[36928] <= 16'b0000_0000_0000_0000;
array[36929] <= 16'b0000_0000_0000_0000;
array[36930] <= 16'b0000_0000_0000_0000;
array[36931] <= 16'b0000_0000_0000_0000;
array[36932] <= 16'b0000_0000_0000_0000;
array[36933] <= 16'b0000_0000_0000_0000;
array[36934] <= 16'b0000_0000_0000_0000;
array[36935] <= 16'b0000_0000_0000_0000;
array[36936] <= 16'b0000_0000_0000_0000;
array[36937] <= 16'b0000_0000_0000_0000;
array[36938] <= 16'b0000_0000_0000_0000;
array[36939] <= 16'b0000_0000_0000_0000;
array[36940] <= 16'b0000_0000_0000_0000;
array[36941] <= 16'b0000_0000_0000_0000;
array[36942] <= 16'b0000_0000_0000_0000;
array[36943] <= 16'b0000_0000_0000_0000;
array[36944] <= 16'b0000_0000_0000_0000;
array[36945] <= 16'b0000_0000_0000_0000;
array[36946] <= 16'b0000_0000_0000_0000;
array[36947] <= 16'b0000_0000_0000_0000;
array[36948] <= 16'b0000_0000_0000_0000;
array[36949] <= 16'b0000_0000_0000_0000;
array[36950] <= 16'b0000_0000_0000_0000;
array[36951] <= 16'b0000_0000_0000_0000;
array[36952] <= 16'b0000_0000_0000_0000;
array[36953] <= 16'b0000_0000_0000_0000;
array[36954] <= 16'b0000_0000_0000_0000;
array[36955] <= 16'b0000_0000_0000_0000;
array[36956] <= 16'b0000_0000_0000_0000;
array[36957] <= 16'b0000_0000_0000_0000;
array[36958] <= 16'b0000_0000_0000_0000;
array[36959] <= 16'b0000_0000_0000_0000;
array[36960] <= 16'b0000_0000_0000_0000;
array[36961] <= 16'b0000_0000_0000_0000;
array[36962] <= 16'b0000_0000_0000_0000;
array[36963] <= 16'b0000_0000_0000_0000;
array[36964] <= 16'b0000_0000_0000_0000;
array[36965] <= 16'b0000_0000_0000_0000;
array[36966] <= 16'b0000_0000_0000_0000;
array[36967] <= 16'b0000_0000_0000_0000;
array[36968] <= 16'b0000_0000_0000_0000;
array[36969] <= 16'b0000_0000_0000_0000;
array[36970] <= 16'b0000_0000_0000_0000;
array[36971] <= 16'b0000_0000_0000_0000;
array[36972] <= 16'b0000_0000_0000_0000;
array[36973] <= 16'b0000_0000_0000_0000;
array[36974] <= 16'b0000_0000_0000_0000;
array[36975] <= 16'b0000_0000_0000_0000;
array[36976] <= 16'b0000_0000_0000_0000;
array[36977] <= 16'b0000_0000_0000_0000;
array[36978] <= 16'b0000_0000_0000_0000;
array[36979] <= 16'b0000_0000_0000_0000;
array[36980] <= 16'b0000_0000_0000_0000;
array[36981] <= 16'b0000_0000_0000_0000;
array[36982] <= 16'b0000_0000_0000_0000;
array[36983] <= 16'b0000_0000_0000_0000;
array[36984] <= 16'b0000_0000_0000_0000;
array[36985] <= 16'b0000_0000_0000_0000;
array[36986] <= 16'b0000_0000_0000_0000;
array[36987] <= 16'b0000_0000_0000_0000;
array[36988] <= 16'b0000_0000_0000_0000;
array[36989] <= 16'b0000_0000_0000_0000;
array[36990] <= 16'b0000_0000_0000_0000;
array[36991] <= 16'b0000_0000_0000_0000;
array[36992] <= 16'b0000_0000_0000_0000;
array[36993] <= 16'b0000_0000_0000_0000;
array[36994] <= 16'b0000_0000_0000_0000;
array[36995] <= 16'b0000_0000_0000_0000;
array[36996] <= 16'b0000_0000_0000_0000;
array[36997] <= 16'b0000_0000_0000_0000;
array[36998] <= 16'b0000_0000_0000_0000;
array[36999] <= 16'b0000_0000_0000_0000;
array[37000] <= 16'b0000_0000_0000_0000;
array[37001] <= 16'b0000_0000_0000_0000;
array[37002] <= 16'b0000_0000_0000_0000;
array[37003] <= 16'b0000_0000_0000_0000;
array[37004] <= 16'b0000_0000_0000_0000;
array[37005] <= 16'b0000_0000_0000_0000;
array[37006] <= 16'b0000_0000_0000_0000;
array[37007] <= 16'b0000_0000_0000_0000;
array[37008] <= 16'b0000_0000_0000_0000;
array[37009] <= 16'b0000_0000_0000_0000;
array[37010] <= 16'b0000_0000_0000_0000;
array[37011] <= 16'b0000_0000_0000_0000;
array[37012] <= 16'b0000_0000_0000_0000;
array[37013] <= 16'b0000_0000_0000_0000;
array[37014] <= 16'b0000_0000_0000_0000;
array[37015] <= 16'b0000_0000_0000_0000;
array[37016] <= 16'b0000_0000_0000_0000;
array[37017] <= 16'b0000_0000_0000_0000;
array[37018] <= 16'b0000_0000_0000_0000;
array[37019] <= 16'b0000_0000_0000_0000;
array[37020] <= 16'b0000_0000_0000_0000;
array[37021] <= 16'b0000_0000_0000_0000;
array[37022] <= 16'b0000_0000_0000_0000;
array[37023] <= 16'b0000_0000_0000_0000;
array[37024] <= 16'b0000_0000_0000_0000;
array[37025] <= 16'b0000_0000_0000_0000;
array[37026] <= 16'b0000_0000_0000_0000;
array[37027] <= 16'b0000_0000_0000_0000;
array[37028] <= 16'b0000_0000_0000_0000;
array[37029] <= 16'b0000_0000_0000_0000;
array[37030] <= 16'b0000_0000_0000_0000;
array[37031] <= 16'b0000_0000_0000_0000;
array[37032] <= 16'b0000_0000_0000_0000;
array[37033] <= 16'b0000_0000_0000_0000;
array[37034] <= 16'b0000_0000_0000_0000;
array[37035] <= 16'b0000_0000_0000_0000;
array[37036] <= 16'b0000_0000_0000_0000;
array[37037] <= 16'b0000_0000_0000_0000;
array[37038] <= 16'b0000_0000_0000_0000;
array[37039] <= 16'b0000_0000_0000_0000;
array[37040] <= 16'b0000_0000_0000_0000;
array[37041] <= 16'b0000_0000_0000_0000;
array[37042] <= 16'b0000_0000_0000_0000;
array[37043] <= 16'b0000_0000_0000_0000;
array[37044] <= 16'b0000_0000_0000_0000;
array[37045] <= 16'b0000_0000_0000_0000;
array[37046] <= 16'b0000_0000_0000_0000;
array[37047] <= 16'b0000_0000_0000_0000;
array[37048] <= 16'b0000_0000_0000_0000;
array[37049] <= 16'b0000_0000_0000_0000;
array[37050] <= 16'b0000_0000_0000_0000;
array[37051] <= 16'b0000_0000_0000_0000;
array[37052] <= 16'b0000_0000_0000_0000;
array[37053] <= 16'b0000_0000_0000_0000;
array[37054] <= 16'b0000_0000_0000_0000;
array[37055] <= 16'b0000_0000_0000_0000;
array[37056] <= 16'b0000_0000_0000_0000;
array[37057] <= 16'b0000_0000_0000_0000;
array[37058] <= 16'b0000_0000_0000_0000;
array[37059] <= 16'b0000_0000_0000_0000;
array[37060] <= 16'b0000_0000_0000_0000;
array[37061] <= 16'b0000_0000_0000_0000;
array[37062] <= 16'b0000_0000_0000_0000;
array[37063] <= 16'b0000_0000_0000_0000;
array[37064] <= 16'b0000_0000_0000_0000;
array[37065] <= 16'b0000_0000_0000_0000;
array[37066] <= 16'b0000_0000_0000_0000;
array[37067] <= 16'b0000_0000_0000_0000;
array[37068] <= 16'b0000_0000_0000_0000;
array[37069] <= 16'b0000_0000_0000_0000;
array[37070] <= 16'b0000_0000_0000_0000;
array[37071] <= 16'b0000_0000_0000_0000;
array[37072] <= 16'b0000_0000_0000_0000;
array[37073] <= 16'b0000_0000_0000_0000;
array[37074] <= 16'b0000_0000_0000_0000;
array[37075] <= 16'b0000_0000_0000_0000;
array[37076] <= 16'b0000_0000_0000_0000;
array[37077] <= 16'b0000_0000_0000_0000;
array[37078] <= 16'b0000_0000_0000_0000;
array[37079] <= 16'b0000_0000_0000_0000;
array[37080] <= 16'b0000_0000_0000_0000;
array[37081] <= 16'b0000_0000_0000_0000;
array[37082] <= 16'b0000_0000_0000_0000;
array[37083] <= 16'b0000_0000_0000_0000;
array[37084] <= 16'b0000_0000_0000_0000;
array[37085] <= 16'b0000_0000_0000_0000;
array[37086] <= 16'b0000_0000_0000_0000;
array[37087] <= 16'b0000_0000_0000_0000;
array[37088] <= 16'b0000_0000_0000_0000;
array[37089] <= 16'b0000_0000_0000_0000;
array[37090] <= 16'b0000_0000_0000_0000;
array[37091] <= 16'b0000_0000_0000_0000;
array[37092] <= 16'b0000_0000_0000_0000;
array[37093] <= 16'b0000_0000_0000_0000;
array[37094] <= 16'b0000_0000_0000_0000;
array[37095] <= 16'b0000_0000_0000_0000;
array[37096] <= 16'b0000_0000_0000_0000;
array[37097] <= 16'b0000_0000_0000_0000;
array[37098] <= 16'b0000_0000_0000_0000;
array[37099] <= 16'b0000_0000_0000_0000;
array[37100] <= 16'b0000_0000_0000_0000;
array[37101] <= 16'b0000_0000_0000_0000;
array[37102] <= 16'b0000_0000_0000_0000;
array[37103] <= 16'b0000_0000_0000_0000;
array[37104] <= 16'b0000_0000_0000_0000;
array[37105] <= 16'b0000_0000_0000_0000;
array[37106] <= 16'b0000_0000_0000_0000;
array[37107] <= 16'b0000_0000_0000_0000;
array[37108] <= 16'b0000_0000_0000_0000;
array[37109] <= 16'b0000_0000_0000_0000;
array[37110] <= 16'b0000_0000_0000_0000;
array[37111] <= 16'b0000_0000_0000_0000;
array[37112] <= 16'b0000_0000_0000_0000;
array[37113] <= 16'b0000_0000_0000_0000;
array[37114] <= 16'b0000_0000_0000_0000;
array[37115] <= 16'b0000_0000_0000_0000;
array[37116] <= 16'b0000_0000_0000_0000;
array[37117] <= 16'b0000_0000_0000_0000;
array[37118] <= 16'b0000_0000_0000_0000;
array[37119] <= 16'b0000_0000_0000_0000;
array[37120] <= 16'b0000_0000_0000_0000;
array[37121] <= 16'b0000_0000_0000_0000;
array[37122] <= 16'b0000_0000_0000_0000;
array[37123] <= 16'b0000_0000_0000_0000;
array[37124] <= 16'b0000_0000_0000_0000;
array[37125] <= 16'b0000_0000_0000_0000;
array[37126] <= 16'b0000_0000_0000_0000;
array[37127] <= 16'b0000_0000_0000_0000;
array[37128] <= 16'b0000_0000_0000_0000;
array[37129] <= 16'b0000_0000_0000_0000;
array[37130] <= 16'b0000_0000_0000_0000;
array[37131] <= 16'b0000_0000_0000_0000;
array[37132] <= 16'b0000_0000_0000_0000;
array[37133] <= 16'b0000_0000_0000_0000;
array[37134] <= 16'b0000_0000_0000_0000;
array[37135] <= 16'b0000_0000_0000_0000;
array[37136] <= 16'b0000_0000_0000_0000;
array[37137] <= 16'b0000_0000_0000_0000;
array[37138] <= 16'b0000_0000_0000_0000;
array[37139] <= 16'b0000_0000_0000_0000;
array[37140] <= 16'b0000_0000_0000_0000;
array[37141] <= 16'b0000_0000_0000_0000;
array[37142] <= 16'b0000_0000_0000_0000;
array[37143] <= 16'b0000_0000_0000_0000;
array[37144] <= 16'b0000_0000_0000_0000;
array[37145] <= 16'b0000_0000_0000_0000;
array[37146] <= 16'b0000_0000_0000_0000;
array[37147] <= 16'b0000_0000_0000_0000;
array[37148] <= 16'b0000_0000_0000_0000;
array[37149] <= 16'b0000_0000_0000_0000;
array[37150] <= 16'b0000_0000_0000_0000;
array[37151] <= 16'b0000_0000_0000_0000;
array[37152] <= 16'b0000_0000_0000_0000;
array[37153] <= 16'b0000_0000_0000_0000;
array[37154] <= 16'b0000_0000_0000_0000;
array[37155] <= 16'b0000_0000_0000_0000;
array[37156] <= 16'b0000_0000_0000_0000;
array[37157] <= 16'b0000_0000_0000_0000;
array[37158] <= 16'b0000_0000_0000_0000;
array[37159] <= 16'b0000_0000_0000_0000;
array[37160] <= 16'b0000_0000_0000_0000;
array[37161] <= 16'b0000_0000_0000_0000;
array[37162] <= 16'b0000_0000_0000_0000;
array[37163] <= 16'b0000_0000_0000_0000;
array[37164] <= 16'b0000_0000_0000_0000;
array[37165] <= 16'b0000_0000_0000_0000;
array[37166] <= 16'b0000_0000_0000_0000;
array[37167] <= 16'b0000_0000_0000_0000;
array[37168] <= 16'b0000_0000_0000_0000;
array[37169] <= 16'b0000_0000_0000_0000;
array[37170] <= 16'b0000_0000_0000_0000;
array[37171] <= 16'b0000_0000_0000_0000;
array[37172] <= 16'b0000_0000_0000_0000;
array[37173] <= 16'b0000_0000_0000_0000;
array[37174] <= 16'b0000_0000_0000_0000;
array[37175] <= 16'b0000_0000_0000_0000;
array[37176] <= 16'b0000_0000_0000_0000;
array[37177] <= 16'b0000_0000_0000_0000;
array[37178] <= 16'b0000_0000_0000_0000;
array[37179] <= 16'b0000_0000_0000_0000;
array[37180] <= 16'b0000_0000_0000_0000;
array[37181] <= 16'b0000_0000_0000_0000;
array[37182] <= 16'b0000_0000_0000_0000;
array[37183] <= 16'b0000_0000_0000_0000;
array[37184] <= 16'b0000_0000_0000_0000;
array[37185] <= 16'b0000_0000_0000_0000;
array[37186] <= 16'b0000_0000_0000_0000;
array[37187] <= 16'b0000_0000_0000_0000;
array[37188] <= 16'b0000_0000_0000_0000;
array[37189] <= 16'b0000_0000_0000_0000;
array[37190] <= 16'b0000_0000_0000_0000;
array[37191] <= 16'b0000_0000_0000_0000;
array[37192] <= 16'b0000_0000_0000_0000;
array[37193] <= 16'b0000_0000_0000_0000;
array[37194] <= 16'b0000_0000_0000_0000;
array[37195] <= 16'b0000_0000_0000_0000;
array[37196] <= 16'b0000_0000_0000_0000;
array[37197] <= 16'b0000_0000_0000_0000;
array[37198] <= 16'b0000_0000_0000_0000;
array[37199] <= 16'b0000_0000_0000_0000;
array[37200] <= 16'b0000_0000_0000_0000;
array[37201] <= 16'b0000_0000_0000_0000;
array[37202] <= 16'b0000_0000_0000_0000;
array[37203] <= 16'b0000_0000_0000_0000;
array[37204] <= 16'b0000_0000_0000_0000;
array[37205] <= 16'b0000_0000_0000_0000;
array[37206] <= 16'b0000_0000_0000_0000;
array[37207] <= 16'b0000_0000_0000_0000;
array[37208] <= 16'b0000_0000_0000_0000;
array[37209] <= 16'b0000_0000_0000_0000;
array[37210] <= 16'b0000_0000_0000_0000;
array[37211] <= 16'b0000_0000_0000_0000;
array[37212] <= 16'b0000_0000_0000_0000;
array[37213] <= 16'b0000_0000_0000_0000;
array[37214] <= 16'b0000_0000_0000_0000;
array[37215] <= 16'b0000_0000_0000_0000;
array[37216] <= 16'b0000_0000_0000_0000;
array[37217] <= 16'b0000_0000_0000_0000;
array[37218] <= 16'b0000_0000_0000_0000;
array[37219] <= 16'b0000_0000_0000_0000;
array[37220] <= 16'b0000_0000_0000_0000;
array[37221] <= 16'b0000_0000_0000_0000;
array[37222] <= 16'b0000_0000_0000_0000;
array[37223] <= 16'b0000_0000_0000_0000;
array[37224] <= 16'b0000_0000_0000_0000;
array[37225] <= 16'b0000_0000_0000_0000;
array[37226] <= 16'b0000_0000_0000_0000;
array[37227] <= 16'b0000_0000_0000_0000;
array[37228] <= 16'b0000_0000_0000_0000;
array[37229] <= 16'b0000_0000_0000_0000;
array[37230] <= 16'b0000_0000_0000_0000;
array[37231] <= 16'b0000_0000_0000_0000;
array[37232] <= 16'b0000_0000_0000_0000;
array[37233] <= 16'b0000_0000_0000_0000;
array[37234] <= 16'b0000_0000_0000_0000;
array[37235] <= 16'b0000_0000_0000_0000;
array[37236] <= 16'b0000_0000_0000_0000;
array[37237] <= 16'b0000_0000_0000_0000;
array[37238] <= 16'b0000_0000_0000_0000;
array[37239] <= 16'b0000_0000_0000_0000;
array[37240] <= 16'b0000_0000_0000_0000;
array[37241] <= 16'b0000_0000_0000_0000;
array[37242] <= 16'b0000_0000_0000_0000;
array[37243] <= 16'b0000_0000_0000_0000;
array[37244] <= 16'b0000_0000_0000_0000;
array[37245] <= 16'b0000_0000_0000_0000;
array[37246] <= 16'b0000_0000_0000_0000;
array[37247] <= 16'b0000_0000_0000_0000;
array[37248] <= 16'b0000_0000_0000_0000;
array[37249] <= 16'b0000_0000_0000_0000;
array[37250] <= 16'b0000_0000_0000_0000;
array[37251] <= 16'b0000_0000_0000_0000;
array[37252] <= 16'b0000_0000_0000_0000;
array[37253] <= 16'b0000_0000_0000_0000;
array[37254] <= 16'b0000_0000_0000_0000;
array[37255] <= 16'b0000_0000_0000_0000;
array[37256] <= 16'b0000_0000_0000_0000;
array[37257] <= 16'b0000_0000_0000_0000;
array[37258] <= 16'b0000_0000_0000_0000;
array[37259] <= 16'b0000_0000_0000_0000;
array[37260] <= 16'b0000_0000_0000_0000;
array[37261] <= 16'b0000_0000_0000_0000;
array[37262] <= 16'b0000_0000_0000_0000;
array[37263] <= 16'b0000_0000_0000_0000;
array[37264] <= 16'b0000_0000_0000_0000;
array[37265] <= 16'b0000_0000_0000_0000;
array[37266] <= 16'b0000_0000_0000_0000;
array[37267] <= 16'b0000_0000_0000_0000;
array[37268] <= 16'b0000_0000_0000_0000;
array[37269] <= 16'b0000_0000_0000_0000;
array[37270] <= 16'b0000_0000_0000_0000;
array[37271] <= 16'b0000_0000_0000_0000;
array[37272] <= 16'b0000_0000_0000_0000;
array[37273] <= 16'b0000_0000_0000_0000;
array[37274] <= 16'b0000_0000_0000_0000;
array[37275] <= 16'b0000_0000_0000_0000;
array[37276] <= 16'b0000_0000_0000_0000;
array[37277] <= 16'b0000_0000_0000_0000;
array[37278] <= 16'b0000_0000_0000_0000;
array[37279] <= 16'b0000_0000_0000_0000;
array[37280] <= 16'b0000_0000_0000_0000;
array[37281] <= 16'b0000_0000_0000_0000;
array[37282] <= 16'b0000_0000_0000_0000;
array[37283] <= 16'b0000_0000_0000_0000;
array[37284] <= 16'b0000_0000_0000_0000;
array[37285] <= 16'b0000_0000_0000_0000;
array[37286] <= 16'b0000_0000_0000_0000;
array[37287] <= 16'b0000_0000_0000_0000;
array[37288] <= 16'b0000_0000_0000_0000;
array[37289] <= 16'b0000_0000_0000_0000;
array[37290] <= 16'b0000_0000_0000_0000;
array[37291] <= 16'b0000_0000_0000_0000;
array[37292] <= 16'b0000_0000_0000_0000;
array[37293] <= 16'b0000_0000_0000_0000;
array[37294] <= 16'b0000_0000_0000_0000;
array[37295] <= 16'b0000_0000_0000_0000;
array[37296] <= 16'b0000_0000_0000_0000;
array[37297] <= 16'b0000_0000_0000_0000;
array[37298] <= 16'b0000_0000_0000_0000;
array[37299] <= 16'b0000_0000_0000_0000;
array[37300] <= 16'b0000_0000_0000_0000;
array[37301] <= 16'b0000_0000_0000_0000;
array[37302] <= 16'b0000_0000_0000_0000;
array[37303] <= 16'b0000_0000_0000_0000;
array[37304] <= 16'b0000_0000_0000_0000;
array[37305] <= 16'b0000_0000_0000_0000;
array[37306] <= 16'b0000_0000_0000_0000;
array[37307] <= 16'b0000_0000_0000_0000;
array[37308] <= 16'b0000_0000_0000_0000;
array[37309] <= 16'b0000_0000_0000_0000;
array[37310] <= 16'b0000_0000_0000_0000;
array[37311] <= 16'b0000_0000_0000_0000;
array[37312] <= 16'b0000_0000_0000_0000;
array[37313] <= 16'b0000_0000_0000_0000;
array[37314] <= 16'b0000_0000_0000_0000;
array[37315] <= 16'b0000_0000_0000_0000;
array[37316] <= 16'b0000_0000_0000_0000;
array[37317] <= 16'b0000_0000_0000_0000;
array[37318] <= 16'b0000_0000_0000_0000;
array[37319] <= 16'b0000_0000_0000_0000;
array[37320] <= 16'b0000_0000_0000_0000;
array[37321] <= 16'b0000_0000_0000_0000;
array[37322] <= 16'b0000_0000_0000_0000;
array[37323] <= 16'b0000_0000_0000_0000;
array[37324] <= 16'b0000_0000_0000_0000;
array[37325] <= 16'b0000_0000_0000_0000;
array[37326] <= 16'b0000_0000_0000_0000;
array[37327] <= 16'b0000_0000_0000_0000;
array[37328] <= 16'b0000_0000_0000_0000;
array[37329] <= 16'b0000_0000_0000_0000;
array[37330] <= 16'b0000_0000_0000_0000;
array[37331] <= 16'b0000_0000_0000_0000;
array[37332] <= 16'b0000_0000_0000_0000;
array[37333] <= 16'b0000_0000_0000_0000;
array[37334] <= 16'b0000_0000_0000_0000;
array[37335] <= 16'b0000_0000_0000_0000;
array[37336] <= 16'b0000_0000_0000_0000;
array[37337] <= 16'b0000_0000_0000_0000;
array[37338] <= 16'b0000_0000_0000_0000;
array[37339] <= 16'b0000_0000_0000_0000;
array[37340] <= 16'b0000_0000_0000_0000;
array[37341] <= 16'b0000_0000_0000_0000;
array[37342] <= 16'b0000_0000_0000_0000;
array[37343] <= 16'b0000_0000_0000_0000;
array[37344] <= 16'b0000_0000_0000_0000;
array[37345] <= 16'b0000_0000_0000_0000;
array[37346] <= 16'b0000_0000_0000_0000;
array[37347] <= 16'b0000_0000_0000_0000;
array[37348] <= 16'b0000_0000_0000_0000;
array[37349] <= 16'b0000_0000_0000_0000;
array[37350] <= 16'b0000_0000_0000_0000;
array[37351] <= 16'b0000_0000_0000_0000;
array[37352] <= 16'b0000_0000_0000_0000;
array[37353] <= 16'b0000_0000_0000_0000;
array[37354] <= 16'b0000_0000_0000_0000;
array[37355] <= 16'b0000_0000_0000_0000;
array[37356] <= 16'b0000_0000_0000_0000;
array[37357] <= 16'b0000_0000_0000_0000;
array[37358] <= 16'b0000_0000_0000_0000;
array[37359] <= 16'b0000_0000_0000_0000;
array[37360] <= 16'b0000_0000_0000_0000;
array[37361] <= 16'b0000_0000_0000_0000;
array[37362] <= 16'b0000_0000_0000_0000;
array[37363] <= 16'b0000_0000_0000_0000;
array[37364] <= 16'b0000_0000_0000_0000;
array[37365] <= 16'b0000_0000_0000_0000;
array[37366] <= 16'b0000_0000_0000_0000;
array[37367] <= 16'b0000_0000_0000_0000;
array[37368] <= 16'b0000_0000_0000_0000;
array[37369] <= 16'b0000_0000_0000_0000;
array[37370] <= 16'b0000_0000_0000_0000;
array[37371] <= 16'b0000_0000_0000_0000;
array[37372] <= 16'b0000_0000_0000_0000;
array[37373] <= 16'b0000_0000_0000_0000;
array[37374] <= 16'b0000_0000_0000_0000;
array[37375] <= 16'b0000_0000_0000_0000;
array[37376] <= 16'b0000_0000_0000_0000;
array[37377] <= 16'b0000_0000_0000_0000;
array[37378] <= 16'b0000_0000_0000_0000;
array[37379] <= 16'b0000_0000_0000_0000;
array[37380] <= 16'b0000_0000_0000_0000;
array[37381] <= 16'b0000_0000_0000_0000;
array[37382] <= 16'b0000_0000_0000_0000;
array[37383] <= 16'b0000_0000_0000_0000;
array[37384] <= 16'b0000_0000_0000_0000;
array[37385] <= 16'b0000_0000_0000_0000;
array[37386] <= 16'b0000_0000_0000_0000;
array[37387] <= 16'b0000_0000_0000_0000;
array[37388] <= 16'b0000_0000_0000_0000;
array[37389] <= 16'b0000_0000_0000_0000;
array[37390] <= 16'b0000_0000_0000_0000;
array[37391] <= 16'b0000_0000_0000_0000;
array[37392] <= 16'b0000_0000_0000_0000;
array[37393] <= 16'b0000_0000_0000_0000;
array[37394] <= 16'b0000_0000_0000_0000;
array[37395] <= 16'b0000_0000_0000_0000;
array[37396] <= 16'b0000_0000_0000_0000;
array[37397] <= 16'b0000_0000_0000_0000;
array[37398] <= 16'b0000_0000_0000_0000;
array[37399] <= 16'b0000_0000_0000_0000;
array[37400] <= 16'b0000_0000_0000_0000;
array[37401] <= 16'b0000_0000_0000_0000;
array[37402] <= 16'b0000_0000_0000_0000;
array[37403] <= 16'b0000_0000_0000_0000;
array[37404] <= 16'b0000_0000_0000_0000;
array[37405] <= 16'b0000_0000_0000_0000;
array[37406] <= 16'b0000_0000_0000_0000;
array[37407] <= 16'b0000_0000_0000_0000;
array[37408] <= 16'b0000_0000_0000_0000;
array[37409] <= 16'b0000_0000_0000_0000;
array[37410] <= 16'b0000_0000_0000_0000;
array[37411] <= 16'b0000_0000_0000_0000;
array[37412] <= 16'b0000_0000_0000_0000;
array[37413] <= 16'b0000_0000_0000_0000;
array[37414] <= 16'b0000_0000_0000_0000;
array[37415] <= 16'b0000_0000_0000_0000;
array[37416] <= 16'b0000_0000_0000_0000;
array[37417] <= 16'b0000_0000_0000_0000;
array[37418] <= 16'b0000_0000_0000_0000;
array[37419] <= 16'b0000_0000_0000_0000;
array[37420] <= 16'b0000_0000_0000_0000;
array[37421] <= 16'b0000_0000_0000_0000;
array[37422] <= 16'b0000_0000_0000_0000;
array[37423] <= 16'b0000_0000_0000_0000;
array[37424] <= 16'b0000_0000_0000_0000;
array[37425] <= 16'b0000_0000_0000_0000;
array[37426] <= 16'b0000_0000_0000_0000;
array[37427] <= 16'b0000_0000_0000_0000;
array[37428] <= 16'b0000_0000_0000_0000;
array[37429] <= 16'b0000_0000_0000_0000;
array[37430] <= 16'b0000_0000_0000_0000;
array[37431] <= 16'b0000_0000_0000_0000;
array[37432] <= 16'b0000_0000_0000_0000;
array[37433] <= 16'b0000_0000_0000_0000;
array[37434] <= 16'b0000_0000_0000_0000;
array[37435] <= 16'b0000_0000_0000_0000;
array[37436] <= 16'b0000_0000_0000_0000;
array[37437] <= 16'b0000_0000_0000_0000;
array[37438] <= 16'b0000_0000_0000_0000;
array[37439] <= 16'b0000_0000_0000_0000;
array[37440] <= 16'b0000_0000_0000_0000;
array[37441] <= 16'b0000_0000_0000_0000;
array[37442] <= 16'b0000_0000_0000_0000;
array[37443] <= 16'b0000_0000_0000_0000;
array[37444] <= 16'b0000_0000_0000_0000;
array[37445] <= 16'b0000_0000_0000_0000;
array[37446] <= 16'b0000_0000_0000_0000;
array[37447] <= 16'b0000_0000_0000_0000;
array[37448] <= 16'b0000_0000_0000_0000;
array[37449] <= 16'b0000_0000_0000_0000;
array[37450] <= 16'b0000_0000_0000_0000;
array[37451] <= 16'b0000_0000_0000_0000;
array[37452] <= 16'b0000_0000_0000_0000;
array[37453] <= 16'b0000_0000_0000_0000;
array[37454] <= 16'b0000_0000_0000_0000;
array[37455] <= 16'b0000_0000_0000_0000;
array[37456] <= 16'b0000_0000_0000_0000;
array[37457] <= 16'b0000_0000_0000_0000;
array[37458] <= 16'b0000_0000_0000_0000;
array[37459] <= 16'b0000_0000_0000_0000;
array[37460] <= 16'b0000_0000_0000_0000;
array[37461] <= 16'b0000_0000_0000_0000;
array[37462] <= 16'b0000_0000_0000_0000;
array[37463] <= 16'b0000_0000_0000_0000;
array[37464] <= 16'b0000_0000_0000_0000;
array[37465] <= 16'b0000_0000_0000_0000;
array[37466] <= 16'b0000_0000_0000_0000;
array[37467] <= 16'b0000_0000_0000_0000;
array[37468] <= 16'b0000_0000_0000_0000;
array[37469] <= 16'b0000_0000_0000_0000;
array[37470] <= 16'b0000_0000_0000_0000;
array[37471] <= 16'b0000_0000_0000_0000;
array[37472] <= 16'b0000_0000_0000_0000;
array[37473] <= 16'b0000_0000_0000_0000;
array[37474] <= 16'b0000_0000_0000_0000;
array[37475] <= 16'b0000_0000_0000_0000;
array[37476] <= 16'b0000_0000_0000_0000;
array[37477] <= 16'b0000_0000_0000_0000;
array[37478] <= 16'b0000_0000_0000_0000;
array[37479] <= 16'b0000_0000_0000_0000;
array[37480] <= 16'b0000_0000_0000_0000;
array[37481] <= 16'b0000_0000_0000_0000;
array[37482] <= 16'b0000_0000_0000_0000;
array[37483] <= 16'b0000_0000_0000_0000;
array[37484] <= 16'b0000_0000_0000_0000;
array[37485] <= 16'b0000_0000_0000_0000;
array[37486] <= 16'b0000_0000_0000_0000;
array[37487] <= 16'b0000_0000_0000_0000;
array[37488] <= 16'b0000_0000_0000_0000;
array[37489] <= 16'b0000_0000_0000_0000;
array[37490] <= 16'b0000_0000_0000_0000;
array[37491] <= 16'b0000_0000_0000_0000;
array[37492] <= 16'b0000_0000_0000_0000;
array[37493] <= 16'b0000_0000_0000_0000;
array[37494] <= 16'b0000_0000_0000_0000;
array[37495] <= 16'b0000_0000_0000_0000;
array[37496] <= 16'b0000_0000_0000_0000;
array[37497] <= 16'b0000_0000_0000_0000;
array[37498] <= 16'b0000_0000_0000_0000;
array[37499] <= 16'b0000_0000_0000_0000;
array[37500] <= 16'b0000_0000_0000_0000;
array[37501] <= 16'b0000_0000_0000_0000;
array[37502] <= 16'b0000_0000_0000_0000;
array[37503] <= 16'b0000_0000_0000_0000;
array[37504] <= 16'b0000_0000_0000_0000;
array[37505] <= 16'b0000_0000_0000_0000;
array[37506] <= 16'b0000_0000_0000_0000;
array[37507] <= 16'b0000_0000_0000_0000;
array[37508] <= 16'b0000_0000_0000_0000;
array[37509] <= 16'b0000_0000_0000_0000;
array[37510] <= 16'b0000_0000_0000_0000;
array[37511] <= 16'b0000_0000_0000_0000;
array[37512] <= 16'b0000_0000_0000_0000;
array[37513] <= 16'b0000_0000_0000_0000;
array[37514] <= 16'b0000_0000_0000_0000;
array[37515] <= 16'b0000_0000_0000_0000;
array[37516] <= 16'b0000_0000_0000_0000;
array[37517] <= 16'b0000_0000_0000_0000;
array[37518] <= 16'b0000_0000_0000_0000;
array[37519] <= 16'b0000_0000_0000_0000;
array[37520] <= 16'b0000_0000_0000_0000;
array[37521] <= 16'b0000_0000_0000_0000;
array[37522] <= 16'b0000_0000_0000_0000;
array[37523] <= 16'b0000_0000_0000_0000;
array[37524] <= 16'b0000_0000_0000_0000;
array[37525] <= 16'b0000_0000_0000_0000;
array[37526] <= 16'b0000_0000_0000_0000;
array[37527] <= 16'b0000_0000_0000_0000;
array[37528] <= 16'b0000_0000_0000_0000;
array[37529] <= 16'b0000_0000_0000_0000;
array[37530] <= 16'b0000_0000_0000_0000;
array[37531] <= 16'b0000_0000_0000_0000;
array[37532] <= 16'b0000_0000_0000_0000;
array[37533] <= 16'b0000_0000_0000_0000;
array[37534] <= 16'b0000_0000_0000_0000;
array[37535] <= 16'b0000_0000_0000_0000;
array[37536] <= 16'b0000_0000_0000_0000;
array[37537] <= 16'b0000_0000_0000_0000;
array[37538] <= 16'b0000_0000_0000_0000;
array[37539] <= 16'b0000_0000_0000_0000;
array[37540] <= 16'b0000_0000_0000_0000;
array[37541] <= 16'b0000_0000_0000_0000;
array[37542] <= 16'b0000_0000_0000_0000;
array[37543] <= 16'b0000_0000_0000_0000;
array[37544] <= 16'b0000_0000_0000_0000;
array[37545] <= 16'b0000_0000_0000_0000;
array[37546] <= 16'b0000_0000_0000_0000;
array[37547] <= 16'b0000_0000_0000_0000;
array[37548] <= 16'b0000_0000_0000_0000;
array[37549] <= 16'b0000_0000_0000_0000;
array[37550] <= 16'b0000_0000_0000_0000;
array[37551] <= 16'b0000_0000_0000_0000;
array[37552] <= 16'b0000_0000_0000_0000;
array[37553] <= 16'b0000_0000_0000_0000;
array[37554] <= 16'b0000_0000_0000_0000;
array[37555] <= 16'b0000_0000_0000_0000;
array[37556] <= 16'b0000_0000_0000_0000;
array[37557] <= 16'b0000_0000_0000_0000;
array[37558] <= 16'b0000_0000_0000_0000;
array[37559] <= 16'b0000_0000_0000_0000;
array[37560] <= 16'b0000_0000_0000_0000;
array[37561] <= 16'b0000_0000_0000_0000;
array[37562] <= 16'b0000_0000_0000_0000;
array[37563] <= 16'b0000_0000_0000_0000;
array[37564] <= 16'b0000_0000_0000_0000;
array[37565] <= 16'b0000_0000_0000_0000;
array[37566] <= 16'b0000_0000_0000_0000;
array[37567] <= 16'b0000_0000_0000_0000;
array[37568] <= 16'b0000_0000_0000_0000;
array[37569] <= 16'b0000_0000_0000_0000;
array[37570] <= 16'b0000_0000_0000_0000;
array[37571] <= 16'b0000_0000_0000_0000;
array[37572] <= 16'b0000_0000_0000_0000;
array[37573] <= 16'b0000_0000_0000_0000;
array[37574] <= 16'b0000_0000_0000_0000;
array[37575] <= 16'b0000_0000_0000_0000;
array[37576] <= 16'b0000_0000_0000_0000;
array[37577] <= 16'b0000_0000_0000_0000;
array[37578] <= 16'b0000_0000_0000_0000;
array[37579] <= 16'b0000_0000_0000_0000;
array[37580] <= 16'b0000_0000_0000_0000;
array[37581] <= 16'b0000_0000_0000_0000;
array[37582] <= 16'b0000_0000_0000_0000;
array[37583] <= 16'b0000_0000_0000_0000;
array[37584] <= 16'b0000_0000_0000_0000;
array[37585] <= 16'b0000_0000_0000_0000;
array[37586] <= 16'b0000_0000_0000_0000;
array[37587] <= 16'b0000_0000_0000_0000;
array[37588] <= 16'b0000_0000_0000_0000;
array[37589] <= 16'b0000_0000_0000_0000;
array[37590] <= 16'b0000_0000_0000_0000;
array[37591] <= 16'b0000_0000_0000_0000;
array[37592] <= 16'b0000_0000_0000_0000;
array[37593] <= 16'b0000_0000_0000_0000;
array[37594] <= 16'b0000_0000_0000_0000;
array[37595] <= 16'b0000_0000_0000_0000;
array[37596] <= 16'b0000_0000_0000_0000;
array[37597] <= 16'b0000_0000_0000_0000;
array[37598] <= 16'b0000_0000_0000_0000;
array[37599] <= 16'b0000_0000_0000_0000;
array[37600] <= 16'b0000_0000_0000_0000;
array[37601] <= 16'b0000_0000_0000_0000;
array[37602] <= 16'b0000_0000_0000_0000;
array[37603] <= 16'b0000_0000_0000_0000;
array[37604] <= 16'b0000_0000_0000_0000;
array[37605] <= 16'b0000_0000_0000_0000;
array[37606] <= 16'b0000_0000_0000_0000;
array[37607] <= 16'b0000_0000_0000_0000;
array[37608] <= 16'b0000_0000_0000_0000;
array[37609] <= 16'b0000_0000_0000_0000;
array[37610] <= 16'b0000_0000_0000_0000;
array[37611] <= 16'b0000_0000_0000_0000;
array[37612] <= 16'b0000_0000_0000_0000;
array[37613] <= 16'b0000_0000_0000_0000;
array[37614] <= 16'b0000_0000_0000_0000;
array[37615] <= 16'b0000_0000_0000_0000;
array[37616] <= 16'b0000_0000_0000_0000;
array[37617] <= 16'b0000_0000_0000_0000;
array[37618] <= 16'b0000_0000_0000_0000;
array[37619] <= 16'b0000_0000_0000_0000;
array[37620] <= 16'b0000_0000_0000_0000;
array[37621] <= 16'b0000_0000_0000_0000;
array[37622] <= 16'b0000_0000_0000_0000;
array[37623] <= 16'b0000_0000_0000_0000;
array[37624] <= 16'b0000_0000_0000_0000;
array[37625] <= 16'b0000_0000_0000_0000;
array[37626] <= 16'b0000_0000_0000_0000;
array[37627] <= 16'b0000_0000_0000_0000;
array[37628] <= 16'b0000_0000_0000_0000;
array[37629] <= 16'b0000_0000_0000_0000;
array[37630] <= 16'b0000_0000_0000_0000;
array[37631] <= 16'b0000_0000_0000_0000;
array[37632] <= 16'b0000_0000_0000_0000;
array[37633] <= 16'b0000_0000_0000_0000;
array[37634] <= 16'b0000_0000_0000_0000;
array[37635] <= 16'b0000_0000_0000_0000;
array[37636] <= 16'b0000_0000_0000_0000;
array[37637] <= 16'b0000_0000_0000_0000;
array[37638] <= 16'b0000_0000_0000_0000;
array[37639] <= 16'b0000_0000_0000_0000;
array[37640] <= 16'b0000_0000_0000_0000;
array[37641] <= 16'b0000_0000_0000_0000;
array[37642] <= 16'b0000_0000_0000_0000;
array[37643] <= 16'b0000_0000_0000_0000;
array[37644] <= 16'b0000_0000_0000_0000;
array[37645] <= 16'b0000_0000_0000_0000;
array[37646] <= 16'b0000_0000_0000_0000;
array[37647] <= 16'b0000_0000_0000_0000;
array[37648] <= 16'b0000_0000_0000_0000;
array[37649] <= 16'b0000_0000_0000_0000;
array[37650] <= 16'b0000_0000_0000_0000;
array[37651] <= 16'b0000_0000_0000_0000;
array[37652] <= 16'b0000_0000_0000_0000;
array[37653] <= 16'b0000_0000_0000_0000;
array[37654] <= 16'b0000_0000_0000_0000;
array[37655] <= 16'b0000_0000_0000_0000;
array[37656] <= 16'b0000_0000_0000_0000;
array[37657] <= 16'b0000_0000_0000_0000;
array[37658] <= 16'b0000_0000_0000_0000;
array[37659] <= 16'b0000_0000_0000_0000;
array[37660] <= 16'b0000_0000_0000_0000;
array[37661] <= 16'b0000_0000_0000_0000;
array[37662] <= 16'b0000_0000_0000_0000;
array[37663] <= 16'b0000_0000_0000_0000;
array[37664] <= 16'b0000_0000_0000_0000;
array[37665] <= 16'b0000_0000_0000_0000;
array[37666] <= 16'b0000_0000_0000_0000;
array[37667] <= 16'b0000_0000_0000_0000;
array[37668] <= 16'b0000_0000_0000_0000;
array[37669] <= 16'b0000_0000_0000_0000;
array[37670] <= 16'b0000_0000_0000_0000;
array[37671] <= 16'b0000_0000_0000_0000;
array[37672] <= 16'b0000_0000_0000_0000;
array[37673] <= 16'b0000_0000_0000_0000;
array[37674] <= 16'b0000_0000_0000_0000;
array[37675] <= 16'b0000_0000_0000_0000;
array[37676] <= 16'b0000_0000_0000_0000;
array[37677] <= 16'b0000_0000_0000_0000;
array[37678] <= 16'b0000_0000_0000_0000;
array[37679] <= 16'b0000_0000_0000_0000;
array[37680] <= 16'b0000_0000_0000_0000;
array[37681] <= 16'b0000_0000_0000_0000;
array[37682] <= 16'b0000_0000_0000_0000;
array[37683] <= 16'b0000_0000_0000_0000;
array[37684] <= 16'b0000_0000_0000_0000;
array[37685] <= 16'b0000_0000_0000_0000;
array[37686] <= 16'b0000_0000_0000_0000;
array[37687] <= 16'b0000_0000_0000_0000;
array[37688] <= 16'b0000_0000_0000_0000;
array[37689] <= 16'b0000_0000_0000_0000;
array[37690] <= 16'b0000_0000_0000_0000;
array[37691] <= 16'b0000_0000_0000_0000;
array[37692] <= 16'b0000_0000_0000_0000;
array[37693] <= 16'b0000_0000_0000_0000;
array[37694] <= 16'b0000_0000_0000_0000;
array[37695] <= 16'b0000_0000_0000_0000;
array[37696] <= 16'b0000_0000_0000_0000;
array[37697] <= 16'b0000_0000_0000_0000;
array[37698] <= 16'b0000_0000_0000_0000;
array[37699] <= 16'b0000_0000_0000_0000;
array[37700] <= 16'b0000_0000_0000_0000;
array[37701] <= 16'b0000_0000_0000_0000;
array[37702] <= 16'b0000_0000_0000_0000;
array[37703] <= 16'b0000_0000_0000_0000;
array[37704] <= 16'b0000_0000_0000_0000;
array[37705] <= 16'b0000_0000_0000_0000;
array[37706] <= 16'b0000_0000_0000_0000;
array[37707] <= 16'b0000_0000_0000_0000;
array[37708] <= 16'b0000_0000_0000_0000;
array[37709] <= 16'b0000_0000_0000_0000;
array[37710] <= 16'b0000_0000_0000_0000;
array[37711] <= 16'b0000_0000_0000_0000;
array[37712] <= 16'b0000_0000_0000_0000;
array[37713] <= 16'b0000_0000_0000_0000;
array[37714] <= 16'b0000_0000_0000_0000;
array[37715] <= 16'b0000_0000_0000_0000;
array[37716] <= 16'b0000_0000_0000_0000;
array[37717] <= 16'b0000_0000_0000_0000;
array[37718] <= 16'b0000_0000_0000_0000;
array[37719] <= 16'b0000_0000_0000_0000;
array[37720] <= 16'b0000_0000_0000_0000;
array[37721] <= 16'b0000_0000_0000_0000;
array[37722] <= 16'b0000_0000_0000_0000;
array[37723] <= 16'b0000_0000_0000_0000;
array[37724] <= 16'b0000_0000_0000_0000;
array[37725] <= 16'b0000_0000_0000_0000;
array[37726] <= 16'b0000_0000_0000_0000;
array[37727] <= 16'b0000_0000_0000_0000;
array[37728] <= 16'b0000_0000_0000_0000;
array[37729] <= 16'b0000_0000_0000_0000;
array[37730] <= 16'b0000_0000_0000_0000;
array[37731] <= 16'b0000_0000_0000_0000;
array[37732] <= 16'b0000_0000_0000_0000;
array[37733] <= 16'b0000_0000_0000_0000;
array[37734] <= 16'b0000_0000_0000_0000;
array[37735] <= 16'b0000_0000_0000_0000;
array[37736] <= 16'b0000_0000_0000_0000;
array[37737] <= 16'b0000_0000_0000_0000;
array[37738] <= 16'b0000_0000_0000_0000;
array[37739] <= 16'b0000_0000_0000_0000;
array[37740] <= 16'b0000_0000_0000_0000;
array[37741] <= 16'b0000_0000_0000_0000;
array[37742] <= 16'b0000_0000_0000_0000;
array[37743] <= 16'b0000_0000_0000_0000;
array[37744] <= 16'b0000_0000_0000_0000;
array[37745] <= 16'b0000_0000_0000_0000;
array[37746] <= 16'b0000_0000_0000_0000;
array[37747] <= 16'b0000_0000_0000_0000;
array[37748] <= 16'b0000_0000_0000_0000;
array[37749] <= 16'b0000_0000_0000_0000;
array[37750] <= 16'b0000_0000_0000_0000;
array[37751] <= 16'b0000_0000_0000_0000;
array[37752] <= 16'b0000_0000_0000_0000;
array[37753] <= 16'b0000_0000_0000_0000;
array[37754] <= 16'b0000_0000_0000_0000;
array[37755] <= 16'b0000_0000_0000_0000;
array[37756] <= 16'b0000_0000_0000_0000;
array[37757] <= 16'b0000_0000_0000_0000;
array[37758] <= 16'b0000_0000_0000_0000;
array[37759] <= 16'b0000_0000_0000_0000;
array[37760] <= 16'b0000_0000_0000_0000;
array[37761] <= 16'b0000_0000_0000_0000;
array[37762] <= 16'b0000_0000_0000_0000;
array[37763] <= 16'b0000_0000_0000_0000;
array[37764] <= 16'b0000_0000_0000_0000;
array[37765] <= 16'b0000_0000_0000_0000;
array[37766] <= 16'b0000_0000_0000_0000;
array[37767] <= 16'b0000_0000_0000_0000;
array[37768] <= 16'b0000_0000_0000_0000;
array[37769] <= 16'b0000_0000_0000_0000;
array[37770] <= 16'b0000_0000_0000_0000;
array[37771] <= 16'b0000_0000_0000_0000;
array[37772] <= 16'b0000_0000_0000_0000;
array[37773] <= 16'b0000_0000_0000_0000;
array[37774] <= 16'b0000_0000_0000_0000;
array[37775] <= 16'b0000_0000_0000_0000;
array[37776] <= 16'b0000_0000_0000_0000;
array[37777] <= 16'b0000_0000_0000_0000;
array[37778] <= 16'b0000_0000_0000_0000;
array[37779] <= 16'b0000_0000_0000_0000;
array[37780] <= 16'b0000_0000_0000_0000;
array[37781] <= 16'b0000_0000_0000_0000;
array[37782] <= 16'b0000_0000_0000_0000;
array[37783] <= 16'b0000_0000_0000_0000;
array[37784] <= 16'b0000_0000_0000_0000;
array[37785] <= 16'b0000_0000_0000_0000;
array[37786] <= 16'b0000_0000_0000_0000;
array[37787] <= 16'b0000_0000_0000_0000;
array[37788] <= 16'b0000_0000_0000_0000;
array[37789] <= 16'b0000_0000_0000_0000;
array[37790] <= 16'b0000_0000_0000_0000;
array[37791] <= 16'b0000_0000_0000_0000;
array[37792] <= 16'b0000_0000_0000_0000;
array[37793] <= 16'b0000_0000_0000_0000;
array[37794] <= 16'b0000_0000_0000_0000;
array[37795] <= 16'b0000_0000_0000_0000;
array[37796] <= 16'b0000_0000_0000_0000;
array[37797] <= 16'b0000_0000_0000_0000;
array[37798] <= 16'b0000_0000_0000_0000;
array[37799] <= 16'b0000_0000_0000_0000;
array[37800] <= 16'b0000_0000_0000_0000;
array[37801] <= 16'b0000_0000_0000_0000;
array[37802] <= 16'b0000_0000_0000_0000;
array[37803] <= 16'b0000_0000_0000_0000;
array[37804] <= 16'b0000_0000_0000_0000;
array[37805] <= 16'b0000_0000_0000_0000;
array[37806] <= 16'b0000_0000_0000_0000;
array[37807] <= 16'b0000_0000_0000_0000;
array[37808] <= 16'b0000_0000_0000_0000;
array[37809] <= 16'b0000_0000_0000_0000;
array[37810] <= 16'b0000_0000_0000_0000;
array[37811] <= 16'b0000_0000_0000_0000;
array[37812] <= 16'b0000_0000_0000_0000;
array[37813] <= 16'b0000_0000_0000_0000;
array[37814] <= 16'b0000_0000_0000_0000;
array[37815] <= 16'b0000_0000_0000_0000;
array[37816] <= 16'b0000_0000_0000_0000;
array[37817] <= 16'b0000_0000_0000_0000;
array[37818] <= 16'b0000_0000_0000_0000;
array[37819] <= 16'b0000_0000_0000_0000;
array[37820] <= 16'b0000_0000_0000_0000;
array[37821] <= 16'b0000_0000_0000_0000;
array[37822] <= 16'b0000_0000_0000_0000;
array[37823] <= 16'b0000_0000_0000_0000;
array[37824] <= 16'b0000_0000_0000_0000;
array[37825] <= 16'b0000_0000_0000_0000;
array[37826] <= 16'b0000_0000_0000_0000;
array[37827] <= 16'b0000_0000_0000_0000;
array[37828] <= 16'b0000_0000_0000_0000;
array[37829] <= 16'b0000_0000_0000_0000;
array[37830] <= 16'b0000_0000_0000_0000;
array[37831] <= 16'b0000_0000_0000_0000;
array[37832] <= 16'b0000_0000_0000_0000;
array[37833] <= 16'b0000_0000_0000_0000;
array[37834] <= 16'b0000_0000_0000_0000;
array[37835] <= 16'b0000_0000_0000_0000;
array[37836] <= 16'b0000_0000_0000_0000;
array[37837] <= 16'b0000_0000_0000_0000;
array[37838] <= 16'b0000_0000_0000_0000;
array[37839] <= 16'b0000_0000_0000_0000;
array[37840] <= 16'b0000_0000_0000_0000;
array[37841] <= 16'b0000_0000_0000_0000;
array[37842] <= 16'b0000_0000_0000_0000;
array[37843] <= 16'b0000_0000_0000_0000;
array[37844] <= 16'b0000_0000_0000_0000;
array[37845] <= 16'b0000_0000_0000_0000;
array[37846] <= 16'b0000_0000_0000_0000;
array[37847] <= 16'b0000_0000_0000_0000;
array[37848] <= 16'b0000_0000_0000_0000;
array[37849] <= 16'b0000_0000_0000_0000;
array[37850] <= 16'b0000_0000_0000_0000;
array[37851] <= 16'b0000_0000_0000_0000;
array[37852] <= 16'b0000_0000_0000_0000;
array[37853] <= 16'b0000_0000_0000_0000;
array[37854] <= 16'b0000_0000_0000_0000;
array[37855] <= 16'b0000_0000_0000_0000;
array[37856] <= 16'b0000_0000_0000_0000;
array[37857] <= 16'b0000_0000_0000_0000;
array[37858] <= 16'b0000_0000_0000_0000;
array[37859] <= 16'b0000_0000_0000_0000;
array[37860] <= 16'b0000_0000_0000_0000;
array[37861] <= 16'b0000_0000_0000_0000;
array[37862] <= 16'b0000_0000_0000_0000;
array[37863] <= 16'b0000_0000_0000_0000;
array[37864] <= 16'b0000_0000_0000_0000;
array[37865] <= 16'b0000_0000_0000_0000;
array[37866] <= 16'b0000_0000_0000_0000;
array[37867] <= 16'b0000_0000_0000_0000;
array[37868] <= 16'b0000_0000_0000_0000;
array[37869] <= 16'b0000_0000_0000_0000;
array[37870] <= 16'b0000_0000_0000_0000;
array[37871] <= 16'b0000_0000_0000_0000;
array[37872] <= 16'b0000_0000_0000_0000;
array[37873] <= 16'b0000_0000_0000_0000;
array[37874] <= 16'b0000_0000_0000_0000;
array[37875] <= 16'b0000_0000_0000_0000;
array[37876] <= 16'b0000_0000_0000_0000;
array[37877] <= 16'b0000_0000_0000_0000;
array[37878] <= 16'b0000_0000_0000_0000;
array[37879] <= 16'b0000_0000_0000_0000;
array[37880] <= 16'b0000_0000_0000_0000;
array[37881] <= 16'b0000_0000_0000_0000;
array[37882] <= 16'b0000_0000_0000_0000;
array[37883] <= 16'b0000_0000_0000_0000;
array[37884] <= 16'b0000_0000_0000_0000;
array[37885] <= 16'b0000_0000_0000_0000;
array[37886] <= 16'b0000_0000_0000_0000;
array[37887] <= 16'b0000_0000_0000_0000;
array[37888] <= 16'b0000_0000_0000_0000;
array[37889] <= 16'b0000_0000_0000_0000;
array[37890] <= 16'b0000_0000_0000_0000;
array[37891] <= 16'b0000_0000_0000_0000;
array[37892] <= 16'b0000_0000_0000_0000;
array[37893] <= 16'b0000_0000_0000_0000;
array[37894] <= 16'b0000_0000_0000_0000;
array[37895] <= 16'b0000_0000_0000_0000;
array[37896] <= 16'b0000_0000_0000_0000;
array[37897] <= 16'b0000_0000_0000_0000;
array[37898] <= 16'b0000_0000_0000_0000;
array[37899] <= 16'b0000_0000_0000_0000;
array[37900] <= 16'b0000_0000_0000_0000;
array[37901] <= 16'b0000_0000_0000_0000;
array[37902] <= 16'b0000_0000_0000_0000;
array[37903] <= 16'b0000_0000_0000_0000;
array[37904] <= 16'b0000_0000_0000_0000;
array[37905] <= 16'b0000_0000_0000_0000;
array[37906] <= 16'b0000_0000_0000_0000;
array[37907] <= 16'b0000_0000_0000_0000;
array[37908] <= 16'b0000_0000_0000_0000;
array[37909] <= 16'b0000_0000_0000_0000;
array[37910] <= 16'b0000_0000_0000_0000;
array[37911] <= 16'b0000_0000_0000_0000;
array[37912] <= 16'b0000_0000_0000_0000;
array[37913] <= 16'b0000_0000_0000_0000;
array[37914] <= 16'b0000_0000_0000_0000;
array[37915] <= 16'b0000_0000_0000_0000;
array[37916] <= 16'b0000_0000_0000_0000;
array[37917] <= 16'b0000_0000_0000_0000;
array[37918] <= 16'b0000_0000_0000_0000;
array[37919] <= 16'b0000_0000_0000_0000;
array[37920] <= 16'b0000_0000_0000_0000;
array[37921] <= 16'b0000_0000_0000_0000;
array[37922] <= 16'b0000_0000_0000_0000;
array[37923] <= 16'b0000_0000_0000_0000;
array[37924] <= 16'b0000_0000_0000_0000;
array[37925] <= 16'b0000_0000_0000_0000;
array[37926] <= 16'b0000_0000_0000_0000;
array[37927] <= 16'b0000_0000_0000_0000;
array[37928] <= 16'b0000_0000_0000_0000;
array[37929] <= 16'b0000_0000_0000_0000;
array[37930] <= 16'b0000_0000_0000_0000;
array[37931] <= 16'b0000_0000_0000_0000;
array[37932] <= 16'b0000_0000_0000_0000;
array[37933] <= 16'b0000_0000_0000_0000;
array[37934] <= 16'b0000_0000_0000_0000;
array[37935] <= 16'b0000_0000_0000_0000;
array[37936] <= 16'b0000_0000_0000_0000;
array[37937] <= 16'b0000_0000_0000_0000;
array[37938] <= 16'b0000_0000_0000_0000;
array[37939] <= 16'b0000_0000_0000_0000;
array[37940] <= 16'b0000_0000_0000_0000;
array[37941] <= 16'b0000_0000_0000_0000;
array[37942] <= 16'b0000_0000_0000_0000;
array[37943] <= 16'b0000_0000_0000_0000;
array[37944] <= 16'b0000_0000_0000_0000;
array[37945] <= 16'b0000_0000_0000_0000;
array[37946] <= 16'b0000_0000_0000_0000;
array[37947] <= 16'b0000_0000_0000_0000;
array[37948] <= 16'b0000_0000_0000_0000;
array[37949] <= 16'b0000_0000_0000_0000;
array[37950] <= 16'b0000_0000_0000_0000;
array[37951] <= 16'b0000_0000_0000_0000;
array[37952] <= 16'b0000_0000_0000_0000;
array[37953] <= 16'b0000_0000_0000_0000;
array[37954] <= 16'b0000_0000_0000_0000;
array[37955] <= 16'b0000_0000_0000_0000;
array[37956] <= 16'b0000_0000_0000_0000;
array[37957] <= 16'b0000_0000_0000_0000;
array[37958] <= 16'b0000_0000_0000_0000;
array[37959] <= 16'b0000_0000_0000_0000;
array[37960] <= 16'b0000_0000_0000_0000;
array[37961] <= 16'b0000_0000_0000_0000;
array[37962] <= 16'b0000_0000_0000_0000;
array[37963] <= 16'b0000_0000_0000_0000;
array[37964] <= 16'b0000_0000_0000_0000;
array[37965] <= 16'b0000_0000_0000_0000;
array[37966] <= 16'b0000_0000_0000_0000;
array[37967] <= 16'b0000_0000_0000_0000;
array[37968] <= 16'b0000_0000_0000_0000;
array[37969] <= 16'b0000_0000_0000_0000;
array[37970] <= 16'b0000_0000_0000_0000;
array[37971] <= 16'b0000_0000_0000_0000;
array[37972] <= 16'b0000_0000_0000_0000;
array[37973] <= 16'b0000_0000_0000_0000;
array[37974] <= 16'b0000_0000_0000_0000;
array[37975] <= 16'b0000_0000_0000_0000;
array[37976] <= 16'b0000_0000_0000_0000;
array[37977] <= 16'b0000_0000_0000_0000;
array[37978] <= 16'b0000_0000_0000_0000;
array[37979] <= 16'b0000_0000_0000_0000;
array[37980] <= 16'b0000_0000_0000_0000;
array[37981] <= 16'b0000_0000_0000_0000;
array[37982] <= 16'b0000_0000_0000_0000;
array[37983] <= 16'b0000_0000_0000_0000;
array[37984] <= 16'b0000_0000_0000_0000;
array[37985] <= 16'b0000_0000_0000_0000;
array[37986] <= 16'b0000_0000_0000_0000;
array[37987] <= 16'b0000_0000_0000_0000;
array[37988] <= 16'b0000_0000_0000_0000;
array[37989] <= 16'b0000_0000_0000_0000;
array[37990] <= 16'b0000_0000_0000_0000;
array[37991] <= 16'b0000_0000_0000_0000;
array[37992] <= 16'b0000_0000_0000_0000;
array[37993] <= 16'b0000_0000_0000_0000;
array[37994] <= 16'b0000_0000_0000_0000;
array[37995] <= 16'b0000_0000_0000_0000;
array[37996] <= 16'b0000_0000_0000_0000;
array[37997] <= 16'b0000_0000_0000_0000;
array[37998] <= 16'b0000_0000_0000_0000;
array[37999] <= 16'b0000_0000_0000_0000;
array[38000] <= 16'b0000_0000_0000_0000;
array[38001] <= 16'b0000_0000_0000_0000;
array[38002] <= 16'b0000_0000_0000_0000;
array[38003] <= 16'b0000_0000_0000_0000;
array[38004] <= 16'b0000_0000_0000_0000;
array[38005] <= 16'b0000_0000_0000_0000;
array[38006] <= 16'b0000_0000_0000_0000;
array[38007] <= 16'b0000_0000_0000_0000;
array[38008] <= 16'b0000_0000_0000_0000;
array[38009] <= 16'b0000_0000_0000_0000;
array[38010] <= 16'b0000_0000_0000_0000;
array[38011] <= 16'b0000_0000_0000_0000;
array[38012] <= 16'b0000_0000_0000_0000;
array[38013] <= 16'b0000_0000_0000_0000;
array[38014] <= 16'b0000_0000_0000_0000;
array[38015] <= 16'b0000_0000_0000_0000;
array[38016] <= 16'b0000_0000_0000_0000;
array[38017] <= 16'b0000_0000_0000_0000;
array[38018] <= 16'b0000_0000_0000_0000;
array[38019] <= 16'b0000_0000_0000_0000;
array[38020] <= 16'b0000_0000_0000_0000;
array[38021] <= 16'b0000_0000_0000_0000;
array[38022] <= 16'b0000_0000_0000_0000;
array[38023] <= 16'b0000_0000_0000_0000;
array[38024] <= 16'b0000_0000_0000_0000;
array[38025] <= 16'b0000_0000_0000_0000;
array[38026] <= 16'b0000_0000_0000_0000;
array[38027] <= 16'b0000_0000_0000_0000;
array[38028] <= 16'b0000_0000_0000_0000;
array[38029] <= 16'b0000_0000_0000_0000;
array[38030] <= 16'b0000_0000_0000_0000;
array[38031] <= 16'b0000_0000_0000_0000;
array[38032] <= 16'b0000_0000_0000_0000;
array[38033] <= 16'b0000_0000_0000_0000;
array[38034] <= 16'b0000_0000_0000_0000;
array[38035] <= 16'b0000_0000_0000_0000;
array[38036] <= 16'b0000_0000_0000_0000;
array[38037] <= 16'b0000_0000_0000_0000;
array[38038] <= 16'b0000_0000_0000_0000;
array[38039] <= 16'b0000_0000_0000_0000;
array[38040] <= 16'b0000_0000_0000_0000;
array[38041] <= 16'b0000_0000_0000_0000;
array[38042] <= 16'b0000_0000_0000_0000;
array[38043] <= 16'b0000_0000_0000_0000;
array[38044] <= 16'b0000_0000_0000_0000;
array[38045] <= 16'b0000_0000_0000_0000;
array[38046] <= 16'b0000_0000_0000_0000;
array[38047] <= 16'b0000_0000_0000_0000;
array[38048] <= 16'b0000_0000_0000_0000;
array[38049] <= 16'b0000_0000_0000_0000;
array[38050] <= 16'b0000_0000_0000_0000;
array[38051] <= 16'b0000_0000_0000_0000;
array[38052] <= 16'b0000_0000_0000_0000;
array[38053] <= 16'b0000_0000_0000_0000;
array[38054] <= 16'b0000_0000_0000_0000;
array[38055] <= 16'b0000_0000_0000_0000;
array[38056] <= 16'b0000_0000_0000_0000;
array[38057] <= 16'b0000_0000_0000_0000;
array[38058] <= 16'b0000_0000_0000_0000;
array[38059] <= 16'b0000_0000_0000_0000;
array[38060] <= 16'b0000_0000_0000_0000;
array[38061] <= 16'b0000_0000_0000_0000;
array[38062] <= 16'b0000_0000_0000_0000;
array[38063] <= 16'b0000_0000_0000_0000;
array[38064] <= 16'b0000_0000_0000_0000;
array[38065] <= 16'b0000_0000_0000_0000;
array[38066] <= 16'b0000_0000_0000_0000;
array[38067] <= 16'b0000_0000_0000_0000;
array[38068] <= 16'b0000_0000_0000_0000;
array[38069] <= 16'b0000_0000_0000_0000;
array[38070] <= 16'b0000_0000_0000_0000;
array[38071] <= 16'b0000_0000_0000_0000;
array[38072] <= 16'b0000_0000_0000_0000;
array[38073] <= 16'b0000_0000_0000_0000;
array[38074] <= 16'b0000_0000_0000_0000;
array[38075] <= 16'b0000_0000_0000_0000;
array[38076] <= 16'b0000_0000_0000_0000;
array[38077] <= 16'b0000_0000_0000_0000;
array[38078] <= 16'b0000_0000_0000_0000;
array[38079] <= 16'b0000_0000_0000_0000;
array[38080] <= 16'b0000_0000_0000_0000;
array[38081] <= 16'b0000_0000_0000_0000;
array[38082] <= 16'b0000_0000_0000_0000;
array[38083] <= 16'b0000_0000_0000_0000;
array[38084] <= 16'b0000_0000_0000_0000;
array[38085] <= 16'b0000_0000_0000_0000;
array[38086] <= 16'b0000_0000_0000_0000;
array[38087] <= 16'b0000_0000_0000_0000;
array[38088] <= 16'b0000_0000_0000_0000;
array[38089] <= 16'b0000_0000_0000_0000;
array[38090] <= 16'b0000_0000_0000_0000;
array[38091] <= 16'b0000_0000_0000_0000;
array[38092] <= 16'b0000_0000_0000_0000;
array[38093] <= 16'b0000_0000_0000_0000;
array[38094] <= 16'b0000_0000_0000_0000;
array[38095] <= 16'b0000_0000_0000_0000;
array[38096] <= 16'b0000_0000_0000_0000;
array[38097] <= 16'b0000_0000_0000_0000;
array[38098] <= 16'b0000_0000_0000_0000;
array[38099] <= 16'b0000_0000_0000_0000;
array[38100] <= 16'b0000_0000_0000_0000;
array[38101] <= 16'b0000_0000_0000_0000;
array[38102] <= 16'b0000_0000_0000_0000;
array[38103] <= 16'b0000_0000_0000_0000;
array[38104] <= 16'b0000_0000_0000_0000;
array[38105] <= 16'b0000_0000_0000_0000;
array[38106] <= 16'b0000_0000_0000_0000;
array[38107] <= 16'b0000_0000_0000_0000;
array[38108] <= 16'b0000_0000_0000_0000;
array[38109] <= 16'b0000_0000_0000_0000;
array[38110] <= 16'b0000_0000_0000_0000;
array[38111] <= 16'b0000_0000_0000_0000;
array[38112] <= 16'b0000_0000_0000_0000;
array[38113] <= 16'b0000_0000_0000_0000;
array[38114] <= 16'b0000_0000_0000_0000;
array[38115] <= 16'b0000_0000_0000_0000;
array[38116] <= 16'b0000_0000_0000_0000;
array[38117] <= 16'b0000_0000_0000_0000;
array[38118] <= 16'b0000_0000_0000_0000;
array[38119] <= 16'b0000_0000_0000_0000;
array[38120] <= 16'b0000_0000_0000_0000;
array[38121] <= 16'b0000_0000_0000_0000;
array[38122] <= 16'b0000_0000_0000_0000;
array[38123] <= 16'b0000_0000_0000_0000;
array[38124] <= 16'b0000_0000_0000_0000;
array[38125] <= 16'b0000_0000_0000_0000;
array[38126] <= 16'b0000_0000_0000_0000;
array[38127] <= 16'b0000_0000_0000_0000;
array[38128] <= 16'b0000_0000_0000_0000;
array[38129] <= 16'b0000_0000_0000_0000;
array[38130] <= 16'b0000_0000_0000_0000;
array[38131] <= 16'b0000_0000_0000_0000;
array[38132] <= 16'b0000_0000_0000_0000;
array[38133] <= 16'b0000_0000_0000_0000;
array[38134] <= 16'b0000_0000_0000_0000;
array[38135] <= 16'b0000_0000_0000_0000;
array[38136] <= 16'b0000_0000_0000_0000;
array[38137] <= 16'b0000_0000_0000_0000;
array[38138] <= 16'b0000_0000_0000_0000;
array[38139] <= 16'b0000_0000_0000_0000;
array[38140] <= 16'b0000_0000_0000_0000;
array[38141] <= 16'b0000_0000_0000_0000;
array[38142] <= 16'b0000_0000_0000_0000;
array[38143] <= 16'b0000_0000_0000_0000;
array[38144] <= 16'b0000_0000_0000_0000;
array[38145] <= 16'b0000_0000_0000_0000;
array[38146] <= 16'b0000_0000_0000_0000;
array[38147] <= 16'b0000_0000_0000_0000;
array[38148] <= 16'b0000_0000_0000_0000;
array[38149] <= 16'b0000_0000_0000_0000;
array[38150] <= 16'b0000_0000_0000_0000;
array[38151] <= 16'b0000_0000_0000_0000;
array[38152] <= 16'b0000_0000_0000_0000;
array[38153] <= 16'b0000_0000_0000_0000;
array[38154] <= 16'b0000_0000_0000_0000;
array[38155] <= 16'b0000_0000_0000_0000;
array[38156] <= 16'b0000_0000_0000_0000;
array[38157] <= 16'b0000_0000_0000_0000;
array[38158] <= 16'b0000_0000_0000_0000;
array[38159] <= 16'b0000_0000_0000_0000;
array[38160] <= 16'b0000_0000_0000_0000;
array[38161] <= 16'b0000_0000_0000_0000;
array[38162] <= 16'b0000_0000_0000_0000;
array[38163] <= 16'b0000_0000_0000_0000;
array[38164] <= 16'b0000_0000_0000_0000;
array[38165] <= 16'b0000_0000_0000_0000;
array[38166] <= 16'b0000_0000_0000_0000;
array[38167] <= 16'b0000_0000_0000_0000;
array[38168] <= 16'b0000_0000_0000_0000;
array[38169] <= 16'b0000_0000_0000_0000;
array[38170] <= 16'b0000_0000_0000_0000;
array[38171] <= 16'b0000_0000_0000_0000;
array[38172] <= 16'b0000_0000_0000_0000;
array[38173] <= 16'b0000_0000_0000_0000;
array[38174] <= 16'b0000_0000_0000_0000;
array[38175] <= 16'b0000_0000_0000_0000;
array[38176] <= 16'b0000_0000_0000_0000;
array[38177] <= 16'b0000_0000_0000_0000;
array[38178] <= 16'b0000_0000_0000_0000;
array[38179] <= 16'b0000_0000_0000_0000;
array[38180] <= 16'b0000_0000_0000_0000;
array[38181] <= 16'b0000_0000_0000_0000;
array[38182] <= 16'b0000_0000_0000_0000;
array[38183] <= 16'b0000_0000_0000_0000;
array[38184] <= 16'b0000_0000_0000_0000;
array[38185] <= 16'b0000_0000_0000_0000;
array[38186] <= 16'b0000_0000_0000_0000;
array[38187] <= 16'b0000_0000_0000_0000;
array[38188] <= 16'b0000_0000_0000_0000;
array[38189] <= 16'b0000_0000_0000_0000;
array[38190] <= 16'b0000_0000_0000_0000;
array[38191] <= 16'b0000_0000_0000_0000;
array[38192] <= 16'b0000_0000_0000_0000;
array[38193] <= 16'b0000_0000_0000_0000;
array[38194] <= 16'b0000_0000_0000_0000;
array[38195] <= 16'b0000_0000_0000_0000;
array[38196] <= 16'b0000_0000_0000_0000;
array[38197] <= 16'b0000_0000_0000_0000;
array[38198] <= 16'b0000_0000_0000_0000;
array[38199] <= 16'b0000_0000_0000_0000;
array[38200] <= 16'b0000_0000_0000_0000;
array[38201] <= 16'b0000_0000_0000_0000;
array[38202] <= 16'b0000_0000_0000_0000;
array[38203] <= 16'b0000_0000_0000_0000;
array[38204] <= 16'b0000_0000_0000_0000;
array[38205] <= 16'b0000_0000_0000_0000;
array[38206] <= 16'b0000_0000_0000_0000;
array[38207] <= 16'b0000_0000_0000_0000;
array[38208] <= 16'b0000_0000_0000_0000;
array[38209] <= 16'b0000_0000_0000_0000;
array[38210] <= 16'b0000_0000_0000_0000;
array[38211] <= 16'b0000_0000_0000_0000;
array[38212] <= 16'b0000_0000_0000_0000;
array[38213] <= 16'b0000_0000_0000_0000;
array[38214] <= 16'b0000_0000_0000_0000;
array[38215] <= 16'b0000_0000_0000_0000;
array[38216] <= 16'b0000_0000_0000_0000;
array[38217] <= 16'b0000_0000_0000_0000;
array[38218] <= 16'b0000_0000_0000_0000;
array[38219] <= 16'b0000_0000_0000_0000;
array[38220] <= 16'b0000_0000_0000_0000;
array[38221] <= 16'b0000_0000_0000_0000;
array[38222] <= 16'b0000_0000_0000_0000;
array[38223] <= 16'b0000_0000_0000_0000;
array[38224] <= 16'b0000_0000_0000_0000;
array[38225] <= 16'b0000_0000_0000_0000;
array[38226] <= 16'b0000_0000_0000_0000;
array[38227] <= 16'b0000_0000_0000_0000;
array[38228] <= 16'b0000_0000_0000_0000;
array[38229] <= 16'b0000_0000_0000_0000;
array[38230] <= 16'b0000_0000_0000_0000;
array[38231] <= 16'b0000_0000_0000_0000;
array[38232] <= 16'b0000_0000_0000_0000;
array[38233] <= 16'b0000_0000_0000_0000;
array[38234] <= 16'b0000_0000_0000_0000;
array[38235] <= 16'b0000_0000_0000_0000;
array[38236] <= 16'b0000_0000_0000_0000;
array[38237] <= 16'b0000_0000_0000_0000;
array[38238] <= 16'b0000_0000_0000_0000;
array[38239] <= 16'b0000_0000_0000_0000;
array[38240] <= 16'b0000_0000_0000_0000;
array[38241] <= 16'b0000_0000_0000_0000;
array[38242] <= 16'b0000_0000_0000_0000;
array[38243] <= 16'b0000_0000_0000_0000;
array[38244] <= 16'b0000_0000_0000_0000;
array[38245] <= 16'b0000_0000_0000_0000;
array[38246] <= 16'b0000_0000_0000_0000;
array[38247] <= 16'b0000_0000_0000_0000;
array[38248] <= 16'b0000_0000_0000_0000;
array[38249] <= 16'b0000_0000_0000_0000;
array[38250] <= 16'b0000_0000_0000_0000;
array[38251] <= 16'b0000_0000_0000_0000;
array[38252] <= 16'b0000_0000_0000_0000;
array[38253] <= 16'b0000_0000_0000_0000;
array[38254] <= 16'b0000_0000_0000_0000;
array[38255] <= 16'b0000_0000_0000_0000;
array[38256] <= 16'b0000_0000_0000_0000;
array[38257] <= 16'b0000_0000_0000_0000;
array[38258] <= 16'b0000_0000_0000_0000;
array[38259] <= 16'b0000_0000_0000_0000;
array[38260] <= 16'b0000_0000_0000_0000;
array[38261] <= 16'b0000_0000_0000_0000;
array[38262] <= 16'b0000_0000_0000_0000;
array[38263] <= 16'b0000_0000_0000_0000;
array[38264] <= 16'b0000_0000_0000_0000;
array[38265] <= 16'b0000_0000_0000_0000;
array[38266] <= 16'b0000_0000_0000_0000;
array[38267] <= 16'b0000_0000_0000_0000;
array[38268] <= 16'b0000_0000_0000_0000;
array[38269] <= 16'b0000_0000_0000_0000;
array[38270] <= 16'b0000_0000_0000_0000;
array[38271] <= 16'b0000_0000_0000_0000;
array[38272] <= 16'b0000_0000_0000_0000;
array[38273] <= 16'b0000_0000_0000_0000;
array[38274] <= 16'b0000_0000_0000_0000;
array[38275] <= 16'b0000_0000_0000_0000;
array[38276] <= 16'b0000_0000_0000_0000;
array[38277] <= 16'b0000_0000_0000_0000;
array[38278] <= 16'b0000_0000_0000_0000;
array[38279] <= 16'b0000_0000_0000_0000;
array[38280] <= 16'b0000_0000_0000_0000;
array[38281] <= 16'b0000_0000_0000_0000;
array[38282] <= 16'b0000_0000_0000_0000;
array[38283] <= 16'b0000_0000_0000_0000;
array[38284] <= 16'b0000_0000_0000_0000;
array[38285] <= 16'b0000_0000_0000_0000;
array[38286] <= 16'b0000_0000_0000_0000;
array[38287] <= 16'b0000_0000_0000_0000;
array[38288] <= 16'b0000_0000_0000_0000;
array[38289] <= 16'b0000_0000_0000_0000;
array[38290] <= 16'b0000_0000_0000_0000;
array[38291] <= 16'b0000_0000_0000_0000;
array[38292] <= 16'b0000_0000_0000_0000;
array[38293] <= 16'b0000_0000_0000_0000;
array[38294] <= 16'b0000_0000_0000_0000;
array[38295] <= 16'b0000_0000_0000_0000;
array[38296] <= 16'b0000_0000_0000_0000;
array[38297] <= 16'b0000_0000_0000_0000;
array[38298] <= 16'b0000_0000_0000_0000;
array[38299] <= 16'b0000_0000_0000_0000;
array[38300] <= 16'b0000_0000_0000_0000;
array[38301] <= 16'b0000_0000_0000_0000;
array[38302] <= 16'b0000_0000_0000_0000;
array[38303] <= 16'b0000_0000_0000_0000;
array[38304] <= 16'b0000_0000_0000_0000;
array[38305] <= 16'b0000_0000_0000_0000;
array[38306] <= 16'b0000_0000_0000_0000;
array[38307] <= 16'b0000_0000_0000_0000;
array[38308] <= 16'b0000_0000_0000_0000;
array[38309] <= 16'b0000_0000_0000_0000;
array[38310] <= 16'b0000_0000_0000_0000;
array[38311] <= 16'b0000_0000_0000_0000;
array[38312] <= 16'b0000_0000_0000_0000;
array[38313] <= 16'b0000_0000_0000_0000;
array[38314] <= 16'b0000_0000_0000_0000;
array[38315] <= 16'b0000_0000_0000_0000;
array[38316] <= 16'b0000_0000_0000_0000;
array[38317] <= 16'b0000_0000_0000_0000;
array[38318] <= 16'b0000_0000_0000_0000;
array[38319] <= 16'b0000_0000_0000_0000;
array[38320] <= 16'b0000_0000_0000_0000;
array[38321] <= 16'b0000_0000_0000_0000;
array[38322] <= 16'b0000_0000_0000_0000;
array[38323] <= 16'b0000_0000_0000_0000;
array[38324] <= 16'b0000_0000_0000_0000;
array[38325] <= 16'b0000_0000_0000_0000;
array[38326] <= 16'b0000_0000_0000_0000;
array[38327] <= 16'b0000_0000_0000_0000;
array[38328] <= 16'b0000_0000_0000_0000;
array[38329] <= 16'b0000_0000_0000_0000;
array[38330] <= 16'b0000_0000_0000_0000;
array[38331] <= 16'b0000_0000_0000_0000;
array[38332] <= 16'b0000_0000_0000_0000;
array[38333] <= 16'b0000_0000_0000_0000;
array[38334] <= 16'b0000_0000_0000_0000;
array[38335] <= 16'b0000_0000_0000_0000;
array[38336] <= 16'b0000_0000_0000_0000;
array[38337] <= 16'b0000_0000_0000_0000;
array[38338] <= 16'b0000_0000_0000_0000;
array[38339] <= 16'b0000_0000_0000_0000;
array[38340] <= 16'b0000_0000_0000_0000;
array[38341] <= 16'b0000_0000_0000_0000;
array[38342] <= 16'b0000_0000_0000_0000;
array[38343] <= 16'b0000_0000_0000_0000;
array[38344] <= 16'b0000_0000_0000_0000;
array[38345] <= 16'b0000_0000_0000_0000;
array[38346] <= 16'b0000_0000_0000_0000;
array[38347] <= 16'b0000_0000_0000_0000;
array[38348] <= 16'b0000_0000_0000_0000;
array[38349] <= 16'b0000_0000_0000_0000;
array[38350] <= 16'b0000_0000_0000_0000;
array[38351] <= 16'b0000_0000_0000_0000;
array[38352] <= 16'b0000_0000_0000_0000;
array[38353] <= 16'b0000_0000_0000_0000;
array[38354] <= 16'b0000_0000_0000_0000;
array[38355] <= 16'b0000_0000_0000_0000;
array[38356] <= 16'b0000_0000_0000_0000;
array[38357] <= 16'b0000_0000_0000_0000;
array[38358] <= 16'b0000_0000_0000_0000;
array[38359] <= 16'b0000_0000_0000_0000;
array[38360] <= 16'b0000_0000_0000_0000;
array[38361] <= 16'b0000_0000_0000_0000;
array[38362] <= 16'b0000_0000_0000_0000;
array[38363] <= 16'b0000_0000_0000_0000;
array[38364] <= 16'b0000_0000_0000_0000;
array[38365] <= 16'b0000_0000_0000_0000;
array[38366] <= 16'b0000_0000_0000_0000;
array[38367] <= 16'b0000_0000_0000_0000;
array[38368] <= 16'b0000_0000_0000_0000;
array[38369] <= 16'b0000_0000_0000_0000;
array[38370] <= 16'b0000_0000_0000_0000;
array[38371] <= 16'b0000_0000_0000_0000;
array[38372] <= 16'b0000_0000_0000_0000;
array[38373] <= 16'b0000_0000_0000_0000;
array[38374] <= 16'b0000_0000_0000_0000;
array[38375] <= 16'b0000_0000_0000_0000;
array[38376] <= 16'b0000_0000_0000_0000;
array[38377] <= 16'b0000_0000_0000_0000;
array[38378] <= 16'b0000_0000_0000_0000;
array[38379] <= 16'b0000_0000_0000_0000;
array[38380] <= 16'b0000_0000_0000_0000;
array[38381] <= 16'b0000_0000_0000_0000;
array[38382] <= 16'b0000_0000_0000_0000;
array[38383] <= 16'b0000_0000_0000_0000;
array[38384] <= 16'b0000_0000_0000_0000;
array[38385] <= 16'b0000_0000_0000_0000;
array[38386] <= 16'b0000_0000_0000_0000;
array[38387] <= 16'b0000_0000_0000_0000;
array[38388] <= 16'b0000_0000_0000_0000;
array[38389] <= 16'b0000_0000_0000_0000;
array[38390] <= 16'b0000_0000_0000_0000;
array[38391] <= 16'b0000_0000_0000_0000;
array[38392] <= 16'b0000_0000_0000_0000;
array[38393] <= 16'b0000_0000_0000_0000;
array[38394] <= 16'b0000_0000_0000_0000;
array[38395] <= 16'b0000_0000_0000_0000;
array[38396] <= 16'b0000_0000_0000_0000;
array[38397] <= 16'b0000_0000_0000_0000;
array[38398] <= 16'b0000_0000_0000_0000;
array[38399] <= 16'b0000_0000_0000_0000;
array[38400] <= 16'b0000_0000_0000_0000;
array[38401] <= 16'b0000_0000_0000_0000;
array[38402] <= 16'b0000_0000_0000_0000;
array[38403] <= 16'b0000_0000_0000_0000;
array[38404] <= 16'b0000_0000_0000_0000;
array[38405] <= 16'b0000_0000_0000_0000;
array[38406] <= 16'b0000_0000_0000_0000;
array[38407] <= 16'b0000_0000_0000_0000;
array[38408] <= 16'b0000_0000_0000_0000;
array[38409] <= 16'b0000_0000_0000_0000;
array[38410] <= 16'b0000_0000_0000_0000;
array[38411] <= 16'b0000_0000_0000_0000;
array[38412] <= 16'b0000_0000_0000_0000;
array[38413] <= 16'b0000_0000_0000_0000;
array[38414] <= 16'b0000_0000_0000_0000;
array[38415] <= 16'b0000_0000_0000_0000;
array[38416] <= 16'b0000_0000_0000_0000;
array[38417] <= 16'b0000_0000_0000_0000;
array[38418] <= 16'b0000_0000_0000_0000;
array[38419] <= 16'b0000_0000_0000_0000;
array[38420] <= 16'b0000_0000_0000_0000;
array[38421] <= 16'b0000_0000_0000_0000;
array[38422] <= 16'b0000_0000_0000_0000;
array[38423] <= 16'b0000_0000_0000_0000;
array[38424] <= 16'b0000_0000_0000_0000;
array[38425] <= 16'b0000_0000_0000_0000;
array[38426] <= 16'b0000_0000_0000_0000;
array[38427] <= 16'b0000_0000_0000_0000;
array[38428] <= 16'b0000_0000_0000_0000;
array[38429] <= 16'b0000_0000_0000_0000;
array[38430] <= 16'b0000_0000_0000_0000;
array[38431] <= 16'b0000_0000_0000_0000;
array[38432] <= 16'b0000_0000_0000_0000;
array[38433] <= 16'b0000_0000_0000_0000;
array[38434] <= 16'b0000_0000_0000_0000;
array[38435] <= 16'b0000_0000_0000_0000;
array[38436] <= 16'b0000_0000_0000_0000;
array[38437] <= 16'b0000_0000_0000_0000;
array[38438] <= 16'b0000_0000_0000_0000;
array[38439] <= 16'b0000_0000_0000_0000;
array[38440] <= 16'b0000_0000_0000_0000;
array[38441] <= 16'b0000_0000_0000_0000;
array[38442] <= 16'b0000_0000_0000_0000;
array[38443] <= 16'b0000_0000_0000_0000;
array[38444] <= 16'b0000_0000_0000_0000;
array[38445] <= 16'b0000_0000_0000_0000;
array[38446] <= 16'b0000_0000_0000_0000;
array[38447] <= 16'b0000_0000_0000_0000;
array[38448] <= 16'b0000_0000_0000_0000;
array[38449] <= 16'b0000_0000_0000_0000;
array[38450] <= 16'b0000_0000_0000_0000;
array[38451] <= 16'b0000_0000_0000_0000;
array[38452] <= 16'b0000_0000_0000_0000;
array[38453] <= 16'b0000_0000_0000_0000;
array[38454] <= 16'b0000_0000_0000_0000;
array[38455] <= 16'b0000_0000_0000_0000;
array[38456] <= 16'b0000_0000_0000_0000;
array[38457] <= 16'b0000_0000_0000_0000;
array[38458] <= 16'b0000_0000_0000_0000;
array[38459] <= 16'b0000_0000_0000_0000;
array[38460] <= 16'b0000_0000_0000_0000;
array[38461] <= 16'b0000_0000_0000_0000;
array[38462] <= 16'b0000_0000_0000_0000;
array[38463] <= 16'b0000_0000_0000_0000;
array[38464] <= 16'b0000_0000_0000_0000;
array[38465] <= 16'b0000_0000_0000_0000;
array[38466] <= 16'b0000_0000_0000_0000;
array[38467] <= 16'b0000_0000_0000_0000;
array[38468] <= 16'b0000_0000_0000_0000;
array[38469] <= 16'b0000_0000_0000_0000;
array[38470] <= 16'b0000_0000_0000_0000;
array[38471] <= 16'b0000_0000_0000_0000;
array[38472] <= 16'b0000_0000_0000_0000;
array[38473] <= 16'b0000_0000_0000_0000;
array[38474] <= 16'b0000_0000_0000_0000;
array[38475] <= 16'b0000_0000_0000_0000;
array[38476] <= 16'b0000_0000_0000_0000;
array[38477] <= 16'b0000_0000_0000_0000;
array[38478] <= 16'b0000_0000_0000_0000;
array[38479] <= 16'b0000_0000_0000_0000;
array[38480] <= 16'b0000_0000_0000_0000;
array[38481] <= 16'b0000_0000_0000_0000;
array[38482] <= 16'b0000_0000_0000_0000;
array[38483] <= 16'b0000_0000_0000_0000;
array[38484] <= 16'b0000_0000_0000_0000;
array[38485] <= 16'b0000_0000_0000_0000;
array[38486] <= 16'b0000_0000_0000_0000;
array[38487] <= 16'b0000_0000_0000_0000;
array[38488] <= 16'b0000_0000_0000_0000;
array[38489] <= 16'b0000_0000_0000_0000;
array[38490] <= 16'b0000_0000_0000_0000;
array[38491] <= 16'b0000_0000_0000_0000;
array[38492] <= 16'b0000_0000_0000_0000;
array[38493] <= 16'b0000_0000_0000_0000;
array[38494] <= 16'b0000_0000_0000_0000;
array[38495] <= 16'b0000_0000_0000_0000;
array[38496] <= 16'b0000_0000_0000_0000;
array[38497] <= 16'b0000_0000_0000_0000;
array[38498] <= 16'b0000_0000_0000_0000;
array[38499] <= 16'b0000_0000_0000_0000;
array[38500] <= 16'b0000_0000_0000_0000;
array[38501] <= 16'b0000_0000_0000_0000;
array[38502] <= 16'b0000_0000_0000_0000;
array[38503] <= 16'b0000_0000_0000_0000;
array[38504] <= 16'b0000_0000_0000_0000;
array[38505] <= 16'b0000_0000_0000_0000;
array[38506] <= 16'b0000_0000_0000_0000;
array[38507] <= 16'b0000_0000_0000_0000;
array[38508] <= 16'b0000_0000_0000_0000;
array[38509] <= 16'b0000_0000_0000_0000;
array[38510] <= 16'b0000_0000_0000_0000;
array[38511] <= 16'b0000_0000_0000_0000;
array[38512] <= 16'b0000_0000_0000_0000;
array[38513] <= 16'b0000_0000_0000_0000;
array[38514] <= 16'b0000_0000_0000_0000;
array[38515] <= 16'b0000_0000_0000_0000;
array[38516] <= 16'b0000_0000_0000_0000;
array[38517] <= 16'b0000_0000_0000_0000;
array[38518] <= 16'b0000_0000_0000_0000;
array[38519] <= 16'b0000_0000_0000_0000;
array[38520] <= 16'b0000_0000_0000_0000;
array[38521] <= 16'b0000_0000_0000_0000;
array[38522] <= 16'b0000_0000_0000_0000;
array[38523] <= 16'b0000_0000_0000_0000;
array[38524] <= 16'b0000_0000_0000_0000;
array[38525] <= 16'b0000_0000_0000_0000;
array[38526] <= 16'b0000_0000_0000_0000;
array[38527] <= 16'b0000_0000_0000_0000;
array[38528] <= 16'b0000_0000_0000_0000;
array[38529] <= 16'b0000_0000_0000_0000;
array[38530] <= 16'b0000_0000_0000_0000;
array[38531] <= 16'b0000_0000_0000_0000;
array[38532] <= 16'b0000_0000_0000_0000;
array[38533] <= 16'b0000_0000_0000_0000;
array[38534] <= 16'b0000_0000_0000_0000;
array[38535] <= 16'b0000_0000_0000_0000;
array[38536] <= 16'b0000_0000_0000_0000;
array[38537] <= 16'b0000_0000_0000_0000;
array[38538] <= 16'b0000_0000_0000_0000;
array[38539] <= 16'b0000_0000_0000_0000;
array[38540] <= 16'b0000_0000_0000_0000;
array[38541] <= 16'b0000_0000_0000_0000;
array[38542] <= 16'b0000_0000_0000_0000;
array[38543] <= 16'b0000_0000_0000_0000;
array[38544] <= 16'b0000_0000_0000_0000;
array[38545] <= 16'b0000_0000_0000_0000;
array[38546] <= 16'b0000_0000_0000_0000;
array[38547] <= 16'b0000_0000_0000_0000;
array[38548] <= 16'b0000_0000_0000_0000;
array[38549] <= 16'b0000_0000_0000_0000;
array[38550] <= 16'b0000_0000_0000_0000;
array[38551] <= 16'b0000_0000_0000_0000;
array[38552] <= 16'b0000_0000_0000_0000;
array[38553] <= 16'b0000_0000_0000_0000;
array[38554] <= 16'b0000_0000_0000_0000;
array[38555] <= 16'b0000_0000_0000_0000;
array[38556] <= 16'b0000_0000_0000_0000;
array[38557] <= 16'b0000_0000_0000_0000;
array[38558] <= 16'b0000_0000_0000_0000;
array[38559] <= 16'b0000_0000_0000_0000;
array[38560] <= 16'b0000_0000_0000_0000;
array[38561] <= 16'b0000_0000_0000_0000;
array[38562] <= 16'b0000_0000_0000_0000;
array[38563] <= 16'b0000_0000_0000_0000;
array[38564] <= 16'b0000_0000_0000_0000;
array[38565] <= 16'b0000_0000_0000_0000;
array[38566] <= 16'b0000_0000_0000_0000;
array[38567] <= 16'b0000_0000_0000_0000;
array[38568] <= 16'b0000_0000_0000_0000;
array[38569] <= 16'b0000_0000_0000_0000;
array[38570] <= 16'b0000_0000_0000_0000;
array[38571] <= 16'b0000_0000_0000_0000;
array[38572] <= 16'b0000_0000_0000_0000;
array[38573] <= 16'b0000_0000_0000_0000;
array[38574] <= 16'b0000_0000_0000_0000;
array[38575] <= 16'b0000_0000_0000_0000;
array[38576] <= 16'b0000_0000_0000_0000;
array[38577] <= 16'b0000_0000_0000_0000;
array[38578] <= 16'b0000_0000_0000_0000;
array[38579] <= 16'b0000_0000_0000_0000;
array[38580] <= 16'b0000_0000_0000_0000;
array[38581] <= 16'b0000_0000_0000_0000;
array[38582] <= 16'b0000_0000_0000_0000;
array[38583] <= 16'b0000_0000_0000_0000;
array[38584] <= 16'b0000_0000_0000_0000;
array[38585] <= 16'b0000_0000_0000_0000;
array[38586] <= 16'b0000_0000_0000_0000;
array[38587] <= 16'b0000_0000_0000_0000;
array[38588] <= 16'b0000_0000_0000_0000;
array[38589] <= 16'b0000_0000_0000_0000;
array[38590] <= 16'b0000_0000_0000_0000;
array[38591] <= 16'b0000_0000_0000_0000;
array[38592] <= 16'b0000_0000_0000_0000;
array[38593] <= 16'b0000_0000_0000_0000;
array[38594] <= 16'b0000_0000_0000_0000;
array[38595] <= 16'b0000_0000_0000_0000;
array[38596] <= 16'b0000_0000_0000_0000;
array[38597] <= 16'b0000_0000_0000_0000;
array[38598] <= 16'b0000_0000_0000_0000;
array[38599] <= 16'b0000_0000_0000_0000;
array[38600] <= 16'b0000_0000_0000_0000;
array[38601] <= 16'b0000_0000_0000_0000;
array[38602] <= 16'b0000_0000_0000_0000;
array[38603] <= 16'b0000_0000_0000_0000;
array[38604] <= 16'b0000_0000_0000_0000;
array[38605] <= 16'b0000_0000_0000_0000;
array[38606] <= 16'b0000_0000_0000_0000;
array[38607] <= 16'b0000_0000_0000_0000;
array[38608] <= 16'b0000_0000_0000_0000;
array[38609] <= 16'b0000_0000_0000_0000;
array[38610] <= 16'b0000_0000_0000_0000;
array[38611] <= 16'b0000_0000_0000_0000;
array[38612] <= 16'b0000_0000_0000_0000;
array[38613] <= 16'b0000_0000_0000_0000;
array[38614] <= 16'b0000_0000_0000_0000;
array[38615] <= 16'b0000_0000_0000_0000;
array[38616] <= 16'b0000_0000_0000_0000;
array[38617] <= 16'b0000_0000_0000_0000;
array[38618] <= 16'b0000_0000_0000_0000;
array[38619] <= 16'b0000_0000_0000_0000;
array[38620] <= 16'b0000_0000_0000_0000;
array[38621] <= 16'b0000_0000_0000_0000;
array[38622] <= 16'b0000_0000_0000_0000;
array[38623] <= 16'b0000_0000_0000_0000;
array[38624] <= 16'b0000_0000_0000_0000;
array[38625] <= 16'b0000_0000_0000_0000;
array[38626] <= 16'b0000_0000_0000_0000;
array[38627] <= 16'b0000_0000_0000_0000;
array[38628] <= 16'b0000_0000_0000_0000;
array[38629] <= 16'b0000_0000_0000_0000;
array[38630] <= 16'b0000_0000_0000_0000;
array[38631] <= 16'b0000_0000_0000_0000;
array[38632] <= 16'b0000_0000_0000_0000;
array[38633] <= 16'b0000_0000_0000_0000;
array[38634] <= 16'b0000_0000_0000_0000;
array[38635] <= 16'b0000_0000_0000_0000;
array[38636] <= 16'b0000_0000_0000_0000;
array[38637] <= 16'b0000_0000_0000_0000;
array[38638] <= 16'b0000_0000_0000_0000;
array[38639] <= 16'b0000_0000_0000_0000;
array[38640] <= 16'b0000_0000_0000_0000;
array[38641] <= 16'b0000_0000_0000_0000;
array[38642] <= 16'b0000_0000_0000_0000;
array[38643] <= 16'b0000_0000_0000_0000;
array[38644] <= 16'b0000_0000_0000_0000;
array[38645] <= 16'b0000_0000_0000_0000;
array[38646] <= 16'b0000_0000_0000_0000;
array[38647] <= 16'b0000_0000_0000_0000;
array[38648] <= 16'b0000_0000_0000_0000;
array[38649] <= 16'b0000_0000_0000_0000;
array[38650] <= 16'b0000_0000_0000_0000;
array[38651] <= 16'b0000_0000_0000_0000;
array[38652] <= 16'b0000_0000_0000_0000;
array[38653] <= 16'b0000_0000_0000_0000;
array[38654] <= 16'b0000_0000_0000_0000;
array[38655] <= 16'b0000_0000_0000_0000;
array[38656] <= 16'b0000_0000_0000_0000;
array[38657] <= 16'b0000_0000_0000_0000;
array[38658] <= 16'b0000_0000_0000_0000;
array[38659] <= 16'b0000_0000_0000_0000;
array[38660] <= 16'b0000_0000_0000_0000;
array[38661] <= 16'b0000_0000_0000_0000;
array[38662] <= 16'b0000_0000_0000_0000;
array[38663] <= 16'b0000_0000_0000_0000;
array[38664] <= 16'b0000_0000_0000_0000;
array[38665] <= 16'b0000_0000_0000_0000;
array[38666] <= 16'b0000_0000_0000_0000;
array[38667] <= 16'b0000_0000_0000_0000;
array[38668] <= 16'b0000_0000_0000_0000;
array[38669] <= 16'b0000_0000_0000_0000;
array[38670] <= 16'b0000_0000_0000_0000;
array[38671] <= 16'b0000_0000_0000_0000;
array[38672] <= 16'b0000_0000_0000_0000;
array[38673] <= 16'b0000_0000_0000_0000;
array[38674] <= 16'b0000_0000_0000_0000;
array[38675] <= 16'b0000_0000_0000_0000;
array[38676] <= 16'b0000_0000_0000_0000;
array[38677] <= 16'b0000_0000_0000_0000;
array[38678] <= 16'b0000_0000_0000_0000;
array[38679] <= 16'b0000_0000_0000_0000;
array[38680] <= 16'b0000_0000_0000_0000;
array[38681] <= 16'b0000_0000_0000_0000;
array[38682] <= 16'b0000_0000_0000_0000;
array[38683] <= 16'b0000_0000_0000_0000;
array[38684] <= 16'b0000_0000_0000_0000;
array[38685] <= 16'b0000_0000_0000_0000;
array[38686] <= 16'b0000_0000_0000_0000;
array[38687] <= 16'b0000_0000_0000_0000;
array[38688] <= 16'b0000_0000_0000_0000;
array[38689] <= 16'b0000_0000_0000_0000;
array[38690] <= 16'b0000_0000_0000_0000;
array[38691] <= 16'b0000_0000_0000_0000;
array[38692] <= 16'b0000_0000_0000_0000;
array[38693] <= 16'b0000_0000_0000_0000;
array[38694] <= 16'b0000_0000_0000_0000;
array[38695] <= 16'b0000_0000_0000_0000;
array[38696] <= 16'b0000_0000_0000_0000;
array[38697] <= 16'b0000_0000_0000_0000;
array[38698] <= 16'b0000_0000_0000_0000;
array[38699] <= 16'b0000_0000_0000_0000;
array[38700] <= 16'b0000_0000_0000_0000;
array[38701] <= 16'b0000_0000_0000_0000;
array[38702] <= 16'b0000_0000_0000_0000;
array[38703] <= 16'b0000_0000_0000_0000;
array[38704] <= 16'b0000_0000_0000_0000;
array[38705] <= 16'b0000_0000_0000_0000;
array[38706] <= 16'b0000_0000_0000_0000;
array[38707] <= 16'b0000_0000_0000_0000;
array[38708] <= 16'b0000_0000_0000_0000;
array[38709] <= 16'b0000_0000_0000_0000;
array[38710] <= 16'b0000_0000_0000_0000;
array[38711] <= 16'b0000_0000_0000_0000;
array[38712] <= 16'b0000_0000_0000_0000;
array[38713] <= 16'b0000_0000_0000_0000;
array[38714] <= 16'b0000_0000_0000_0000;
array[38715] <= 16'b0000_0000_0000_0000;
array[38716] <= 16'b0000_0000_0000_0000;
array[38717] <= 16'b0000_0000_0000_0000;
array[38718] <= 16'b0000_0000_0000_0000;
array[38719] <= 16'b0000_0000_0000_0000;
array[38720] <= 16'b0000_0000_0000_0000;
array[38721] <= 16'b0000_0000_0000_0000;
array[38722] <= 16'b0000_0000_0000_0000;
array[38723] <= 16'b0000_0000_0000_0000;
array[38724] <= 16'b0000_0000_0000_0000;
array[38725] <= 16'b0000_0000_0000_0000;
array[38726] <= 16'b0000_0000_0000_0000;
array[38727] <= 16'b0000_0000_0000_0000;
array[38728] <= 16'b0000_0000_0000_0000;
array[38729] <= 16'b0000_0000_0000_0000;
array[38730] <= 16'b0000_0000_0000_0000;
array[38731] <= 16'b0000_0000_0000_0000;
array[38732] <= 16'b0000_0000_0000_0000;
array[38733] <= 16'b0000_0000_0000_0000;
array[38734] <= 16'b0000_0000_0000_0000;
array[38735] <= 16'b0000_0000_0000_0000;
array[38736] <= 16'b0000_0000_0000_0000;
array[38737] <= 16'b0000_0000_0000_0000;
array[38738] <= 16'b0000_0000_0000_0000;
array[38739] <= 16'b0000_0000_0000_0000;
array[38740] <= 16'b0000_0000_0000_0000;
array[38741] <= 16'b0000_0000_0000_0000;
array[38742] <= 16'b0000_0000_0000_0000;
array[38743] <= 16'b0000_0000_0000_0000;
array[38744] <= 16'b0000_0000_0000_0000;
array[38745] <= 16'b0000_0000_0000_0000;
array[38746] <= 16'b0000_0000_0000_0000;
array[38747] <= 16'b0000_0000_0000_0000;
array[38748] <= 16'b0000_0000_0000_0000;
array[38749] <= 16'b0000_0000_0000_0000;
array[38750] <= 16'b0000_0000_0000_0000;
array[38751] <= 16'b0000_0000_0000_0000;
array[38752] <= 16'b0000_0000_0000_0000;
array[38753] <= 16'b0000_0000_0000_0000;
array[38754] <= 16'b0000_0000_0000_0000;
array[38755] <= 16'b0000_0000_0000_0000;
array[38756] <= 16'b0000_0000_0000_0000;
array[38757] <= 16'b0000_0000_0000_0000;
array[38758] <= 16'b0000_0000_0000_0000;
array[38759] <= 16'b0000_0000_0000_0000;
array[38760] <= 16'b0000_0000_0000_0000;
array[38761] <= 16'b0000_0000_0000_0000;
array[38762] <= 16'b0000_0000_0000_0000;
array[38763] <= 16'b0000_0000_0000_0000;
array[38764] <= 16'b0000_0000_0000_0000;
array[38765] <= 16'b0000_0000_0000_0000;
array[38766] <= 16'b0000_0000_0000_0000;
array[38767] <= 16'b0000_0000_0000_0000;
array[38768] <= 16'b0000_0000_0000_0000;
array[38769] <= 16'b0000_0000_0000_0000;
array[38770] <= 16'b0000_0000_0000_0000;
array[38771] <= 16'b0000_0000_0000_0000;
array[38772] <= 16'b0000_0000_0000_0000;
array[38773] <= 16'b0000_0000_0000_0000;
array[38774] <= 16'b0000_0000_0000_0000;
array[38775] <= 16'b0000_0000_0000_0000;
array[38776] <= 16'b0000_0000_0000_0000;
array[38777] <= 16'b0000_0000_0000_0000;
array[38778] <= 16'b0000_0000_0000_0000;
array[38779] <= 16'b0000_0000_0000_0000;
array[38780] <= 16'b0000_0000_0000_0000;
array[38781] <= 16'b0000_0000_0000_0000;
array[38782] <= 16'b0000_0000_0000_0000;
array[38783] <= 16'b0000_0000_0000_0000;
array[38784] <= 16'b0000_0000_0000_0000;
array[38785] <= 16'b0000_0000_0000_0000;
array[38786] <= 16'b0000_0000_0000_0000;
array[38787] <= 16'b0000_0000_0000_0000;
array[38788] <= 16'b0000_0000_0000_0000;
array[38789] <= 16'b0000_0000_0000_0000;
array[38790] <= 16'b0000_0000_0000_0000;
array[38791] <= 16'b0000_0000_0000_0000;
array[38792] <= 16'b0000_0000_0000_0000;
array[38793] <= 16'b0000_0000_0000_0000;
array[38794] <= 16'b0000_0000_0000_0000;
array[38795] <= 16'b0000_0000_0000_0000;
array[38796] <= 16'b0000_0000_0000_0000;
array[38797] <= 16'b0000_0000_0000_0000;
array[38798] <= 16'b0000_0000_0000_0000;
array[38799] <= 16'b0000_0000_0000_0000;
array[38800] <= 16'b0000_0000_0000_0000;
array[38801] <= 16'b0000_0000_0000_0000;
array[38802] <= 16'b0000_0000_0000_0000;
array[38803] <= 16'b0000_0000_0000_0000;
array[38804] <= 16'b0000_0000_0000_0000;
array[38805] <= 16'b0000_0000_0000_0000;
array[38806] <= 16'b0000_0000_0000_0000;
array[38807] <= 16'b0000_0000_0000_0000;
array[38808] <= 16'b0000_0000_0000_0000;
array[38809] <= 16'b0000_0000_0000_0000;
array[38810] <= 16'b0000_0000_0000_0000;
array[38811] <= 16'b0000_0000_0000_0000;
array[38812] <= 16'b0000_0000_0000_0000;
array[38813] <= 16'b0000_0000_0000_0000;
array[38814] <= 16'b0000_0000_0000_0000;
array[38815] <= 16'b0000_0000_0000_0000;
array[38816] <= 16'b0000_0000_0000_0000;
array[38817] <= 16'b0000_0000_0000_0000;
array[38818] <= 16'b0000_0000_0000_0000;
array[38819] <= 16'b0000_0000_0000_0000;
array[38820] <= 16'b0000_0000_0000_0000;
array[38821] <= 16'b0000_0000_0000_0000;
array[38822] <= 16'b0000_0000_0000_0000;
array[38823] <= 16'b0000_0000_0000_0000;
array[38824] <= 16'b0000_0000_0000_0000;
array[38825] <= 16'b0000_0000_0000_0000;
array[38826] <= 16'b0000_0000_0000_0000;
array[38827] <= 16'b0000_0000_0000_0000;
array[38828] <= 16'b0000_0000_0000_0000;
array[38829] <= 16'b0000_0000_0000_0000;
array[38830] <= 16'b0000_0000_0000_0000;
array[38831] <= 16'b0000_0000_0000_0000;
array[38832] <= 16'b0000_0000_0000_0000;
array[38833] <= 16'b0000_0000_0000_0000;
array[38834] <= 16'b0000_0000_0000_0000;
array[38835] <= 16'b0000_0000_0000_0000;
array[38836] <= 16'b0000_0000_0000_0000;
array[38837] <= 16'b0000_0000_0000_0000;
array[38838] <= 16'b0000_0000_0000_0000;
array[38839] <= 16'b0000_0000_0000_0000;
array[38840] <= 16'b0000_0000_0000_0000;
array[38841] <= 16'b0000_0000_0000_0000;
array[38842] <= 16'b0000_0000_0000_0000;
array[38843] <= 16'b0000_0000_0000_0000;
array[38844] <= 16'b0000_0000_0000_0000;
array[38845] <= 16'b0000_0000_0000_0000;
array[38846] <= 16'b0000_0000_0000_0000;
array[38847] <= 16'b0000_0000_0000_0000;
array[38848] <= 16'b0000_0000_0000_0000;
array[38849] <= 16'b0000_0000_0000_0000;
array[38850] <= 16'b0000_0000_0000_0000;
array[38851] <= 16'b0000_0000_0000_0000;
array[38852] <= 16'b0000_0000_0000_0000;
array[38853] <= 16'b0000_0000_0000_0000;
array[38854] <= 16'b0000_0000_0000_0000;
array[38855] <= 16'b0000_0000_0000_0000;
array[38856] <= 16'b0000_0000_0000_0000;
array[38857] <= 16'b0000_0000_0000_0000;
array[38858] <= 16'b0000_0000_0000_0000;
array[38859] <= 16'b0000_0000_0000_0000;
array[38860] <= 16'b0000_0000_0000_0000;
array[38861] <= 16'b0000_0000_0000_0000;
array[38862] <= 16'b0000_0000_0000_0000;
array[38863] <= 16'b0000_0000_0000_0000;
array[38864] <= 16'b0000_0000_0000_0000;
array[38865] <= 16'b0000_0000_0000_0000;
array[38866] <= 16'b0000_0000_0000_0000;
array[38867] <= 16'b0000_0000_0000_0000;
array[38868] <= 16'b0000_0000_0000_0000;
array[38869] <= 16'b0000_0000_0000_0000;
array[38870] <= 16'b0000_0000_0000_0000;
array[38871] <= 16'b0000_0000_0000_0000;
array[38872] <= 16'b0000_0000_0000_0000;
array[38873] <= 16'b0000_0000_0000_0000;
array[38874] <= 16'b0000_0000_0000_0000;
array[38875] <= 16'b0000_0000_0000_0000;
array[38876] <= 16'b0000_0000_0000_0000;
array[38877] <= 16'b0000_0000_0000_0000;
array[38878] <= 16'b0000_0000_0000_0000;
array[38879] <= 16'b0000_0000_0000_0000;
array[38880] <= 16'b0000_0000_0000_0000;
array[38881] <= 16'b0000_0000_0000_0000;
array[38882] <= 16'b0000_0000_0000_0000;
array[38883] <= 16'b0000_0000_0000_0000;
array[38884] <= 16'b0000_0000_0000_0000;
array[38885] <= 16'b0000_0000_0000_0000;
array[38886] <= 16'b0000_0000_0000_0000;
array[38887] <= 16'b0000_0000_0000_0000;
array[38888] <= 16'b0000_0000_0000_0000;
array[38889] <= 16'b0000_0000_0000_0000;
array[38890] <= 16'b0000_0000_0000_0000;
array[38891] <= 16'b0000_0000_0000_0000;
array[38892] <= 16'b0000_0000_0000_0000;
array[38893] <= 16'b0000_0000_0000_0000;
array[38894] <= 16'b0000_0000_0000_0000;
array[38895] <= 16'b0000_0000_0000_0000;
array[38896] <= 16'b0000_0000_0000_0000;
array[38897] <= 16'b0000_0000_0000_0000;
array[38898] <= 16'b0000_0000_0000_0000;
array[38899] <= 16'b0000_0000_0000_0000;
array[38900] <= 16'b0000_0000_0000_0000;
array[38901] <= 16'b0000_0000_0000_0000;
array[38902] <= 16'b0000_0000_0000_0000;
array[38903] <= 16'b0000_0000_0000_0000;
array[38904] <= 16'b0000_0000_0000_0000;
array[38905] <= 16'b0000_0000_0000_0000;
array[38906] <= 16'b0000_0000_0000_0000;
array[38907] <= 16'b0000_0000_0000_0000;
array[38908] <= 16'b0000_0000_0000_0000;
array[38909] <= 16'b0000_0000_0000_0000;
array[38910] <= 16'b0000_0000_0000_0000;
array[38911] <= 16'b0000_0000_0000_0000;
array[38912] <= 16'b0000_0000_0000_0000;
array[38913] <= 16'b0000_0000_0000_0000;
array[38914] <= 16'b0000_0000_0000_0000;
array[38915] <= 16'b0000_0000_0000_0000;
array[38916] <= 16'b0000_0000_0000_0000;
array[38917] <= 16'b0000_0000_0000_0000;
array[38918] <= 16'b0000_0000_0000_0000;
array[38919] <= 16'b0000_0000_0000_0000;
array[38920] <= 16'b0000_0000_0000_0000;
array[38921] <= 16'b0000_0000_0000_0000;
array[38922] <= 16'b0000_0000_0000_0000;
array[38923] <= 16'b0000_0000_0000_0000;
array[38924] <= 16'b0000_0000_0000_0000;
array[38925] <= 16'b0000_0000_0000_0000;
array[38926] <= 16'b0000_0000_0000_0000;
array[38927] <= 16'b0000_0000_0000_0000;
array[38928] <= 16'b0000_0000_0000_0000;
array[38929] <= 16'b0000_0000_0000_0000;
array[38930] <= 16'b0000_0000_0000_0000;
array[38931] <= 16'b0000_0000_0000_0000;
array[38932] <= 16'b0000_0000_0000_0000;
array[38933] <= 16'b0000_0000_0000_0000;
array[38934] <= 16'b0000_0000_0000_0000;
array[38935] <= 16'b0000_0000_0000_0000;
array[38936] <= 16'b0000_0000_0000_0000;
array[38937] <= 16'b0000_0000_0000_0000;
array[38938] <= 16'b0000_0000_0000_0000;
array[38939] <= 16'b0000_0000_0000_0000;
array[38940] <= 16'b0000_0000_0000_0000;
array[38941] <= 16'b0000_0000_0000_0000;
array[38942] <= 16'b0000_0000_0000_0000;
array[38943] <= 16'b0000_0000_0000_0000;
array[38944] <= 16'b0000_0000_0000_0000;
array[38945] <= 16'b0000_0000_0000_0000;
array[38946] <= 16'b0000_0000_0000_0000;
array[38947] <= 16'b0000_0000_0000_0000;
array[38948] <= 16'b0000_0000_0000_0000;
array[38949] <= 16'b0000_0000_0000_0000;
array[38950] <= 16'b0000_0000_0000_0000;
array[38951] <= 16'b0000_0000_0000_0000;
array[38952] <= 16'b0000_0000_0000_0000;
array[38953] <= 16'b0000_0000_0000_0000;
array[38954] <= 16'b0000_0000_0000_0000;
array[38955] <= 16'b0000_0000_0000_0000;
array[38956] <= 16'b0000_0000_0000_0000;
array[38957] <= 16'b0000_0000_0000_0000;
array[38958] <= 16'b0000_0000_0000_0000;
array[38959] <= 16'b0000_0000_0000_0000;
array[38960] <= 16'b0000_0000_0000_0000;
array[38961] <= 16'b0000_0000_0000_0000;
array[38962] <= 16'b0000_0000_0000_0000;
array[38963] <= 16'b0000_0000_0000_0000;
array[38964] <= 16'b0000_0000_0000_0000;
array[38965] <= 16'b0000_0000_0000_0000;
array[38966] <= 16'b0000_0000_0000_0000;
array[38967] <= 16'b0000_0000_0000_0000;
array[38968] <= 16'b0000_0000_0000_0000;
array[38969] <= 16'b0000_0000_0000_0000;
array[38970] <= 16'b0000_0000_0000_0000;
array[38971] <= 16'b0000_0000_0000_0000;
array[38972] <= 16'b0000_0000_0000_0000;
array[38973] <= 16'b0000_0000_0000_0000;
array[38974] <= 16'b0000_0000_0000_0000;
array[38975] <= 16'b0000_0000_0000_0000;
array[38976] <= 16'b0000_0000_0000_0000;
array[38977] <= 16'b0000_0000_0000_0000;
array[38978] <= 16'b0000_0000_0000_0000;
array[38979] <= 16'b0000_0000_0000_0000;
array[38980] <= 16'b0000_0000_0000_0000;
array[38981] <= 16'b0000_0000_0000_0000;
array[38982] <= 16'b0000_0000_0000_0000;
array[38983] <= 16'b0000_0000_0000_0000;
array[38984] <= 16'b0000_0000_0000_0000;
array[38985] <= 16'b0000_0000_0000_0000;
array[38986] <= 16'b0000_0000_0000_0000;
array[38987] <= 16'b0000_0000_0000_0000;
array[38988] <= 16'b0000_0000_0000_0000;
array[38989] <= 16'b0000_0000_0000_0000;
array[38990] <= 16'b0000_0000_0000_0000;
array[38991] <= 16'b0000_0000_0000_0000;
array[38992] <= 16'b0000_0000_0000_0000;
array[38993] <= 16'b0000_0000_0000_0000;
array[38994] <= 16'b0000_0000_0000_0000;
array[38995] <= 16'b0000_0000_0000_0000;
array[38996] <= 16'b0000_0000_0000_0000;
array[38997] <= 16'b0000_0000_0000_0000;
array[38998] <= 16'b0000_0000_0000_0000;
array[38999] <= 16'b0000_0000_0000_0000;
array[39000] <= 16'b0000_0000_0000_0000;
array[39001] <= 16'b0000_0000_0000_0000;
array[39002] <= 16'b0000_0000_0000_0000;
array[39003] <= 16'b0000_0000_0000_0000;
array[39004] <= 16'b0000_0000_0000_0000;
array[39005] <= 16'b0000_0000_0000_0000;
array[39006] <= 16'b0000_0000_0000_0000;
array[39007] <= 16'b0000_0000_0000_0000;
array[39008] <= 16'b0000_0000_0000_0000;
array[39009] <= 16'b0000_0000_0000_0000;
array[39010] <= 16'b0000_0000_0000_0000;
array[39011] <= 16'b0000_0000_0000_0000;
array[39012] <= 16'b0000_0000_0000_0000;
array[39013] <= 16'b0000_0000_0000_0000;
array[39014] <= 16'b0000_0000_0000_0000;
array[39015] <= 16'b0000_0000_0000_0000;
array[39016] <= 16'b0000_0000_0000_0000;
array[39017] <= 16'b0000_0000_0000_0000;
array[39018] <= 16'b0000_0000_0000_0000;
array[39019] <= 16'b0000_0000_0000_0000;
array[39020] <= 16'b0000_0000_0000_0000;
array[39021] <= 16'b0000_0000_0000_0000;
array[39022] <= 16'b0000_0000_0000_0000;
array[39023] <= 16'b0000_0000_0000_0000;
array[39024] <= 16'b0000_0000_0000_0000;
array[39025] <= 16'b0000_0000_0000_0000;
array[39026] <= 16'b0000_0000_0000_0000;
array[39027] <= 16'b0000_0000_0000_0000;
array[39028] <= 16'b0000_0000_0000_0000;
array[39029] <= 16'b0000_0000_0000_0000;
array[39030] <= 16'b0000_0000_0000_0000;
array[39031] <= 16'b0000_0000_0000_0000;
array[39032] <= 16'b0000_0000_0000_0000;
array[39033] <= 16'b0000_0000_0000_0000;
array[39034] <= 16'b0000_0000_0000_0000;
array[39035] <= 16'b0000_0000_0000_0000;
array[39036] <= 16'b0000_0000_0000_0000;
array[39037] <= 16'b0000_0000_0000_0000;
array[39038] <= 16'b0000_0000_0000_0000;
array[39039] <= 16'b0000_0000_0000_0000;
array[39040] <= 16'b0000_0000_0000_0000;
array[39041] <= 16'b0000_0000_0000_0000;
array[39042] <= 16'b0000_0000_0000_0000;
array[39043] <= 16'b0000_0000_0000_0000;
array[39044] <= 16'b0000_0000_0000_0000;
array[39045] <= 16'b0000_0000_0000_0000;
array[39046] <= 16'b0000_0000_0000_0000;
array[39047] <= 16'b0000_0000_0000_0000;
array[39048] <= 16'b0000_0000_0000_0000;
array[39049] <= 16'b0000_0000_0000_0000;
array[39050] <= 16'b0000_0000_0000_0000;
array[39051] <= 16'b0000_0000_0000_0000;
array[39052] <= 16'b0000_0000_0000_0000;
array[39053] <= 16'b0000_0000_0000_0000;
array[39054] <= 16'b0000_0000_0000_0000;
array[39055] <= 16'b0000_0000_0000_0000;
array[39056] <= 16'b0000_0000_0000_0000;
array[39057] <= 16'b0000_0000_0000_0000;
array[39058] <= 16'b0000_0000_0000_0000;
array[39059] <= 16'b0000_0000_0000_0000;
array[39060] <= 16'b0000_0000_0000_0000;
array[39061] <= 16'b0000_0000_0000_0000;
array[39062] <= 16'b0000_0000_0000_0000;
array[39063] <= 16'b0000_0000_0000_0000;
array[39064] <= 16'b0000_0000_0000_0000;
array[39065] <= 16'b0000_0000_0000_0000;
array[39066] <= 16'b0000_0000_0000_0000;
array[39067] <= 16'b0000_0000_0000_0000;
array[39068] <= 16'b0000_0000_0000_0000;
array[39069] <= 16'b0000_0000_0000_0000;
array[39070] <= 16'b0000_0000_0000_0000;
array[39071] <= 16'b0000_0000_0000_0000;
array[39072] <= 16'b0000_0000_0000_0000;
array[39073] <= 16'b0000_0000_0000_0000;
array[39074] <= 16'b0000_0000_0000_0000;
array[39075] <= 16'b0000_0000_0000_0000;
array[39076] <= 16'b0000_0000_0000_0000;
array[39077] <= 16'b0000_0000_0000_0000;
array[39078] <= 16'b0000_0000_0000_0000;
array[39079] <= 16'b0000_0000_0000_0000;
array[39080] <= 16'b0000_0000_0000_0000;
array[39081] <= 16'b0000_0000_0000_0000;
array[39082] <= 16'b0000_0000_0000_0000;
array[39083] <= 16'b0000_0000_0000_0000;
array[39084] <= 16'b0000_0000_0000_0000;
array[39085] <= 16'b0000_0000_0000_0000;
array[39086] <= 16'b0000_0000_0000_0000;
array[39087] <= 16'b0000_0000_0000_0000;
array[39088] <= 16'b0000_0000_0000_0000;
array[39089] <= 16'b0000_0000_0000_0000;
array[39090] <= 16'b0000_0000_0000_0000;
array[39091] <= 16'b0000_0000_0000_0000;
array[39092] <= 16'b0000_0000_0000_0000;
array[39093] <= 16'b0000_0000_0000_0000;
array[39094] <= 16'b0000_0000_0000_0000;
array[39095] <= 16'b0000_0000_0000_0000;
array[39096] <= 16'b0000_0000_0000_0000;
array[39097] <= 16'b0000_0000_0000_0000;
array[39098] <= 16'b0000_0000_0000_0000;
array[39099] <= 16'b0000_0000_0000_0000;
array[39100] <= 16'b0000_0000_0000_0000;
array[39101] <= 16'b0000_0000_0000_0000;
array[39102] <= 16'b0000_0000_0000_0000;
array[39103] <= 16'b0000_0000_0000_0000;
array[39104] <= 16'b0000_0000_0000_0000;
array[39105] <= 16'b0000_0000_0000_0000;
array[39106] <= 16'b0000_0000_0000_0000;
array[39107] <= 16'b0000_0000_0000_0000;
array[39108] <= 16'b0000_0000_0000_0000;
array[39109] <= 16'b0000_0000_0000_0000;
array[39110] <= 16'b0000_0000_0000_0000;
array[39111] <= 16'b0000_0000_0000_0000;
array[39112] <= 16'b0000_0000_0000_0000;
array[39113] <= 16'b0000_0000_0000_0000;
array[39114] <= 16'b0000_0000_0000_0000;
array[39115] <= 16'b0000_0000_0000_0000;
array[39116] <= 16'b0000_0000_0000_0000;
array[39117] <= 16'b0000_0000_0000_0000;
array[39118] <= 16'b0000_0000_0000_0000;
array[39119] <= 16'b0000_0000_0000_0000;
array[39120] <= 16'b0000_0000_0000_0000;
array[39121] <= 16'b0000_0000_0000_0000;
array[39122] <= 16'b0000_0000_0000_0000;
array[39123] <= 16'b0000_0000_0000_0000;
array[39124] <= 16'b0000_0000_0000_0000;
array[39125] <= 16'b0000_0000_0000_0000;
array[39126] <= 16'b0000_0000_0000_0000;
array[39127] <= 16'b0000_0000_0000_0000;
array[39128] <= 16'b0000_0000_0000_0000;
array[39129] <= 16'b0000_0000_0000_0000;
array[39130] <= 16'b0000_0000_0000_0000;
array[39131] <= 16'b0000_0000_0000_0000;
array[39132] <= 16'b0000_0000_0000_0000;
array[39133] <= 16'b0000_0000_0000_0000;
array[39134] <= 16'b0000_0000_0000_0000;
array[39135] <= 16'b0000_0000_0000_0000;
array[39136] <= 16'b0000_0000_0000_0000;
array[39137] <= 16'b0000_0000_0000_0000;
array[39138] <= 16'b0000_0000_0000_0000;
array[39139] <= 16'b0000_0000_0000_0000;
array[39140] <= 16'b0000_0000_0000_0000;
array[39141] <= 16'b0000_0000_0000_0000;
array[39142] <= 16'b0000_0000_0000_0000;
array[39143] <= 16'b0000_0000_0000_0000;
array[39144] <= 16'b0000_0000_0000_0000;
array[39145] <= 16'b0000_0000_0000_0000;
array[39146] <= 16'b0000_0000_0000_0000;
array[39147] <= 16'b0000_0000_0000_0000;
array[39148] <= 16'b0000_0000_0000_0000;
array[39149] <= 16'b0000_0000_0000_0000;
array[39150] <= 16'b0000_0000_0000_0000;
array[39151] <= 16'b0000_0000_0000_0000;
array[39152] <= 16'b0000_0000_0000_0000;
array[39153] <= 16'b0000_0000_0000_0000;
array[39154] <= 16'b0000_0000_0000_0000;
array[39155] <= 16'b0000_0000_0000_0000;
array[39156] <= 16'b0000_0000_0000_0000;
array[39157] <= 16'b0000_0000_0000_0000;
array[39158] <= 16'b0000_0000_0000_0000;
array[39159] <= 16'b0000_0000_0000_0000;
array[39160] <= 16'b0000_0000_0000_0000;
array[39161] <= 16'b0000_0000_0000_0000;
array[39162] <= 16'b0000_0000_0000_0000;
array[39163] <= 16'b0000_0000_0000_0000;
array[39164] <= 16'b0000_0000_0000_0000;
array[39165] <= 16'b0000_0000_0000_0000;
array[39166] <= 16'b0000_0000_0000_0000;
array[39167] <= 16'b0000_0000_0000_0000;
array[39168] <= 16'b0000_0000_0000_0000;
array[39169] <= 16'b0000_0000_0000_0000;
array[39170] <= 16'b0000_0000_0000_0000;
array[39171] <= 16'b0000_0000_0000_0000;
array[39172] <= 16'b0000_0000_0000_0000;
array[39173] <= 16'b0000_0000_0000_0000;
array[39174] <= 16'b0000_0000_0000_0000;
array[39175] <= 16'b0000_0000_0000_0000;
array[39176] <= 16'b0000_0000_0000_0000;
array[39177] <= 16'b0000_0000_0000_0000;
array[39178] <= 16'b0000_0000_0000_0000;
array[39179] <= 16'b0000_0000_0000_0000;
array[39180] <= 16'b0000_0000_0000_0000;
array[39181] <= 16'b0000_0000_0000_0000;
array[39182] <= 16'b0000_0000_0000_0000;
array[39183] <= 16'b0000_0000_0000_0000;
array[39184] <= 16'b0000_0000_0000_0000;
array[39185] <= 16'b0000_0000_0000_0000;
array[39186] <= 16'b0000_0000_0000_0000;
array[39187] <= 16'b0000_0000_0000_0000;
array[39188] <= 16'b0000_0000_0000_0000;
array[39189] <= 16'b0000_0000_0000_0000;
array[39190] <= 16'b0000_0000_0000_0000;
array[39191] <= 16'b0000_0000_0000_0000;
array[39192] <= 16'b0000_0000_0000_0000;
array[39193] <= 16'b0000_0000_0000_0000;
array[39194] <= 16'b0000_0000_0000_0000;
array[39195] <= 16'b0000_0000_0000_0000;
array[39196] <= 16'b0000_0000_0000_0000;
array[39197] <= 16'b0000_0000_0000_0000;
array[39198] <= 16'b0000_0000_0000_0000;
array[39199] <= 16'b0000_0000_0000_0000;
array[39200] <= 16'b0000_0000_0000_0000;
array[39201] <= 16'b0000_0000_0000_0000;
array[39202] <= 16'b0000_0000_0000_0000;
array[39203] <= 16'b0000_0000_0000_0000;
array[39204] <= 16'b0000_0000_0000_0000;
array[39205] <= 16'b0000_0000_0000_0000;
array[39206] <= 16'b0000_0000_0000_0000;
array[39207] <= 16'b0000_0000_0000_0000;
array[39208] <= 16'b0000_0000_0000_0000;
array[39209] <= 16'b0000_0000_0000_0000;
array[39210] <= 16'b0000_0000_0000_0000;
array[39211] <= 16'b0000_0000_0000_0000;
array[39212] <= 16'b0000_0000_0000_0000;
array[39213] <= 16'b0000_0000_0000_0000;
array[39214] <= 16'b0000_0000_0000_0000;
array[39215] <= 16'b0000_0000_0000_0000;
array[39216] <= 16'b0000_0000_0000_0000;
array[39217] <= 16'b0000_0000_0000_0000;
array[39218] <= 16'b0000_0000_0000_0000;
array[39219] <= 16'b0000_0000_0000_0000;
array[39220] <= 16'b0000_0000_0000_0000;
array[39221] <= 16'b0000_0000_0000_0000;
array[39222] <= 16'b0000_0000_0000_0000;
array[39223] <= 16'b0000_0000_0000_0000;
array[39224] <= 16'b0000_0000_0000_0000;
array[39225] <= 16'b0000_0000_0000_0000;
array[39226] <= 16'b0000_0000_0000_0000;
array[39227] <= 16'b0000_0000_0000_0000;
array[39228] <= 16'b0000_0000_0000_0000;
array[39229] <= 16'b0000_0000_0000_0000;
array[39230] <= 16'b0000_0000_0000_0000;
array[39231] <= 16'b0000_0000_0000_0000;
array[39232] <= 16'b0000_0000_0000_0000;
array[39233] <= 16'b0000_0000_0000_0000;
array[39234] <= 16'b0000_0000_0000_0000;
array[39235] <= 16'b0000_0000_0000_0000;
array[39236] <= 16'b0000_0000_0000_0000;
array[39237] <= 16'b0000_0000_0000_0000;
array[39238] <= 16'b0000_0000_0000_0000;
array[39239] <= 16'b0000_0000_0000_0000;
array[39240] <= 16'b0000_0000_0000_0000;
array[39241] <= 16'b0000_0000_0000_0000;
array[39242] <= 16'b0000_0000_0000_0000;
array[39243] <= 16'b0000_0000_0000_0000;
array[39244] <= 16'b0000_0000_0000_0000;
array[39245] <= 16'b0000_0000_0000_0000;
array[39246] <= 16'b0000_0000_0000_0000;
array[39247] <= 16'b0000_0000_0000_0000;
array[39248] <= 16'b0000_0000_0000_0000;
array[39249] <= 16'b0000_0000_0000_0000;
array[39250] <= 16'b0000_0000_0000_0000;
array[39251] <= 16'b0000_0000_0000_0000;
array[39252] <= 16'b0000_0000_0000_0000;
array[39253] <= 16'b0000_0000_0000_0000;
array[39254] <= 16'b0000_0000_0000_0000;
array[39255] <= 16'b0000_0000_0000_0000;
array[39256] <= 16'b0000_0000_0000_0000;
array[39257] <= 16'b0000_0000_0000_0000;
array[39258] <= 16'b0000_0000_0000_0000;
array[39259] <= 16'b0000_0000_0000_0000;
array[39260] <= 16'b0000_0000_0000_0000;
array[39261] <= 16'b0000_0000_0000_0000;
array[39262] <= 16'b0000_0000_0000_0000;
array[39263] <= 16'b0000_0000_0000_0000;
array[39264] <= 16'b0000_0000_0000_0000;
array[39265] <= 16'b0000_0000_0000_0000;
array[39266] <= 16'b0000_0000_0000_0000;
array[39267] <= 16'b0000_0000_0000_0000;
array[39268] <= 16'b0000_0000_0000_0000;
array[39269] <= 16'b0000_0000_0000_0000;
array[39270] <= 16'b0000_0000_0000_0000;
array[39271] <= 16'b0000_0000_0000_0000;
array[39272] <= 16'b0000_0000_0000_0000;
array[39273] <= 16'b0000_0000_0000_0000;
array[39274] <= 16'b0000_0000_0000_0000;
array[39275] <= 16'b0000_0000_0000_0000;
array[39276] <= 16'b0000_0000_0000_0000;
array[39277] <= 16'b0000_0000_0000_0000;
array[39278] <= 16'b0000_0000_0000_0000;
array[39279] <= 16'b0000_0000_0000_0000;
array[39280] <= 16'b0000_0000_0000_0000;
array[39281] <= 16'b0000_0000_0000_0000;
array[39282] <= 16'b0000_0000_0000_0000;
array[39283] <= 16'b0000_0000_0000_0000;
array[39284] <= 16'b0000_0000_0000_0000;
array[39285] <= 16'b0000_0000_0000_0000;
array[39286] <= 16'b0000_0000_0000_0000;
array[39287] <= 16'b0000_0000_0000_0000;
array[39288] <= 16'b0000_0000_0000_0000;
array[39289] <= 16'b0000_0000_0000_0000;
array[39290] <= 16'b0000_0000_0000_0000;
array[39291] <= 16'b0000_0000_0000_0000;
array[39292] <= 16'b0000_0000_0000_0000;
array[39293] <= 16'b0000_0000_0000_0000;
array[39294] <= 16'b0000_0000_0000_0000;
array[39295] <= 16'b0000_0000_0000_0000;
array[39296] <= 16'b0000_0000_0000_0000;
array[39297] <= 16'b0000_0000_0000_0000;
array[39298] <= 16'b0000_0000_0000_0000;
array[39299] <= 16'b0000_0000_0000_0000;
array[39300] <= 16'b0000_0000_0000_0000;
array[39301] <= 16'b0000_0000_0000_0000;
array[39302] <= 16'b0000_0000_0000_0000;
array[39303] <= 16'b0000_0000_0000_0000;
array[39304] <= 16'b0000_0000_0000_0000;
array[39305] <= 16'b0000_0000_0000_0000;
array[39306] <= 16'b0000_0000_0000_0000;
array[39307] <= 16'b0000_0000_0000_0000;
array[39308] <= 16'b0000_0000_0000_0000;
array[39309] <= 16'b0000_0000_0000_0000;
array[39310] <= 16'b0000_0000_0000_0000;
array[39311] <= 16'b0000_0000_0000_0000;
array[39312] <= 16'b0000_0000_0000_0000;
array[39313] <= 16'b0000_0000_0000_0000;
array[39314] <= 16'b0000_0000_0000_0000;
array[39315] <= 16'b0000_0000_0000_0000;
array[39316] <= 16'b0000_0000_0000_0000;
array[39317] <= 16'b0000_0000_0000_0000;
array[39318] <= 16'b0000_0000_0000_0000;
array[39319] <= 16'b0000_0000_0000_0000;
array[39320] <= 16'b0000_0000_0000_0000;
array[39321] <= 16'b0000_0000_0000_0000;
array[39322] <= 16'b0000_0000_0000_0000;
array[39323] <= 16'b0000_0000_0000_0000;
array[39324] <= 16'b0000_0000_0000_0000;
array[39325] <= 16'b0000_0000_0000_0000;
array[39326] <= 16'b0000_0000_0000_0000;
array[39327] <= 16'b0000_0000_0000_0000;
array[39328] <= 16'b0000_0000_0000_0000;
array[39329] <= 16'b0000_0000_0000_0000;
array[39330] <= 16'b0000_0000_0000_0000;
array[39331] <= 16'b0000_0000_0000_0000;
array[39332] <= 16'b0000_0000_0000_0000;
array[39333] <= 16'b0000_0000_0000_0000;
array[39334] <= 16'b0000_0000_0000_0000;
array[39335] <= 16'b0000_0000_0000_0000;
array[39336] <= 16'b0000_0000_0000_0000;
array[39337] <= 16'b0000_0000_0000_0000;
array[39338] <= 16'b0000_0000_0000_0000;
array[39339] <= 16'b0000_0000_0000_0000;
array[39340] <= 16'b0000_0000_0000_0000;
array[39341] <= 16'b0000_0000_0000_0000;
array[39342] <= 16'b0000_0000_0000_0000;
array[39343] <= 16'b0000_0000_0000_0000;
array[39344] <= 16'b0000_0000_0000_0000;
array[39345] <= 16'b0000_0000_0000_0000;
array[39346] <= 16'b0000_0000_0000_0000;
array[39347] <= 16'b0000_0000_0000_0000;
array[39348] <= 16'b0000_0000_0000_0000;
array[39349] <= 16'b0000_0000_0000_0000;
array[39350] <= 16'b0000_0000_0000_0000;
array[39351] <= 16'b0000_0000_0000_0000;
array[39352] <= 16'b0000_0000_0000_0000;
array[39353] <= 16'b0000_0000_0000_0000;
array[39354] <= 16'b0000_0000_0000_0000;
array[39355] <= 16'b0000_0000_0000_0000;
array[39356] <= 16'b0000_0000_0000_0000;
array[39357] <= 16'b0000_0000_0000_0000;
array[39358] <= 16'b0000_0000_0000_0000;
array[39359] <= 16'b0000_0000_0000_0000;
array[39360] <= 16'b0000_0000_0000_0000;
array[39361] <= 16'b0000_0000_0000_0000;
array[39362] <= 16'b0000_0000_0000_0000;
array[39363] <= 16'b0000_0000_0000_0000;
array[39364] <= 16'b0000_0000_0000_0000;
array[39365] <= 16'b0000_0000_0000_0000;
array[39366] <= 16'b0000_0000_0000_0000;
array[39367] <= 16'b0000_0000_0000_0000;
array[39368] <= 16'b0000_0000_0000_0000;
array[39369] <= 16'b0000_0000_0000_0000;
array[39370] <= 16'b0000_0000_0000_0000;
array[39371] <= 16'b0000_0000_0000_0000;
array[39372] <= 16'b0000_0000_0000_0000;
array[39373] <= 16'b0000_0000_0000_0000;
array[39374] <= 16'b0000_0000_0000_0000;
array[39375] <= 16'b0000_0000_0000_0000;
array[39376] <= 16'b0000_0000_0000_0000;
array[39377] <= 16'b0000_0000_0000_0000;
array[39378] <= 16'b0000_0000_0000_0000;
array[39379] <= 16'b0000_0000_0000_0000;
array[39380] <= 16'b0000_0000_0000_0000;
array[39381] <= 16'b0000_0000_0000_0000;
array[39382] <= 16'b0000_0000_0000_0000;
array[39383] <= 16'b0000_0000_0000_0000;
array[39384] <= 16'b0000_0000_0000_0000;
array[39385] <= 16'b0000_0000_0000_0000;
array[39386] <= 16'b0000_0000_0000_0000;
array[39387] <= 16'b0000_0000_0000_0000;
array[39388] <= 16'b0000_0000_0000_0000;
array[39389] <= 16'b0000_0000_0000_0000;
array[39390] <= 16'b0000_0000_0000_0000;
array[39391] <= 16'b0000_0000_0000_0000;
array[39392] <= 16'b0000_0000_0000_0000;
array[39393] <= 16'b0000_0000_0000_0000;
array[39394] <= 16'b0000_0000_0000_0000;
array[39395] <= 16'b0000_0000_0000_0000;
array[39396] <= 16'b0000_0000_0000_0000;
array[39397] <= 16'b0000_0000_0000_0000;
array[39398] <= 16'b0000_0000_0000_0000;
array[39399] <= 16'b0000_0000_0000_0000;
array[39400] <= 16'b0000_0000_0000_0000;
array[39401] <= 16'b0000_0000_0000_0000;
array[39402] <= 16'b0000_0000_0000_0000;
array[39403] <= 16'b0000_0000_0000_0000;
array[39404] <= 16'b0000_0000_0000_0000;
array[39405] <= 16'b0000_0000_0000_0000;
array[39406] <= 16'b0000_0000_0000_0000;
array[39407] <= 16'b0000_0000_0000_0000;
array[39408] <= 16'b0000_0000_0000_0000;
array[39409] <= 16'b0000_0000_0000_0000;
array[39410] <= 16'b0000_0000_0000_0000;
array[39411] <= 16'b0000_0000_0000_0000;
array[39412] <= 16'b0000_0000_0000_0000;
array[39413] <= 16'b0000_0000_0000_0000;
array[39414] <= 16'b0000_0000_0000_0000;
array[39415] <= 16'b0000_0000_0000_0000;
array[39416] <= 16'b0000_0000_0000_0000;
array[39417] <= 16'b0000_0000_0000_0000;
array[39418] <= 16'b0000_0000_0000_0000;
array[39419] <= 16'b0000_0000_0000_0000;
array[39420] <= 16'b0000_0000_0000_0000;
array[39421] <= 16'b0000_0000_0000_0000;
array[39422] <= 16'b0000_0000_0000_0000;
array[39423] <= 16'b0000_0000_0000_0000;
array[39424] <= 16'b0000_0000_0000_0000;
array[39425] <= 16'b0000_0000_0000_0000;
array[39426] <= 16'b0000_0000_0000_0000;
array[39427] <= 16'b0000_0000_0000_0000;
array[39428] <= 16'b0000_0000_0000_0000;
array[39429] <= 16'b0000_0000_0000_0000;
array[39430] <= 16'b0000_0000_0000_0000;
array[39431] <= 16'b0000_0000_0000_0000;
array[39432] <= 16'b0000_0000_0000_0000;
array[39433] <= 16'b0000_0000_0000_0000;
array[39434] <= 16'b0000_0000_0000_0000;
array[39435] <= 16'b0000_0000_0000_0000;
array[39436] <= 16'b0000_0000_0000_0000;
array[39437] <= 16'b0000_0000_0000_0000;
array[39438] <= 16'b0000_0000_0000_0000;
array[39439] <= 16'b0000_0000_0000_0000;
array[39440] <= 16'b0000_0000_0000_0000;
array[39441] <= 16'b0000_0000_0000_0000;
array[39442] <= 16'b0000_0000_0000_0000;
array[39443] <= 16'b0000_0000_0000_0000;
array[39444] <= 16'b0000_0000_0000_0000;
array[39445] <= 16'b0000_0000_0000_0000;
array[39446] <= 16'b0000_0000_0000_0000;
array[39447] <= 16'b0000_0000_0000_0000;
array[39448] <= 16'b0000_0000_0000_0000;
array[39449] <= 16'b0000_0000_0000_0000;
array[39450] <= 16'b0000_0000_0000_0000;
array[39451] <= 16'b0000_0000_0000_0000;
array[39452] <= 16'b0000_0000_0000_0000;
array[39453] <= 16'b0000_0000_0000_0000;
array[39454] <= 16'b0000_0000_0000_0000;
array[39455] <= 16'b0000_0000_0000_0000;
array[39456] <= 16'b0000_0000_0000_0000;
array[39457] <= 16'b0000_0000_0000_0000;
array[39458] <= 16'b0000_0000_0000_0000;
array[39459] <= 16'b0000_0000_0000_0000;
array[39460] <= 16'b0000_0000_0000_0000;
array[39461] <= 16'b0000_0000_0000_0000;
array[39462] <= 16'b0000_0000_0000_0000;
array[39463] <= 16'b0000_0000_0000_0000;
array[39464] <= 16'b0000_0000_0000_0000;
array[39465] <= 16'b0000_0000_0000_0000;
array[39466] <= 16'b0000_0000_0000_0000;
array[39467] <= 16'b0000_0000_0000_0000;
array[39468] <= 16'b0000_0000_0000_0000;
array[39469] <= 16'b0000_0000_0000_0000;
array[39470] <= 16'b0000_0000_0000_0000;
array[39471] <= 16'b0000_0000_0000_0000;
array[39472] <= 16'b0000_0000_0000_0000;
array[39473] <= 16'b0000_0000_0000_0000;
array[39474] <= 16'b0000_0000_0000_0000;
array[39475] <= 16'b0000_0000_0000_0000;
array[39476] <= 16'b0000_0000_0000_0000;
array[39477] <= 16'b0000_0000_0000_0000;
array[39478] <= 16'b0000_0000_0000_0000;
array[39479] <= 16'b0000_0000_0000_0000;
array[39480] <= 16'b0000_0000_0000_0000;
array[39481] <= 16'b0000_0000_0000_0000;
array[39482] <= 16'b0000_0000_0000_0000;
array[39483] <= 16'b0000_0000_0000_0000;
array[39484] <= 16'b0000_0000_0000_0000;
array[39485] <= 16'b0000_0000_0000_0000;
array[39486] <= 16'b0000_0000_0000_0000;
array[39487] <= 16'b0000_0000_0000_0000;
array[39488] <= 16'b0000_0000_0000_0000;
array[39489] <= 16'b0000_0000_0000_0000;
array[39490] <= 16'b0000_0000_0000_0000;
array[39491] <= 16'b0000_0000_0000_0000;
array[39492] <= 16'b0000_0000_0000_0000;
array[39493] <= 16'b0000_0000_0000_0000;
array[39494] <= 16'b0000_0000_0000_0000;
array[39495] <= 16'b0000_0000_0000_0000;
array[39496] <= 16'b0000_0000_0000_0000;
array[39497] <= 16'b0000_0000_0000_0000;
array[39498] <= 16'b0000_0000_0000_0000;
array[39499] <= 16'b0000_0000_0000_0000;
array[39500] <= 16'b0000_0000_0000_0000;
array[39501] <= 16'b0000_0000_0000_0000;
array[39502] <= 16'b0000_0000_0000_0000;
array[39503] <= 16'b0000_0000_0000_0000;
array[39504] <= 16'b0000_0000_0000_0000;
array[39505] <= 16'b0000_0000_0000_0000;
array[39506] <= 16'b0000_0000_0000_0000;
array[39507] <= 16'b0000_0000_0000_0000;
array[39508] <= 16'b0000_0000_0000_0000;
array[39509] <= 16'b0000_0000_0000_0000;
array[39510] <= 16'b0000_0000_0000_0000;
array[39511] <= 16'b0000_0000_0000_0000;
array[39512] <= 16'b0000_0000_0000_0000;
array[39513] <= 16'b0000_0000_0000_0000;
array[39514] <= 16'b0000_0000_0000_0000;
array[39515] <= 16'b0000_0000_0000_0000;
array[39516] <= 16'b0000_0000_0000_0000;
array[39517] <= 16'b0000_0000_0000_0000;
array[39518] <= 16'b0000_0000_0000_0000;
array[39519] <= 16'b0000_0000_0000_0000;
array[39520] <= 16'b0000_0000_0000_0000;
array[39521] <= 16'b0000_0000_0000_0000;
array[39522] <= 16'b0000_0000_0000_0000;
array[39523] <= 16'b0000_0000_0000_0000;
array[39524] <= 16'b0000_0000_0000_0000;
array[39525] <= 16'b0000_0000_0000_0000;
array[39526] <= 16'b0000_0000_0000_0000;
array[39527] <= 16'b0000_0000_0000_0000;
array[39528] <= 16'b0000_0000_0000_0000;
array[39529] <= 16'b0000_0000_0000_0000;
array[39530] <= 16'b0000_0000_0000_0000;
array[39531] <= 16'b0000_0000_0000_0000;
array[39532] <= 16'b0000_0000_0000_0000;
array[39533] <= 16'b0000_0000_0000_0000;
array[39534] <= 16'b0000_0000_0000_0000;
array[39535] <= 16'b0000_0000_0000_0000;
array[39536] <= 16'b0000_0000_0000_0000;
array[39537] <= 16'b0000_0000_0000_0000;
array[39538] <= 16'b0000_0000_0000_0000;
array[39539] <= 16'b0000_0000_0000_0000;
array[39540] <= 16'b0000_0000_0000_0000;
array[39541] <= 16'b0000_0000_0000_0000;
array[39542] <= 16'b0000_0000_0000_0000;
array[39543] <= 16'b0000_0000_0000_0000;
array[39544] <= 16'b0000_0000_0000_0000;
array[39545] <= 16'b0000_0000_0000_0000;
array[39546] <= 16'b0000_0000_0000_0000;
array[39547] <= 16'b0000_0000_0000_0000;
array[39548] <= 16'b0000_0000_0000_0000;
array[39549] <= 16'b0000_0000_0000_0000;
array[39550] <= 16'b0000_0000_0000_0000;
array[39551] <= 16'b0000_0000_0000_0000;
array[39552] <= 16'b0000_0000_0000_0000;
array[39553] <= 16'b0000_0000_0000_0000;
array[39554] <= 16'b0000_0000_0000_0000;
array[39555] <= 16'b0000_0000_0000_0000;
array[39556] <= 16'b0000_0000_0000_0000;
array[39557] <= 16'b0000_0000_0000_0000;
array[39558] <= 16'b0000_0000_0000_0000;
array[39559] <= 16'b0000_0000_0000_0000;
array[39560] <= 16'b0000_0000_0000_0000;
array[39561] <= 16'b0000_0000_0000_0000;
array[39562] <= 16'b0000_0000_0000_0000;
array[39563] <= 16'b0000_0000_0000_0000;
array[39564] <= 16'b0000_0000_0000_0000;
array[39565] <= 16'b0000_0000_0000_0000;
array[39566] <= 16'b0000_0000_0000_0000;
array[39567] <= 16'b0000_0000_0000_0000;
array[39568] <= 16'b0000_0000_0000_0000;
array[39569] <= 16'b0000_0000_0000_0000;
array[39570] <= 16'b0000_0000_0000_0000;
array[39571] <= 16'b0000_0000_0000_0000;
array[39572] <= 16'b0000_0000_0000_0000;
array[39573] <= 16'b0000_0000_0000_0000;
array[39574] <= 16'b0000_0000_0000_0000;
array[39575] <= 16'b0000_0000_0000_0000;
array[39576] <= 16'b0000_0000_0000_0000;
array[39577] <= 16'b0000_0000_0000_0000;
array[39578] <= 16'b0000_0000_0000_0000;
array[39579] <= 16'b0000_0000_0000_0000;
array[39580] <= 16'b0000_0000_0000_0000;
array[39581] <= 16'b0000_0000_0000_0000;
array[39582] <= 16'b0000_0000_0000_0000;
array[39583] <= 16'b0000_0000_0000_0000;
array[39584] <= 16'b0000_0000_0000_0000;
array[39585] <= 16'b0000_0000_0000_0000;
array[39586] <= 16'b0000_0000_0000_0000;
array[39587] <= 16'b0000_0000_0000_0000;
array[39588] <= 16'b0000_0000_0000_0000;
array[39589] <= 16'b0000_0000_0000_0000;
array[39590] <= 16'b0000_0000_0000_0000;
array[39591] <= 16'b0000_0000_0000_0000;
array[39592] <= 16'b0000_0000_0000_0000;
array[39593] <= 16'b0000_0000_0000_0000;
array[39594] <= 16'b0000_0000_0000_0000;
array[39595] <= 16'b0000_0000_0000_0000;
array[39596] <= 16'b0000_0000_0000_0000;
array[39597] <= 16'b0000_0000_0000_0000;
array[39598] <= 16'b0000_0000_0000_0000;
array[39599] <= 16'b0000_0000_0000_0000;
array[39600] <= 16'b0000_0000_0000_0000;
array[39601] <= 16'b0000_0000_0000_0000;
array[39602] <= 16'b0000_0000_0000_0000;
array[39603] <= 16'b0000_0000_0000_0000;
array[39604] <= 16'b0000_0000_0000_0000;
array[39605] <= 16'b0000_0000_0000_0000;
array[39606] <= 16'b0000_0000_0000_0000;
array[39607] <= 16'b0000_0000_0000_0000;
array[39608] <= 16'b0000_0000_0000_0000;
array[39609] <= 16'b0000_0000_0000_0000;
array[39610] <= 16'b0000_0000_0000_0000;
array[39611] <= 16'b0000_0000_0000_0000;
array[39612] <= 16'b0000_0000_0000_0000;
array[39613] <= 16'b0000_0000_0000_0000;
array[39614] <= 16'b0000_0000_0000_0000;
array[39615] <= 16'b0000_0000_0000_0000;
array[39616] <= 16'b0000_0000_0000_0000;
array[39617] <= 16'b0000_0000_0000_0000;
array[39618] <= 16'b0000_0000_0000_0000;
array[39619] <= 16'b0000_0000_0000_0000;
array[39620] <= 16'b0000_0000_0000_0000;
array[39621] <= 16'b0000_0000_0000_0000;
array[39622] <= 16'b0000_0000_0000_0000;
array[39623] <= 16'b0000_0000_0000_0000;
array[39624] <= 16'b0000_0000_0000_0000;
array[39625] <= 16'b0000_0000_0000_0000;
array[39626] <= 16'b0000_0000_0000_0000;
array[39627] <= 16'b0000_0000_0000_0000;
array[39628] <= 16'b0000_0000_0000_0000;
array[39629] <= 16'b0000_0000_0000_0000;
array[39630] <= 16'b0000_0000_0000_0000;
array[39631] <= 16'b0000_0000_0000_0000;
array[39632] <= 16'b0000_0000_0000_0000;
array[39633] <= 16'b0000_0000_0000_0000;
array[39634] <= 16'b0000_0000_0000_0000;
array[39635] <= 16'b0000_0000_0000_0000;
array[39636] <= 16'b0000_0000_0000_0000;
array[39637] <= 16'b0000_0000_0000_0000;
array[39638] <= 16'b0000_0000_0000_0000;
array[39639] <= 16'b0000_0000_0000_0000;
array[39640] <= 16'b0000_0000_0000_0000;
array[39641] <= 16'b0000_0000_0000_0000;
array[39642] <= 16'b0000_0000_0000_0000;
array[39643] <= 16'b0000_0000_0000_0000;
array[39644] <= 16'b0000_0000_0000_0000;
array[39645] <= 16'b0000_0000_0000_0000;
array[39646] <= 16'b0000_0000_0000_0000;
array[39647] <= 16'b0000_0000_0000_0000;
array[39648] <= 16'b0000_0000_0000_0000;
array[39649] <= 16'b0000_0000_0000_0000;
array[39650] <= 16'b0000_0000_0000_0000;
array[39651] <= 16'b0000_0000_0000_0000;
array[39652] <= 16'b0000_0000_0000_0000;
array[39653] <= 16'b0000_0000_0000_0000;
array[39654] <= 16'b0000_0000_0000_0000;
array[39655] <= 16'b0000_0000_0000_0000;
array[39656] <= 16'b0000_0000_0000_0000;
array[39657] <= 16'b0000_0000_0000_0000;
array[39658] <= 16'b0000_0000_0000_0000;
array[39659] <= 16'b0000_0000_0000_0000;
array[39660] <= 16'b0000_0000_0000_0000;
array[39661] <= 16'b0000_0000_0000_0000;
array[39662] <= 16'b0000_0000_0000_0000;
array[39663] <= 16'b0000_0000_0000_0000;
array[39664] <= 16'b0000_0000_0000_0000;
array[39665] <= 16'b0000_0000_0000_0000;
array[39666] <= 16'b0000_0000_0000_0000;
array[39667] <= 16'b0000_0000_0000_0000;
array[39668] <= 16'b0000_0000_0000_0000;
array[39669] <= 16'b0000_0000_0000_0000;
array[39670] <= 16'b0000_0000_0000_0000;
array[39671] <= 16'b0000_0000_0000_0000;
array[39672] <= 16'b0000_0000_0000_0000;
array[39673] <= 16'b0000_0000_0000_0000;
array[39674] <= 16'b0000_0000_0000_0000;
array[39675] <= 16'b0000_0000_0000_0000;
array[39676] <= 16'b0000_0000_0000_0000;
array[39677] <= 16'b0000_0000_0000_0000;
array[39678] <= 16'b0000_0000_0000_0000;
array[39679] <= 16'b0000_0000_0000_0000;
array[39680] <= 16'b0000_0000_0000_0000;
array[39681] <= 16'b0000_0000_0000_0000;
array[39682] <= 16'b0000_0000_0000_0000;
array[39683] <= 16'b0000_0000_0000_0000;
array[39684] <= 16'b0000_0000_0000_0000;
array[39685] <= 16'b0000_0000_0000_0000;
array[39686] <= 16'b0000_0000_0000_0000;
array[39687] <= 16'b0000_0000_0000_0000;
array[39688] <= 16'b0000_0000_0000_0000;
array[39689] <= 16'b0000_0000_0000_0000;
array[39690] <= 16'b0000_0000_0000_0000;
array[39691] <= 16'b0000_0000_0000_0000;
array[39692] <= 16'b0000_0000_0000_0000;
array[39693] <= 16'b0000_0000_0000_0000;
array[39694] <= 16'b0000_0000_0000_0000;
array[39695] <= 16'b0000_0000_0000_0000;
array[39696] <= 16'b0000_0000_0000_0000;
array[39697] <= 16'b0000_0000_0000_0000;
array[39698] <= 16'b0000_0000_0000_0000;
array[39699] <= 16'b0000_0000_0000_0000;
array[39700] <= 16'b0000_0000_0000_0000;
array[39701] <= 16'b0000_0000_0000_0000;
array[39702] <= 16'b0000_0000_0000_0000;
array[39703] <= 16'b0000_0000_0000_0000;
array[39704] <= 16'b0000_0000_0000_0000;
array[39705] <= 16'b0000_0000_0000_0000;
array[39706] <= 16'b0000_0000_0000_0000;
array[39707] <= 16'b0000_0000_0000_0000;
array[39708] <= 16'b0000_0000_0000_0000;
array[39709] <= 16'b0000_0000_0000_0000;
array[39710] <= 16'b0000_0000_0000_0000;
array[39711] <= 16'b0000_0000_0000_0000;
array[39712] <= 16'b0000_0000_0000_0000;
array[39713] <= 16'b0000_0000_0000_0000;
array[39714] <= 16'b0000_0000_0000_0000;
array[39715] <= 16'b0000_0000_0000_0000;
array[39716] <= 16'b0000_0000_0000_0000;
array[39717] <= 16'b0000_0000_0000_0000;
array[39718] <= 16'b0000_0000_0000_0000;
array[39719] <= 16'b0000_0000_0000_0000;
array[39720] <= 16'b0000_0000_0000_0000;
array[39721] <= 16'b0000_0000_0000_0000;
array[39722] <= 16'b0000_0000_0000_0000;
array[39723] <= 16'b0000_0000_0000_0000;
array[39724] <= 16'b0000_0000_0000_0000;
array[39725] <= 16'b0000_0000_0000_0000;
array[39726] <= 16'b0000_0000_0000_0000;
array[39727] <= 16'b0000_0000_0000_0000;
array[39728] <= 16'b0000_0000_0000_0000;
array[39729] <= 16'b0000_0000_0000_0000;
array[39730] <= 16'b0000_0000_0000_0000;
array[39731] <= 16'b0000_0000_0000_0000;
array[39732] <= 16'b0000_0000_0000_0000;
array[39733] <= 16'b0000_0000_0000_0000;
array[39734] <= 16'b0000_0000_0000_0000;
array[39735] <= 16'b0000_0000_0000_0000;
array[39736] <= 16'b0000_0000_0000_0000;
array[39737] <= 16'b0000_0000_0000_0000;
array[39738] <= 16'b0000_0000_0000_0000;
array[39739] <= 16'b0000_0000_0000_0000;
array[39740] <= 16'b0000_0000_0000_0000;
array[39741] <= 16'b0000_0000_0000_0000;
array[39742] <= 16'b0000_0000_0000_0000;
array[39743] <= 16'b0000_0000_0000_0000;
array[39744] <= 16'b0000_0000_0000_0000;
array[39745] <= 16'b0000_0000_0000_0000;
array[39746] <= 16'b0000_0000_0000_0000;
array[39747] <= 16'b0000_0000_0000_0000;
array[39748] <= 16'b0000_0000_0000_0000;
array[39749] <= 16'b0000_0000_0000_0000;
array[39750] <= 16'b0000_0000_0000_0000;
array[39751] <= 16'b0000_0000_0000_0000;
array[39752] <= 16'b0000_0000_0000_0000;
array[39753] <= 16'b0000_0000_0000_0000;
array[39754] <= 16'b0000_0000_0000_0000;
array[39755] <= 16'b0000_0000_0000_0000;
array[39756] <= 16'b0000_0000_0000_0000;
array[39757] <= 16'b0000_0000_0000_0000;
array[39758] <= 16'b0000_0000_0000_0000;
array[39759] <= 16'b0000_0000_0000_0000;
array[39760] <= 16'b0000_0000_0000_0000;
array[39761] <= 16'b0000_0000_0000_0000;
array[39762] <= 16'b0000_0000_0000_0000;
array[39763] <= 16'b0000_0000_0000_0000;
array[39764] <= 16'b0000_0000_0000_0000;
array[39765] <= 16'b0000_0000_0000_0000;
array[39766] <= 16'b0000_0000_0000_0000;
array[39767] <= 16'b0000_0000_0000_0000;
array[39768] <= 16'b0000_0000_0000_0000;
array[39769] <= 16'b0000_0000_0000_0000;
array[39770] <= 16'b0000_0000_0000_0000;
array[39771] <= 16'b0000_0000_0000_0000;
array[39772] <= 16'b0000_0000_0000_0000;
array[39773] <= 16'b0000_0000_0000_0000;
array[39774] <= 16'b0000_0000_0000_0000;
array[39775] <= 16'b0000_0000_0000_0000;
array[39776] <= 16'b0000_0000_0000_0000;
array[39777] <= 16'b0000_0000_0000_0000;
array[39778] <= 16'b0000_0000_0000_0000;
array[39779] <= 16'b0000_0000_0000_0000;
array[39780] <= 16'b0000_0000_0000_0000;
array[39781] <= 16'b0000_0000_0000_0000;
array[39782] <= 16'b0000_0000_0000_0000;
array[39783] <= 16'b0000_0000_0000_0000;
array[39784] <= 16'b0000_0000_0000_0000;
array[39785] <= 16'b0000_0000_0000_0000;
array[39786] <= 16'b0000_0000_0000_0000;
array[39787] <= 16'b0000_0000_0000_0000;
array[39788] <= 16'b0000_0000_0000_0000;
array[39789] <= 16'b0000_0000_0000_0000;
array[39790] <= 16'b0000_0000_0000_0000;
array[39791] <= 16'b0000_0000_0000_0000;
array[39792] <= 16'b0000_0000_0000_0000;
array[39793] <= 16'b0000_0000_0000_0000;
array[39794] <= 16'b0000_0000_0000_0000;
array[39795] <= 16'b0000_0000_0000_0000;
array[39796] <= 16'b0000_0000_0000_0000;
array[39797] <= 16'b0000_0000_0000_0000;
array[39798] <= 16'b0000_0000_0000_0000;
array[39799] <= 16'b0000_0000_0000_0000;
array[39800] <= 16'b0000_0000_0000_0000;
array[39801] <= 16'b0000_0000_0000_0000;
array[39802] <= 16'b0000_0000_0000_0000;
array[39803] <= 16'b0000_0000_0000_0000;
array[39804] <= 16'b0000_0000_0000_0000;
array[39805] <= 16'b0000_0000_0000_0000;
array[39806] <= 16'b0000_0000_0000_0000;
array[39807] <= 16'b0000_0000_0000_0000;
array[39808] <= 16'b0000_0000_0000_0000;
array[39809] <= 16'b0000_0000_0000_0000;
array[39810] <= 16'b0000_0000_0000_0000;
array[39811] <= 16'b0000_0000_0000_0000;
array[39812] <= 16'b0000_0000_0000_0000;
array[39813] <= 16'b0000_0000_0000_0000;
array[39814] <= 16'b0000_0000_0000_0000;
array[39815] <= 16'b0000_0000_0000_0000;
array[39816] <= 16'b0000_0000_0000_0000;
array[39817] <= 16'b0000_0000_0000_0000;
array[39818] <= 16'b0000_0000_0000_0000;
array[39819] <= 16'b0000_0000_0000_0000;
array[39820] <= 16'b0000_0000_0000_0000;
array[39821] <= 16'b0000_0000_0000_0000;
array[39822] <= 16'b0000_0000_0000_0000;
array[39823] <= 16'b0000_0000_0000_0000;
array[39824] <= 16'b0000_0000_0000_0000;
array[39825] <= 16'b0000_0000_0000_0000;
array[39826] <= 16'b0000_0000_0000_0000;
array[39827] <= 16'b0000_0000_0000_0000;
array[39828] <= 16'b0000_0000_0000_0000;
array[39829] <= 16'b0000_0000_0000_0000;
array[39830] <= 16'b0000_0000_0000_0000;
array[39831] <= 16'b0000_0000_0000_0000;
array[39832] <= 16'b0000_0000_0000_0000;
array[39833] <= 16'b0000_0000_0000_0000;
array[39834] <= 16'b0000_0000_0000_0000;
array[39835] <= 16'b0000_0000_0000_0000;
array[39836] <= 16'b0000_0000_0000_0000;
array[39837] <= 16'b0000_0000_0000_0000;
array[39838] <= 16'b0000_0000_0000_0000;
array[39839] <= 16'b0000_0000_0000_0000;
array[39840] <= 16'b0000_0000_0000_0000;
array[39841] <= 16'b0000_0000_0000_0000;
array[39842] <= 16'b0000_0000_0000_0000;
array[39843] <= 16'b0000_0000_0000_0000;
array[39844] <= 16'b0000_0000_0000_0000;
array[39845] <= 16'b0000_0000_0000_0000;
array[39846] <= 16'b0000_0000_0000_0000;
array[39847] <= 16'b0000_0000_0000_0000;
array[39848] <= 16'b0000_0000_0000_0000;
array[39849] <= 16'b0000_0000_0000_0000;
array[39850] <= 16'b0000_0000_0000_0000;
array[39851] <= 16'b0000_0000_0000_0000;
array[39852] <= 16'b0000_0000_0000_0000;
array[39853] <= 16'b0000_0000_0000_0000;
array[39854] <= 16'b0000_0000_0000_0000;
array[39855] <= 16'b0000_0000_0000_0000;
array[39856] <= 16'b0000_0000_0000_0000;
array[39857] <= 16'b0000_0000_0000_0000;
array[39858] <= 16'b0000_0000_0000_0000;
array[39859] <= 16'b0000_0000_0000_0000;
array[39860] <= 16'b0000_0000_0000_0000;
array[39861] <= 16'b0000_0000_0000_0000;
array[39862] <= 16'b0000_0000_0000_0000;
array[39863] <= 16'b0000_0000_0000_0000;
array[39864] <= 16'b0000_0000_0000_0000;
array[39865] <= 16'b0000_0000_0000_0000;
array[39866] <= 16'b0000_0000_0000_0000;
array[39867] <= 16'b0000_0000_0000_0000;
array[39868] <= 16'b0000_0000_0000_0000;
array[39869] <= 16'b0000_0000_0000_0000;
array[39870] <= 16'b0000_0000_0000_0000;
array[39871] <= 16'b0000_0000_0000_0000;
array[39872] <= 16'b0000_0000_0000_0000;
array[39873] <= 16'b0000_0000_0000_0000;
array[39874] <= 16'b0000_0000_0000_0000;
array[39875] <= 16'b0000_0000_0000_0000;
array[39876] <= 16'b0000_0000_0000_0000;
array[39877] <= 16'b0000_0000_0000_0000;
array[39878] <= 16'b0000_0000_0000_0000;
array[39879] <= 16'b0000_0000_0000_0000;
array[39880] <= 16'b0000_0000_0000_0000;
array[39881] <= 16'b0000_0000_0000_0000;
array[39882] <= 16'b0000_0000_0000_0000;
array[39883] <= 16'b0000_0000_0000_0000;
array[39884] <= 16'b0000_0000_0000_0000;
array[39885] <= 16'b0000_0000_0000_0000;
array[39886] <= 16'b0000_0000_0000_0000;
array[39887] <= 16'b0000_0000_0000_0000;
array[39888] <= 16'b0000_0000_0000_0000;
array[39889] <= 16'b0000_0000_0000_0000;
array[39890] <= 16'b0000_0000_0000_0000;
array[39891] <= 16'b0000_0000_0000_0000;
array[39892] <= 16'b0000_0000_0000_0000;
array[39893] <= 16'b0000_0000_0000_0000;
array[39894] <= 16'b0000_0000_0000_0000;
array[39895] <= 16'b0000_0000_0000_0000;
array[39896] <= 16'b0000_0000_0000_0000;
array[39897] <= 16'b0000_0000_0000_0000;
array[39898] <= 16'b0000_0000_0000_0000;
array[39899] <= 16'b0000_0000_0000_0000;
array[39900] <= 16'b0000_0000_0000_0000;
array[39901] <= 16'b0000_0000_0000_0000;
array[39902] <= 16'b0000_0000_0000_0000;
array[39903] <= 16'b0000_0000_0000_0000;
array[39904] <= 16'b0000_0000_0000_0000;
array[39905] <= 16'b0000_0000_0000_0000;
array[39906] <= 16'b0000_0000_0000_0000;
array[39907] <= 16'b0000_0000_0000_0000;
array[39908] <= 16'b0000_0000_0000_0000;
array[39909] <= 16'b0000_0000_0000_0000;
array[39910] <= 16'b0000_0000_0000_0000;
array[39911] <= 16'b0000_0000_0000_0000;
array[39912] <= 16'b0000_0000_0000_0000;
array[39913] <= 16'b0000_0000_0000_0000;
array[39914] <= 16'b0000_0000_0000_0000;
array[39915] <= 16'b0000_0000_0000_0000;
array[39916] <= 16'b0000_0000_0000_0000;
array[39917] <= 16'b0000_0000_0000_0000;
array[39918] <= 16'b0000_0000_0000_0000;
array[39919] <= 16'b0000_0000_0000_0000;
array[39920] <= 16'b0000_0000_0000_0000;
array[39921] <= 16'b0000_0000_0000_0000;
array[39922] <= 16'b0000_0000_0000_0000;
array[39923] <= 16'b0000_0000_0000_0000;
array[39924] <= 16'b0000_0000_0000_0000;
array[39925] <= 16'b0000_0000_0000_0000;
array[39926] <= 16'b0000_0000_0000_0000;
array[39927] <= 16'b0000_0000_0000_0000;
array[39928] <= 16'b0000_0000_0000_0000;
array[39929] <= 16'b0000_0000_0000_0000;
array[39930] <= 16'b0000_0000_0000_0000;
array[39931] <= 16'b0000_0000_0000_0000;
array[39932] <= 16'b0000_0000_0000_0000;
array[39933] <= 16'b0000_0000_0000_0000;
array[39934] <= 16'b0000_0000_0000_0000;
array[39935] <= 16'b0000_0000_0000_0000;
array[39936] <= 16'b0000_0000_0000_0000;
array[39937] <= 16'b0000_0000_0000_0000;
array[39938] <= 16'b0000_0000_0000_0000;
array[39939] <= 16'b0000_0000_0000_0000;
array[39940] <= 16'b0000_0000_0000_0000;
array[39941] <= 16'b0000_0000_0000_0000;
array[39942] <= 16'b0000_0000_0000_0000;
array[39943] <= 16'b0000_0000_0000_0000;
array[39944] <= 16'b0000_0000_0000_0000;
array[39945] <= 16'b0000_0000_0000_0000;
array[39946] <= 16'b0000_0000_0000_0000;
array[39947] <= 16'b0000_0000_0000_0000;
array[39948] <= 16'b0000_0000_0000_0000;
array[39949] <= 16'b0000_0000_0000_0000;
array[39950] <= 16'b0000_0000_0000_0000;
array[39951] <= 16'b0000_0000_0000_0000;
array[39952] <= 16'b0000_0000_0000_0000;
array[39953] <= 16'b0000_0000_0000_0000;
array[39954] <= 16'b0000_0000_0000_0000;
array[39955] <= 16'b0000_0000_0000_0000;
array[39956] <= 16'b0000_0000_0000_0000;
array[39957] <= 16'b0000_0000_0000_0000;
array[39958] <= 16'b0000_0000_0000_0000;
array[39959] <= 16'b0000_0000_0000_0000;
array[39960] <= 16'b0000_0000_0000_0000;
array[39961] <= 16'b0000_0000_0000_0000;
array[39962] <= 16'b0000_0000_0000_0000;
array[39963] <= 16'b0000_0000_0000_0000;
array[39964] <= 16'b0000_0000_0000_0000;
array[39965] <= 16'b0000_0000_0000_0000;
array[39966] <= 16'b0000_0000_0000_0000;
array[39967] <= 16'b0000_0000_0000_0000;
array[39968] <= 16'b0000_0000_0000_0000;
array[39969] <= 16'b0000_0000_0000_0000;
array[39970] <= 16'b0000_0000_0000_0000;
array[39971] <= 16'b0000_0000_0000_0000;
array[39972] <= 16'b0000_0000_0000_0000;
array[39973] <= 16'b0000_0000_0000_0000;
array[39974] <= 16'b0000_0000_0000_0000;
array[39975] <= 16'b0000_0000_0000_0000;
array[39976] <= 16'b0000_0000_0000_0000;
array[39977] <= 16'b0000_0000_0000_0000;
array[39978] <= 16'b0000_0000_0000_0000;
array[39979] <= 16'b0000_0000_0000_0000;
array[39980] <= 16'b0000_0000_0000_0000;
array[39981] <= 16'b0000_0000_0000_0000;
array[39982] <= 16'b0000_0000_0000_0000;
array[39983] <= 16'b0000_0000_0000_0000;
array[39984] <= 16'b0000_0000_0000_0000;
array[39985] <= 16'b0000_0000_0000_0000;
array[39986] <= 16'b0000_0000_0000_0000;
array[39987] <= 16'b0000_0000_0000_0000;
array[39988] <= 16'b0000_0000_0000_0000;
array[39989] <= 16'b0000_0000_0000_0000;
array[39990] <= 16'b0000_0000_0000_0000;
array[39991] <= 16'b0000_0000_0000_0000;
array[39992] <= 16'b0000_0000_0000_0000;
array[39993] <= 16'b0000_0000_0000_0000;
array[39994] <= 16'b0000_0000_0000_0000;
array[39995] <= 16'b0000_0000_0000_0000;
array[39996] <= 16'b0000_0000_0000_0000;
array[39997] <= 16'b0000_0000_0000_0000;
array[39998] <= 16'b0000_0000_0000_0000;
array[39999] <= 16'b0000_0000_0000_0000;
array[40000] <= 16'b0000_0000_0000_0000;
array[40001] <= 16'b0000_0000_0000_0000;
array[40002] <= 16'b0000_0000_0000_0000;
array[40003] <= 16'b0000_0000_0000_0000;
array[40004] <= 16'b0000_0000_0000_0000;
array[40005] <= 16'b0000_0000_0000_0000;
array[40006] <= 16'b0000_0000_0000_0000;
array[40007] <= 16'b0000_0000_0000_0000;
array[40008] <= 16'b0000_0000_0000_0000;
array[40009] <= 16'b0000_0000_0000_0000;
array[40010] <= 16'b0000_0000_0000_0000;
array[40011] <= 16'b0000_0000_0000_0000;
array[40012] <= 16'b0000_0000_0000_0000;
array[40013] <= 16'b0000_0000_0000_0000;
array[40014] <= 16'b0000_0000_0000_0000;
array[40015] <= 16'b0000_0000_0000_0000;
array[40016] <= 16'b0000_0000_0000_0000;
array[40017] <= 16'b0000_0000_0000_0000;
array[40018] <= 16'b0000_0000_0000_0000;
array[40019] <= 16'b0000_0000_0000_0000;
array[40020] <= 16'b0000_0000_0000_0000;
array[40021] <= 16'b0000_0000_0000_0000;
array[40022] <= 16'b0000_0000_0000_0000;
array[40023] <= 16'b0000_0000_0000_0000;
array[40024] <= 16'b0000_0000_0000_0000;
array[40025] <= 16'b0000_0000_0000_0000;
array[40026] <= 16'b0000_0000_0000_0000;
array[40027] <= 16'b0000_0000_0000_0000;
array[40028] <= 16'b0000_0000_0000_0000;
array[40029] <= 16'b0000_0000_0000_0000;
array[40030] <= 16'b0000_0000_0000_0000;
array[40031] <= 16'b0000_0000_0000_0000;
array[40032] <= 16'b0000_0000_0000_0000;
array[40033] <= 16'b0000_0000_0000_0000;
array[40034] <= 16'b0000_0000_0000_0000;
array[40035] <= 16'b0000_0000_0000_0000;
array[40036] <= 16'b0000_0000_0000_0000;
array[40037] <= 16'b0000_0000_0000_0000;
array[40038] <= 16'b0000_0000_0000_0000;
array[40039] <= 16'b0000_0000_0000_0000;
array[40040] <= 16'b0000_0000_0000_0000;
array[40041] <= 16'b0000_0000_0000_0000;
array[40042] <= 16'b0000_0000_0000_0000;
array[40043] <= 16'b0000_0000_0000_0000;
array[40044] <= 16'b0000_0000_0000_0000;
array[40045] <= 16'b0000_0000_0000_0000;
array[40046] <= 16'b0000_0000_0000_0000;
array[40047] <= 16'b0000_0000_0000_0000;
array[40048] <= 16'b0000_0000_0000_0000;
array[40049] <= 16'b0000_0000_0000_0000;
array[40050] <= 16'b0000_0000_0000_0000;
array[40051] <= 16'b0000_0000_0000_0000;
array[40052] <= 16'b0000_0000_0000_0000;
array[40053] <= 16'b0000_0000_0000_0000;
array[40054] <= 16'b0000_0000_0000_0000;
array[40055] <= 16'b0000_0000_0000_0000;
array[40056] <= 16'b0000_0000_0000_0000;
array[40057] <= 16'b0000_0000_0000_0000;
array[40058] <= 16'b0000_0000_0000_0000;
array[40059] <= 16'b0000_0000_0000_0000;
array[40060] <= 16'b0000_0000_0000_0000;
array[40061] <= 16'b0000_0000_0000_0000;
array[40062] <= 16'b0000_0000_0000_0000;
array[40063] <= 16'b0000_0000_0000_0000;
array[40064] <= 16'b0000_0000_0000_0000;
array[40065] <= 16'b0000_0000_0000_0000;
array[40066] <= 16'b0000_0000_0000_0000;
array[40067] <= 16'b0000_0000_0000_0000;
array[40068] <= 16'b0000_0000_0000_0000;
array[40069] <= 16'b0000_0000_0000_0000;
array[40070] <= 16'b0000_0000_0000_0000;
array[40071] <= 16'b0000_0000_0000_0000;
array[40072] <= 16'b0000_0000_0000_0000;
array[40073] <= 16'b0000_0000_0000_0000;
array[40074] <= 16'b0000_0000_0000_0000;
array[40075] <= 16'b0000_0000_0000_0000;
array[40076] <= 16'b0000_0000_0000_0000;
array[40077] <= 16'b0000_0000_0000_0000;
array[40078] <= 16'b0000_0000_0000_0000;
array[40079] <= 16'b0000_0000_0000_0000;
array[40080] <= 16'b0000_0000_0000_0000;
array[40081] <= 16'b0000_0000_0000_0000;
array[40082] <= 16'b0000_0000_0000_0000;
array[40083] <= 16'b0000_0000_0000_0000;
array[40084] <= 16'b0000_0000_0000_0000;
array[40085] <= 16'b0000_0000_0000_0000;
array[40086] <= 16'b0000_0000_0000_0000;
array[40087] <= 16'b0000_0000_0000_0000;
array[40088] <= 16'b0000_0000_0000_0000;
array[40089] <= 16'b0000_0000_0000_0000;
array[40090] <= 16'b0000_0000_0000_0000;
array[40091] <= 16'b0000_0000_0000_0000;
array[40092] <= 16'b0000_0000_0000_0000;
array[40093] <= 16'b0000_0000_0000_0000;
array[40094] <= 16'b0000_0000_0000_0000;
array[40095] <= 16'b0000_0000_0000_0000;
array[40096] <= 16'b0000_0000_0000_0000;
array[40097] <= 16'b0000_0000_0000_0000;
array[40098] <= 16'b0000_0000_0000_0000;
array[40099] <= 16'b0000_0000_0000_0000;
array[40100] <= 16'b0000_0000_0000_0000;
array[40101] <= 16'b0000_0000_0000_0000;
array[40102] <= 16'b0000_0000_0000_0000;
array[40103] <= 16'b0000_0000_0000_0000;
array[40104] <= 16'b0000_0000_0000_0000;
array[40105] <= 16'b0000_0000_0000_0000;
array[40106] <= 16'b0000_0000_0000_0000;
array[40107] <= 16'b0000_0000_0000_0000;
array[40108] <= 16'b0000_0000_0000_0000;
array[40109] <= 16'b0000_0000_0000_0000;
array[40110] <= 16'b0000_0000_0000_0000;
array[40111] <= 16'b0000_0000_0000_0000;
array[40112] <= 16'b0000_0000_0000_0000;
array[40113] <= 16'b0000_0000_0000_0000;
array[40114] <= 16'b0000_0000_0000_0000;
array[40115] <= 16'b0000_0000_0000_0000;
array[40116] <= 16'b0000_0000_0000_0000;
array[40117] <= 16'b0000_0000_0000_0000;
array[40118] <= 16'b0000_0000_0000_0000;
array[40119] <= 16'b0000_0000_0000_0000;
array[40120] <= 16'b0000_0000_0000_0000;
array[40121] <= 16'b0000_0000_0000_0000;
array[40122] <= 16'b0000_0000_0000_0000;
array[40123] <= 16'b0000_0000_0000_0000;
array[40124] <= 16'b0000_0000_0000_0000;
array[40125] <= 16'b0000_0000_0000_0000;
array[40126] <= 16'b0000_0000_0000_0000;
array[40127] <= 16'b0000_0000_0000_0000;
array[40128] <= 16'b0000_0000_0000_0000;
array[40129] <= 16'b0000_0000_0000_0000;
array[40130] <= 16'b0000_0000_0000_0000;
array[40131] <= 16'b0000_0000_0000_0000;
array[40132] <= 16'b0000_0000_0000_0000;
array[40133] <= 16'b0000_0000_0000_0000;
array[40134] <= 16'b0000_0000_0000_0000;
array[40135] <= 16'b0000_0000_0000_0000;
array[40136] <= 16'b0000_0000_0000_0000;
array[40137] <= 16'b0000_0000_0000_0000;
array[40138] <= 16'b0000_0000_0000_0000;
array[40139] <= 16'b0000_0000_0000_0000;
array[40140] <= 16'b0000_0000_0000_0000;
array[40141] <= 16'b0000_0000_0000_0000;
array[40142] <= 16'b0000_0000_0000_0000;
array[40143] <= 16'b0000_0000_0000_0000;
array[40144] <= 16'b0000_0000_0000_0000;
array[40145] <= 16'b0000_0000_0000_0000;
array[40146] <= 16'b0000_0000_0000_0000;
array[40147] <= 16'b0000_0000_0000_0000;
array[40148] <= 16'b0000_0000_0000_0000;
array[40149] <= 16'b0000_0000_0000_0000;
array[40150] <= 16'b0000_0000_0000_0000;
array[40151] <= 16'b0000_0000_0000_0000;
array[40152] <= 16'b0000_0000_0000_0000;
array[40153] <= 16'b0000_0000_0000_0000;
array[40154] <= 16'b0000_0000_0000_0000;
array[40155] <= 16'b0000_0000_0000_0000;
array[40156] <= 16'b0000_0000_0000_0000;
array[40157] <= 16'b0000_0000_0000_0000;
array[40158] <= 16'b0000_0000_0000_0000;
array[40159] <= 16'b0000_0000_0000_0000;
array[40160] <= 16'b0000_0000_0000_0000;
array[40161] <= 16'b0000_0000_0000_0000;
array[40162] <= 16'b0000_0000_0000_0000;
array[40163] <= 16'b0000_0000_0000_0000;
array[40164] <= 16'b0000_0000_0000_0000;
array[40165] <= 16'b0000_0000_0000_0000;
array[40166] <= 16'b0000_0000_0000_0000;
array[40167] <= 16'b0000_0000_0000_0000;
array[40168] <= 16'b0000_0000_0000_0000;
array[40169] <= 16'b0000_0000_0000_0000;
array[40170] <= 16'b0000_0000_0000_0000;
array[40171] <= 16'b0000_0000_0000_0000;
array[40172] <= 16'b0000_0000_0000_0000;
array[40173] <= 16'b0000_0000_0000_0000;
array[40174] <= 16'b0000_0000_0000_0000;
array[40175] <= 16'b0000_0000_0000_0000;
array[40176] <= 16'b0000_0000_0000_0000;
array[40177] <= 16'b0000_0000_0000_0000;
array[40178] <= 16'b0000_0000_0000_0000;
array[40179] <= 16'b0000_0000_0000_0000;
array[40180] <= 16'b0000_0000_0000_0000;
array[40181] <= 16'b0000_0000_0000_0000;
array[40182] <= 16'b0000_0000_0000_0000;
array[40183] <= 16'b0000_0000_0000_0000;
array[40184] <= 16'b0000_0000_0000_0000;
array[40185] <= 16'b0000_0000_0000_0000;
array[40186] <= 16'b0000_0000_0000_0000;
array[40187] <= 16'b0000_0000_0000_0000;
array[40188] <= 16'b0000_0000_0000_0000;
array[40189] <= 16'b0000_0000_0000_0000;
array[40190] <= 16'b0000_0000_0000_0000;
array[40191] <= 16'b0000_0000_0000_0000;
array[40192] <= 16'b0000_0000_0000_0000;
array[40193] <= 16'b0000_0000_0000_0000;
array[40194] <= 16'b0000_0000_0000_0000;
array[40195] <= 16'b0000_0000_0000_0000;
array[40196] <= 16'b0000_0000_0000_0000;
array[40197] <= 16'b0000_0000_0000_0000;
array[40198] <= 16'b0000_0000_0000_0000;
array[40199] <= 16'b0000_0000_0000_0000;
array[40200] <= 16'b0000_0000_0000_0000;
array[40201] <= 16'b0000_0000_0000_0000;
array[40202] <= 16'b0000_0000_0000_0000;
array[40203] <= 16'b0000_0000_0000_0000;
array[40204] <= 16'b0000_0000_0000_0000;
array[40205] <= 16'b0000_0000_0000_0000;
array[40206] <= 16'b0000_0000_0000_0000;
array[40207] <= 16'b0000_0000_0000_0000;
array[40208] <= 16'b0000_0000_0000_0000;
array[40209] <= 16'b0000_0000_0000_0000;
array[40210] <= 16'b0000_0000_0000_0000;
array[40211] <= 16'b0000_0000_0000_0000;
array[40212] <= 16'b0000_0000_0000_0000;
array[40213] <= 16'b0000_0000_0000_0000;
array[40214] <= 16'b0000_0000_0000_0000;
array[40215] <= 16'b0000_0000_0000_0000;
array[40216] <= 16'b0000_0000_0000_0000;
array[40217] <= 16'b0000_0000_0000_0000;
array[40218] <= 16'b0000_0000_0000_0000;
array[40219] <= 16'b0000_0000_0000_0000;
array[40220] <= 16'b0000_0000_0000_0000;
array[40221] <= 16'b0000_0000_0000_0000;
array[40222] <= 16'b0000_0000_0000_0000;
array[40223] <= 16'b0000_0000_0000_0000;
array[40224] <= 16'b0000_0000_0000_0000;
array[40225] <= 16'b0000_0000_0000_0000;
array[40226] <= 16'b0000_0000_0000_0000;
array[40227] <= 16'b0000_0000_0000_0000;
array[40228] <= 16'b0000_0000_0000_0000;
array[40229] <= 16'b0000_0000_0000_0000;
array[40230] <= 16'b0000_0000_0000_0000;
array[40231] <= 16'b0000_0000_0000_0000;
array[40232] <= 16'b0000_0000_0000_0000;
array[40233] <= 16'b0000_0000_0000_0000;
array[40234] <= 16'b0000_0000_0000_0000;
array[40235] <= 16'b0000_0000_0000_0000;
array[40236] <= 16'b0000_0000_0000_0000;
array[40237] <= 16'b0000_0000_0000_0000;
array[40238] <= 16'b0000_0000_0000_0000;
array[40239] <= 16'b0000_0000_0000_0000;
array[40240] <= 16'b0000_0000_0000_0000;
array[40241] <= 16'b0000_0000_0000_0000;
array[40242] <= 16'b0000_0000_0000_0000;
array[40243] <= 16'b0000_0000_0000_0000;
array[40244] <= 16'b0000_0000_0000_0000;
array[40245] <= 16'b0000_0000_0000_0000;
array[40246] <= 16'b0000_0000_0000_0000;
array[40247] <= 16'b0000_0000_0000_0000;
array[40248] <= 16'b0000_0000_0000_0000;
array[40249] <= 16'b0000_0000_0000_0000;
array[40250] <= 16'b0000_0000_0000_0000;
array[40251] <= 16'b0000_0000_0000_0000;
array[40252] <= 16'b0000_0000_0000_0000;
array[40253] <= 16'b0000_0000_0000_0000;
array[40254] <= 16'b0000_0000_0000_0000;
array[40255] <= 16'b0000_0000_0000_0000;
array[40256] <= 16'b0000_0000_0000_0000;
array[40257] <= 16'b0000_0000_0000_0000;
array[40258] <= 16'b0000_0000_0000_0000;
array[40259] <= 16'b0000_0000_0000_0000;
array[40260] <= 16'b0000_0000_0000_0000;
array[40261] <= 16'b0000_0000_0000_0000;
array[40262] <= 16'b0000_0000_0000_0000;
array[40263] <= 16'b0000_0000_0000_0000;
array[40264] <= 16'b0000_0000_0000_0000;
array[40265] <= 16'b0000_0000_0000_0000;
array[40266] <= 16'b0000_0000_0000_0000;
array[40267] <= 16'b0000_0000_0000_0000;
array[40268] <= 16'b0000_0000_0000_0000;
array[40269] <= 16'b0000_0000_0000_0000;
array[40270] <= 16'b0000_0000_0000_0000;
array[40271] <= 16'b0000_0000_0000_0000;
array[40272] <= 16'b0000_0000_0000_0000;
array[40273] <= 16'b0000_0000_0000_0000;
array[40274] <= 16'b0000_0000_0000_0000;
array[40275] <= 16'b0000_0000_0000_0000;
array[40276] <= 16'b0000_0000_0000_0000;
array[40277] <= 16'b0000_0000_0000_0000;
array[40278] <= 16'b0000_0000_0000_0000;
array[40279] <= 16'b0000_0000_0000_0000;
array[40280] <= 16'b0000_0000_0000_0000;
array[40281] <= 16'b0000_0000_0000_0000;
array[40282] <= 16'b0000_0000_0000_0000;
array[40283] <= 16'b0000_0000_0000_0000;
array[40284] <= 16'b0000_0000_0000_0000;
array[40285] <= 16'b0000_0000_0000_0000;
array[40286] <= 16'b0000_0000_0000_0000;
array[40287] <= 16'b0000_0000_0000_0000;
array[40288] <= 16'b0000_0000_0000_0000;
array[40289] <= 16'b0000_0000_0000_0000;
array[40290] <= 16'b0000_0000_0000_0000;
array[40291] <= 16'b0000_0000_0000_0000;
array[40292] <= 16'b0000_0000_0000_0000;
array[40293] <= 16'b0000_0000_0000_0000;
array[40294] <= 16'b0000_0000_0000_0000;
array[40295] <= 16'b0000_0000_0000_0000;
array[40296] <= 16'b0000_0000_0000_0000;
array[40297] <= 16'b0000_0000_0000_0000;
array[40298] <= 16'b0000_0000_0000_0000;
array[40299] <= 16'b0000_0000_0000_0000;
array[40300] <= 16'b0000_0000_0000_0000;
array[40301] <= 16'b0000_0000_0000_0000;
array[40302] <= 16'b0000_0000_0000_0000;
array[40303] <= 16'b0000_0000_0000_0000;
array[40304] <= 16'b0000_0000_0000_0000;
array[40305] <= 16'b0000_0000_0000_0000;
array[40306] <= 16'b0000_0000_0000_0000;
array[40307] <= 16'b0000_0000_0000_0000;
array[40308] <= 16'b0000_0000_0000_0000;
array[40309] <= 16'b0000_0000_0000_0000;
array[40310] <= 16'b0000_0000_0000_0000;
array[40311] <= 16'b0000_0000_0000_0000;
array[40312] <= 16'b0000_0000_0000_0000;
array[40313] <= 16'b0000_0000_0000_0000;
array[40314] <= 16'b0000_0000_0000_0000;
array[40315] <= 16'b0000_0000_0000_0000;
array[40316] <= 16'b0000_0000_0000_0000;
array[40317] <= 16'b0000_0000_0000_0000;
array[40318] <= 16'b0000_0000_0000_0000;
array[40319] <= 16'b0000_0000_0000_0000;
array[40320] <= 16'b0000_0000_0000_0000;
array[40321] <= 16'b0000_0000_0000_0000;
array[40322] <= 16'b0000_0000_0000_0000;
array[40323] <= 16'b0000_0000_0000_0000;
array[40324] <= 16'b0000_0000_0000_0000;
array[40325] <= 16'b0000_0000_0000_0000;
array[40326] <= 16'b0000_0000_0000_0000;
array[40327] <= 16'b0000_0000_0000_0000;
array[40328] <= 16'b0000_0000_0000_0000;
array[40329] <= 16'b0000_0000_0000_0000;
array[40330] <= 16'b0000_0000_0000_0000;
array[40331] <= 16'b0000_0000_0000_0000;
array[40332] <= 16'b0000_0000_0000_0000;
array[40333] <= 16'b0000_0000_0000_0000;
array[40334] <= 16'b0000_0000_0000_0000;
array[40335] <= 16'b0000_0000_0000_0000;
array[40336] <= 16'b0000_0000_0000_0000;
array[40337] <= 16'b0000_0000_0000_0000;
array[40338] <= 16'b0000_0000_0000_0000;
array[40339] <= 16'b0000_0000_0000_0000;
array[40340] <= 16'b0000_0000_0000_0000;
array[40341] <= 16'b0000_0000_0000_0000;
array[40342] <= 16'b0000_0000_0000_0000;
array[40343] <= 16'b0000_0000_0000_0000;
array[40344] <= 16'b0000_0000_0000_0000;
array[40345] <= 16'b0000_0000_0000_0000;
array[40346] <= 16'b0000_0000_0000_0000;
array[40347] <= 16'b0000_0000_0000_0000;
array[40348] <= 16'b0000_0000_0000_0000;
array[40349] <= 16'b0000_0000_0000_0000;
array[40350] <= 16'b0000_0000_0000_0000;
array[40351] <= 16'b0000_0000_0000_0000;
array[40352] <= 16'b0000_0000_0000_0000;
array[40353] <= 16'b0000_0000_0000_0000;
array[40354] <= 16'b0000_0000_0000_0000;
array[40355] <= 16'b0000_0000_0000_0000;
array[40356] <= 16'b0000_0000_0000_0000;
array[40357] <= 16'b0000_0000_0000_0000;
array[40358] <= 16'b0000_0000_0000_0000;
array[40359] <= 16'b0000_0000_0000_0000;
array[40360] <= 16'b0000_0000_0000_0000;
array[40361] <= 16'b0000_0000_0000_0000;
array[40362] <= 16'b0000_0000_0000_0000;
array[40363] <= 16'b0000_0000_0000_0000;
array[40364] <= 16'b0000_0000_0000_0000;
array[40365] <= 16'b0000_0000_0000_0000;
array[40366] <= 16'b0000_0000_0000_0000;
array[40367] <= 16'b0000_0000_0000_0000;
array[40368] <= 16'b0000_0000_0000_0000;
array[40369] <= 16'b0000_0000_0000_0000;
array[40370] <= 16'b0000_0000_0000_0000;
array[40371] <= 16'b0000_0000_0000_0000;
array[40372] <= 16'b0000_0000_0000_0000;
array[40373] <= 16'b0000_0000_0000_0000;
array[40374] <= 16'b0000_0000_0000_0000;
array[40375] <= 16'b0000_0000_0000_0000;
array[40376] <= 16'b0000_0000_0000_0000;
array[40377] <= 16'b0000_0000_0000_0000;
array[40378] <= 16'b0000_0000_0000_0000;
array[40379] <= 16'b0000_0000_0000_0000;
array[40380] <= 16'b0000_0000_0000_0000;
array[40381] <= 16'b0000_0000_0000_0000;
array[40382] <= 16'b0000_0000_0000_0000;
array[40383] <= 16'b0000_0000_0000_0000;
array[40384] <= 16'b0000_0000_0000_0000;
array[40385] <= 16'b0000_0000_0000_0000;
array[40386] <= 16'b0000_0000_0000_0000;
array[40387] <= 16'b0000_0000_0000_0000;
array[40388] <= 16'b0000_0000_0000_0000;
array[40389] <= 16'b0000_0000_0000_0000;
array[40390] <= 16'b0000_0000_0000_0000;
array[40391] <= 16'b0000_0000_0000_0000;
array[40392] <= 16'b0000_0000_0000_0000;
array[40393] <= 16'b0000_0000_0000_0000;
array[40394] <= 16'b0000_0000_0000_0000;
array[40395] <= 16'b0000_0000_0000_0000;
array[40396] <= 16'b0000_0000_0000_0000;
array[40397] <= 16'b0000_0000_0000_0000;
array[40398] <= 16'b0000_0000_0000_0000;
array[40399] <= 16'b0000_0000_0000_0000;
array[40400] <= 16'b0000_0000_0000_0000;
array[40401] <= 16'b0000_0000_0000_0000;
array[40402] <= 16'b0000_0000_0000_0000;
array[40403] <= 16'b0000_0000_0000_0000;
array[40404] <= 16'b0000_0000_0000_0000;
array[40405] <= 16'b0000_0000_0000_0000;
array[40406] <= 16'b0000_0000_0000_0000;
array[40407] <= 16'b0000_0000_0000_0000;
array[40408] <= 16'b0000_0000_0000_0000;
array[40409] <= 16'b0000_0000_0000_0000;
array[40410] <= 16'b0000_0000_0000_0000;
array[40411] <= 16'b0000_0000_0000_0000;
array[40412] <= 16'b0000_0000_0000_0000;
array[40413] <= 16'b0000_0000_0000_0000;
array[40414] <= 16'b0000_0000_0000_0000;
array[40415] <= 16'b0000_0000_0000_0000;
array[40416] <= 16'b0000_0000_0000_0000;
array[40417] <= 16'b0000_0000_0000_0000;
array[40418] <= 16'b0000_0000_0000_0000;
array[40419] <= 16'b0000_0000_0000_0000;
array[40420] <= 16'b0000_0000_0000_0000;
array[40421] <= 16'b0000_0000_0000_0000;
array[40422] <= 16'b0000_0000_0000_0000;
array[40423] <= 16'b0000_0000_0000_0000;
array[40424] <= 16'b0000_0000_0000_0000;
array[40425] <= 16'b0000_0000_0000_0000;
array[40426] <= 16'b0000_0000_0000_0000;
array[40427] <= 16'b0000_0000_0000_0000;
array[40428] <= 16'b0000_0000_0000_0000;
array[40429] <= 16'b0000_0000_0000_0000;
array[40430] <= 16'b0000_0000_0000_0000;
array[40431] <= 16'b0000_0000_0000_0000;
array[40432] <= 16'b0000_0000_0000_0000;
array[40433] <= 16'b0000_0000_0000_0000;
array[40434] <= 16'b0000_0000_0000_0000;
array[40435] <= 16'b0000_0000_0000_0000;
array[40436] <= 16'b0000_0000_0000_0000;
array[40437] <= 16'b0000_0000_0000_0000;
array[40438] <= 16'b0000_0000_0000_0000;
array[40439] <= 16'b0000_0000_0000_0000;
array[40440] <= 16'b0000_0000_0000_0000;
array[40441] <= 16'b0000_0000_0000_0000;
array[40442] <= 16'b0000_0000_0000_0000;
array[40443] <= 16'b0000_0000_0000_0000;
array[40444] <= 16'b0000_0000_0000_0000;
array[40445] <= 16'b0000_0000_0000_0000;
array[40446] <= 16'b0000_0000_0000_0000;
array[40447] <= 16'b0000_0000_0000_0000;
array[40448] <= 16'b0000_0000_0000_0000;
array[40449] <= 16'b0000_0000_0000_0000;
array[40450] <= 16'b0000_0000_0000_0000;
array[40451] <= 16'b0000_0000_0000_0000;
array[40452] <= 16'b0000_0000_0000_0000;
array[40453] <= 16'b0000_0000_0000_0000;
array[40454] <= 16'b0000_0000_0000_0000;
array[40455] <= 16'b0000_0000_0000_0000;
array[40456] <= 16'b0000_0000_0000_0000;
array[40457] <= 16'b0000_0000_0000_0000;
array[40458] <= 16'b0000_0000_0000_0000;
array[40459] <= 16'b0000_0000_0000_0000;
array[40460] <= 16'b0000_0000_0000_0000;
array[40461] <= 16'b0000_0000_0000_0000;
array[40462] <= 16'b0000_0000_0000_0000;
array[40463] <= 16'b0000_0000_0000_0000;
array[40464] <= 16'b0000_0000_0000_0000;
array[40465] <= 16'b0000_0000_0000_0000;
array[40466] <= 16'b0000_0000_0000_0000;
array[40467] <= 16'b0000_0000_0000_0000;
array[40468] <= 16'b0000_0000_0000_0000;
array[40469] <= 16'b0000_0000_0000_0000;
array[40470] <= 16'b0000_0000_0000_0000;
array[40471] <= 16'b0000_0000_0000_0000;
array[40472] <= 16'b0000_0000_0000_0000;
array[40473] <= 16'b0000_0000_0000_0000;
array[40474] <= 16'b0000_0000_0000_0000;
array[40475] <= 16'b0000_0000_0000_0000;
array[40476] <= 16'b0000_0000_0000_0000;
array[40477] <= 16'b0000_0000_0000_0000;
array[40478] <= 16'b0000_0000_0000_0000;
array[40479] <= 16'b0000_0000_0000_0000;
array[40480] <= 16'b0000_0000_0000_0000;
array[40481] <= 16'b0000_0000_0000_0000;
array[40482] <= 16'b0000_0000_0000_0000;
array[40483] <= 16'b0000_0000_0000_0000;
array[40484] <= 16'b0000_0000_0000_0000;
array[40485] <= 16'b0000_0000_0000_0000;
array[40486] <= 16'b0000_0000_0000_0000;
array[40487] <= 16'b0000_0000_0000_0000;
array[40488] <= 16'b0000_0000_0000_0000;
array[40489] <= 16'b0000_0000_0000_0000;
array[40490] <= 16'b0000_0000_0000_0000;
array[40491] <= 16'b0000_0000_0000_0000;
array[40492] <= 16'b0000_0000_0000_0000;
array[40493] <= 16'b0000_0000_0000_0000;
array[40494] <= 16'b0000_0000_0000_0000;
array[40495] <= 16'b0000_0000_0000_0000;
array[40496] <= 16'b0000_0000_0000_0000;
array[40497] <= 16'b0000_0000_0000_0000;
array[40498] <= 16'b0000_0000_0000_0000;
array[40499] <= 16'b0000_0000_0000_0000;
array[40500] <= 16'b0000_0000_0000_0000;
array[40501] <= 16'b0000_0000_0000_0000;
array[40502] <= 16'b0000_0000_0000_0000;
array[40503] <= 16'b0000_0000_0000_0000;
array[40504] <= 16'b0000_0000_0000_0000;
array[40505] <= 16'b0000_0000_0000_0000;
array[40506] <= 16'b0000_0000_0000_0000;
array[40507] <= 16'b0000_0000_0000_0000;
array[40508] <= 16'b0000_0000_0000_0000;
array[40509] <= 16'b0000_0000_0000_0000;
array[40510] <= 16'b0000_0000_0000_0000;
array[40511] <= 16'b0000_0000_0000_0000;
array[40512] <= 16'b0000_0000_0000_0000;
array[40513] <= 16'b0000_0000_0000_0000;
array[40514] <= 16'b0000_0000_0000_0000;
array[40515] <= 16'b0000_0000_0000_0000;
array[40516] <= 16'b0000_0000_0000_0000;
array[40517] <= 16'b0000_0000_0000_0000;
array[40518] <= 16'b0000_0000_0000_0000;
array[40519] <= 16'b0000_0000_0000_0000;
array[40520] <= 16'b0000_0000_0000_0000;
array[40521] <= 16'b0000_0000_0000_0000;
array[40522] <= 16'b0000_0000_0000_0000;
array[40523] <= 16'b0000_0000_0000_0000;
array[40524] <= 16'b0000_0000_0000_0000;
array[40525] <= 16'b0000_0000_0000_0000;
array[40526] <= 16'b0000_0000_0000_0000;
array[40527] <= 16'b0000_0000_0000_0000;
array[40528] <= 16'b0000_0000_0000_0000;
array[40529] <= 16'b0000_0000_0000_0000;
array[40530] <= 16'b0000_0000_0000_0000;
array[40531] <= 16'b0000_0000_0000_0000;
array[40532] <= 16'b0000_0000_0000_0000;
array[40533] <= 16'b0000_0000_0000_0000;
array[40534] <= 16'b0000_0000_0000_0000;
array[40535] <= 16'b0000_0000_0000_0000;
array[40536] <= 16'b0000_0000_0000_0000;
array[40537] <= 16'b0000_0000_0000_0000;
array[40538] <= 16'b0000_0000_0000_0000;
array[40539] <= 16'b0000_0000_0000_0000;
array[40540] <= 16'b0000_0000_0000_0000;
array[40541] <= 16'b0000_0000_0000_0000;
array[40542] <= 16'b0000_0000_0000_0000;
array[40543] <= 16'b0000_0000_0000_0000;
array[40544] <= 16'b0000_0000_0000_0000;
array[40545] <= 16'b0000_0000_0000_0000;
array[40546] <= 16'b0000_0000_0000_0000;
array[40547] <= 16'b0000_0000_0000_0000;
array[40548] <= 16'b0000_0000_0000_0000;
array[40549] <= 16'b0000_0000_0000_0000;
array[40550] <= 16'b0000_0000_0000_0000;
array[40551] <= 16'b0000_0000_0000_0000;
array[40552] <= 16'b0000_0000_0000_0000;
array[40553] <= 16'b0000_0000_0000_0000;
array[40554] <= 16'b0000_0000_0000_0000;
array[40555] <= 16'b0000_0000_0000_0000;
array[40556] <= 16'b0000_0000_0000_0000;
array[40557] <= 16'b0000_0000_0000_0000;
array[40558] <= 16'b0000_0000_0000_0000;
array[40559] <= 16'b0000_0000_0000_0000;
array[40560] <= 16'b0000_0000_0000_0000;
array[40561] <= 16'b0000_0000_0000_0000;
array[40562] <= 16'b0000_0000_0000_0000;
array[40563] <= 16'b0000_0000_0000_0000;
array[40564] <= 16'b0000_0000_0000_0000;
array[40565] <= 16'b0000_0000_0000_0000;
array[40566] <= 16'b0000_0000_0000_0000;
array[40567] <= 16'b0000_0000_0000_0000;
array[40568] <= 16'b0000_0000_0000_0000;
array[40569] <= 16'b0000_0000_0000_0000;
array[40570] <= 16'b0000_0000_0000_0000;
array[40571] <= 16'b0000_0000_0000_0000;
array[40572] <= 16'b0000_0000_0000_0000;
array[40573] <= 16'b0000_0000_0000_0000;
array[40574] <= 16'b0000_0000_0000_0000;
array[40575] <= 16'b0000_0000_0000_0000;
array[40576] <= 16'b0000_0000_0000_0000;
array[40577] <= 16'b0000_0000_0000_0000;
array[40578] <= 16'b0000_0000_0000_0000;
array[40579] <= 16'b0000_0000_0000_0000;
array[40580] <= 16'b0000_0000_0000_0000;
array[40581] <= 16'b0000_0000_0000_0000;
array[40582] <= 16'b0000_0000_0000_0000;
array[40583] <= 16'b0000_0000_0000_0000;
array[40584] <= 16'b0000_0000_0000_0000;
array[40585] <= 16'b0000_0000_0000_0000;
array[40586] <= 16'b0000_0000_0000_0000;
array[40587] <= 16'b0000_0000_0000_0000;
array[40588] <= 16'b0000_0000_0000_0000;
array[40589] <= 16'b0000_0000_0000_0000;
array[40590] <= 16'b0000_0000_0000_0000;
array[40591] <= 16'b0000_0000_0000_0000;
array[40592] <= 16'b0000_0000_0000_0000;
array[40593] <= 16'b0000_0000_0000_0000;
array[40594] <= 16'b0000_0000_0000_0000;
array[40595] <= 16'b0000_0000_0000_0000;
array[40596] <= 16'b0000_0000_0000_0000;
array[40597] <= 16'b0000_0000_0000_0000;
array[40598] <= 16'b0000_0000_0000_0000;
array[40599] <= 16'b0000_0000_0000_0000;
array[40600] <= 16'b0000_0000_0000_0000;
array[40601] <= 16'b0000_0000_0000_0000;
array[40602] <= 16'b0000_0000_0000_0000;
array[40603] <= 16'b0000_0000_0000_0000;
array[40604] <= 16'b0000_0000_0000_0000;
array[40605] <= 16'b0000_0000_0000_0000;
array[40606] <= 16'b0000_0000_0000_0000;
array[40607] <= 16'b0000_0000_0000_0000;
array[40608] <= 16'b0000_0000_0000_0000;
array[40609] <= 16'b0000_0000_0000_0000;
array[40610] <= 16'b0000_0000_0000_0000;
array[40611] <= 16'b0000_0000_0000_0000;
array[40612] <= 16'b0000_0000_0000_0000;
array[40613] <= 16'b0000_0000_0000_0000;
array[40614] <= 16'b0000_0000_0000_0000;
array[40615] <= 16'b0000_0000_0000_0000;
array[40616] <= 16'b0000_0000_0000_0000;
array[40617] <= 16'b0000_0000_0000_0000;
array[40618] <= 16'b0000_0000_0000_0000;
array[40619] <= 16'b0000_0000_0000_0000;
array[40620] <= 16'b0000_0000_0000_0000;
array[40621] <= 16'b0000_0000_0000_0000;
array[40622] <= 16'b0000_0000_0000_0000;
array[40623] <= 16'b0000_0000_0000_0000;
array[40624] <= 16'b0000_0000_0000_0000;
array[40625] <= 16'b0000_0000_0000_0000;
array[40626] <= 16'b0000_0000_0000_0000;
array[40627] <= 16'b0000_0000_0000_0000;
array[40628] <= 16'b0000_0000_0000_0000;
array[40629] <= 16'b0000_0000_0000_0000;
array[40630] <= 16'b0000_0000_0000_0000;
array[40631] <= 16'b0000_0000_0000_0000;
array[40632] <= 16'b0000_0000_0000_0000;
array[40633] <= 16'b0000_0000_0000_0000;
array[40634] <= 16'b0000_0000_0000_0000;
array[40635] <= 16'b0000_0000_0000_0000;
array[40636] <= 16'b0000_0000_0000_0000;
array[40637] <= 16'b0000_0000_0000_0000;
array[40638] <= 16'b0000_0000_0000_0000;
array[40639] <= 16'b0000_0000_0000_0000;
array[40640] <= 16'b0000_0000_0000_0000;
array[40641] <= 16'b0000_0000_0000_0000;
array[40642] <= 16'b0000_0000_0000_0000;
array[40643] <= 16'b0000_0000_0000_0000;
array[40644] <= 16'b0000_0000_0000_0000;
array[40645] <= 16'b0000_0000_0000_0000;
array[40646] <= 16'b0000_0000_0000_0000;
array[40647] <= 16'b0000_0000_0000_0000;
array[40648] <= 16'b0000_0000_0000_0000;
array[40649] <= 16'b0000_0000_0000_0000;
array[40650] <= 16'b0000_0000_0000_0000;
array[40651] <= 16'b0000_0000_0000_0000;
array[40652] <= 16'b0000_0000_0000_0000;
array[40653] <= 16'b0000_0000_0000_0000;
array[40654] <= 16'b0000_0000_0000_0000;
array[40655] <= 16'b0000_0000_0000_0000;
array[40656] <= 16'b0000_0000_0000_0000;
array[40657] <= 16'b0000_0000_0000_0000;
array[40658] <= 16'b0000_0000_0000_0000;
array[40659] <= 16'b0000_0000_0000_0000;
array[40660] <= 16'b0000_0000_0000_0000;
array[40661] <= 16'b0000_0000_0000_0000;
array[40662] <= 16'b0000_0000_0000_0000;
array[40663] <= 16'b0000_0000_0000_0000;
array[40664] <= 16'b0000_0000_0000_0000;
array[40665] <= 16'b0000_0000_0000_0000;
array[40666] <= 16'b0000_0000_0000_0000;
array[40667] <= 16'b0000_0000_0000_0000;
array[40668] <= 16'b0000_0000_0000_0000;
array[40669] <= 16'b0000_0000_0000_0000;
array[40670] <= 16'b0000_0000_0000_0000;
array[40671] <= 16'b0000_0000_0000_0000;
array[40672] <= 16'b0000_0000_0000_0000;
array[40673] <= 16'b0000_0000_0000_0000;
array[40674] <= 16'b0000_0000_0000_0000;
array[40675] <= 16'b0000_0000_0000_0000;
array[40676] <= 16'b0000_0000_0000_0000;
array[40677] <= 16'b0000_0000_0000_0000;
array[40678] <= 16'b0000_0000_0000_0000;
array[40679] <= 16'b0000_0000_0000_0000;
array[40680] <= 16'b0000_0000_0000_0000;
array[40681] <= 16'b0000_0000_0000_0000;
array[40682] <= 16'b0000_0000_0000_0000;
array[40683] <= 16'b0000_0000_0000_0000;
array[40684] <= 16'b0000_0000_0000_0000;
array[40685] <= 16'b0000_0000_0000_0000;
array[40686] <= 16'b0000_0000_0000_0000;
array[40687] <= 16'b0000_0000_0000_0000;
array[40688] <= 16'b0000_0000_0000_0000;
array[40689] <= 16'b0000_0000_0000_0000;
array[40690] <= 16'b0000_0000_0000_0000;
array[40691] <= 16'b0000_0000_0000_0000;
array[40692] <= 16'b0000_0000_0000_0000;
array[40693] <= 16'b0000_0000_0000_0000;
array[40694] <= 16'b0000_0000_0000_0000;
array[40695] <= 16'b0000_0000_0000_0000;
array[40696] <= 16'b0000_0000_0000_0000;
array[40697] <= 16'b0000_0000_0000_0000;
array[40698] <= 16'b0000_0000_0000_0000;
array[40699] <= 16'b0000_0000_0000_0000;
array[40700] <= 16'b0000_0000_0000_0000;
array[40701] <= 16'b0000_0000_0000_0000;
array[40702] <= 16'b0000_0000_0000_0000;
array[40703] <= 16'b0000_0000_0000_0000;
array[40704] <= 16'b0000_0000_0000_0000;
array[40705] <= 16'b0000_0000_0000_0000;
array[40706] <= 16'b0000_0000_0000_0000;
array[40707] <= 16'b0000_0000_0000_0000;
array[40708] <= 16'b0000_0000_0000_0000;
array[40709] <= 16'b0000_0000_0000_0000;
array[40710] <= 16'b0000_0000_0000_0000;
array[40711] <= 16'b0000_0000_0000_0000;
array[40712] <= 16'b0000_0000_0000_0000;
array[40713] <= 16'b0000_0000_0000_0000;
array[40714] <= 16'b0000_0000_0000_0000;
array[40715] <= 16'b0000_0000_0000_0000;
array[40716] <= 16'b0000_0000_0000_0000;
array[40717] <= 16'b0000_0000_0000_0000;
array[40718] <= 16'b0000_0000_0000_0000;
array[40719] <= 16'b0000_0000_0000_0000;
array[40720] <= 16'b0000_0000_0000_0000;
array[40721] <= 16'b0000_0000_0000_0000;
array[40722] <= 16'b0000_0000_0000_0000;
array[40723] <= 16'b0000_0000_0000_0000;
array[40724] <= 16'b0000_0000_0000_0000;
array[40725] <= 16'b0000_0000_0000_0000;
array[40726] <= 16'b0000_0000_0000_0000;
array[40727] <= 16'b0000_0000_0000_0000;
array[40728] <= 16'b0000_0000_0000_0000;
array[40729] <= 16'b0000_0000_0000_0000;
array[40730] <= 16'b0000_0000_0000_0000;
array[40731] <= 16'b0000_0000_0000_0000;
array[40732] <= 16'b0000_0000_0000_0000;
array[40733] <= 16'b0000_0000_0000_0000;
array[40734] <= 16'b0000_0000_0000_0000;
array[40735] <= 16'b0000_0000_0000_0000;
array[40736] <= 16'b0000_0000_0000_0000;
array[40737] <= 16'b0000_0000_0000_0000;
array[40738] <= 16'b0000_0000_0000_0000;
array[40739] <= 16'b0000_0000_0000_0000;
array[40740] <= 16'b0000_0000_0000_0000;
array[40741] <= 16'b0000_0000_0000_0000;
array[40742] <= 16'b0000_0000_0000_0000;
array[40743] <= 16'b0000_0000_0000_0000;
array[40744] <= 16'b0000_0000_0000_0000;
array[40745] <= 16'b0000_0000_0000_0000;
array[40746] <= 16'b0000_0000_0000_0000;
array[40747] <= 16'b0000_0000_0000_0000;
array[40748] <= 16'b0000_0000_0000_0000;
array[40749] <= 16'b0000_0000_0000_0000;
array[40750] <= 16'b0000_0000_0000_0000;
array[40751] <= 16'b0000_0000_0000_0000;
array[40752] <= 16'b0000_0000_0000_0000;
array[40753] <= 16'b0000_0000_0000_0000;
array[40754] <= 16'b0000_0000_0000_0000;
array[40755] <= 16'b0000_0000_0000_0000;
array[40756] <= 16'b0000_0000_0000_0000;
array[40757] <= 16'b0000_0000_0000_0000;
array[40758] <= 16'b0000_0000_0000_0000;
array[40759] <= 16'b0000_0000_0000_0000;
array[40760] <= 16'b0000_0000_0000_0000;
array[40761] <= 16'b0000_0000_0000_0000;
array[40762] <= 16'b0000_0000_0000_0000;
array[40763] <= 16'b0000_0000_0000_0000;
array[40764] <= 16'b0000_0000_0000_0000;
array[40765] <= 16'b0000_0000_0000_0000;
array[40766] <= 16'b0000_0000_0000_0000;
array[40767] <= 16'b0000_0000_0000_0000;
array[40768] <= 16'b0000_0000_0000_0000;
array[40769] <= 16'b0000_0000_0000_0000;
array[40770] <= 16'b0000_0000_0000_0000;
array[40771] <= 16'b0000_0000_0000_0000;
array[40772] <= 16'b0000_0000_0000_0000;
array[40773] <= 16'b0000_0000_0000_0000;
array[40774] <= 16'b0000_0000_0000_0000;
array[40775] <= 16'b0000_0000_0000_0000;
array[40776] <= 16'b0000_0000_0000_0000;
array[40777] <= 16'b0000_0000_0000_0000;
array[40778] <= 16'b0000_0000_0000_0000;
array[40779] <= 16'b0000_0000_0000_0000;
array[40780] <= 16'b0000_0000_0000_0000;
array[40781] <= 16'b0000_0000_0000_0000;
array[40782] <= 16'b0000_0000_0000_0000;
array[40783] <= 16'b0000_0000_0000_0000;
array[40784] <= 16'b0000_0000_0000_0000;
array[40785] <= 16'b0000_0000_0000_0000;
array[40786] <= 16'b0000_0000_0000_0000;
array[40787] <= 16'b0000_0000_0000_0000;
array[40788] <= 16'b0000_0000_0000_0000;
array[40789] <= 16'b0000_0000_0000_0000;
array[40790] <= 16'b0000_0000_0000_0000;
array[40791] <= 16'b0000_0000_0000_0000;
array[40792] <= 16'b0000_0000_0000_0000;
array[40793] <= 16'b0000_0000_0000_0000;
array[40794] <= 16'b0000_0000_0000_0000;
array[40795] <= 16'b0000_0000_0000_0000;
array[40796] <= 16'b0000_0000_0000_0000;
array[40797] <= 16'b0000_0000_0000_0000;
array[40798] <= 16'b0000_0000_0000_0000;
array[40799] <= 16'b0000_0000_0000_0000;
array[40800] <= 16'b0000_0000_0000_0000;
array[40801] <= 16'b0000_0000_0000_0000;
array[40802] <= 16'b0000_0000_0000_0000;
array[40803] <= 16'b0000_0000_0000_0000;
array[40804] <= 16'b0000_0000_0000_0000;
array[40805] <= 16'b0000_0000_0000_0000;
array[40806] <= 16'b0000_0000_0000_0000;
array[40807] <= 16'b0000_0000_0000_0000;
array[40808] <= 16'b0000_0000_0000_0000;
array[40809] <= 16'b0000_0000_0000_0000;
array[40810] <= 16'b0000_0000_0000_0000;
array[40811] <= 16'b0000_0000_0000_0000;
array[40812] <= 16'b0000_0000_0000_0000;
array[40813] <= 16'b0000_0000_0000_0000;
array[40814] <= 16'b0000_0000_0000_0000;
array[40815] <= 16'b0000_0000_0000_0000;
array[40816] <= 16'b0000_0000_0000_0000;
array[40817] <= 16'b0000_0000_0000_0000;
array[40818] <= 16'b0000_0000_0000_0000;
array[40819] <= 16'b0000_0000_0000_0000;
array[40820] <= 16'b0000_0000_0000_0000;
array[40821] <= 16'b0000_0000_0000_0000;
array[40822] <= 16'b0000_0000_0000_0000;
array[40823] <= 16'b0000_0000_0000_0000;
array[40824] <= 16'b0000_0000_0000_0000;
array[40825] <= 16'b0000_0000_0000_0000;
array[40826] <= 16'b0000_0000_0000_0000;
array[40827] <= 16'b0000_0000_0000_0000;
array[40828] <= 16'b0000_0000_0000_0000;
array[40829] <= 16'b0000_0000_0000_0000;
array[40830] <= 16'b0000_0000_0000_0000;
array[40831] <= 16'b0000_0000_0000_0000;
array[40832] <= 16'b0000_0000_0000_0000;
array[40833] <= 16'b0000_0000_0000_0000;
array[40834] <= 16'b0000_0000_0000_0000;
array[40835] <= 16'b0000_0000_0000_0000;
array[40836] <= 16'b0000_0000_0000_0000;
array[40837] <= 16'b0000_0000_0000_0000;
array[40838] <= 16'b0000_0000_0000_0000;
array[40839] <= 16'b0000_0000_0000_0000;
array[40840] <= 16'b0000_0000_0000_0000;
array[40841] <= 16'b0000_0000_0000_0000;
array[40842] <= 16'b0000_0000_0000_0000;
array[40843] <= 16'b0000_0000_0000_0000;
array[40844] <= 16'b0000_0000_0000_0000;
array[40845] <= 16'b0000_0000_0000_0000;
array[40846] <= 16'b0000_0000_0000_0000;
array[40847] <= 16'b0000_0000_0000_0000;
array[40848] <= 16'b0000_0000_0000_0000;
array[40849] <= 16'b0000_0000_0000_0000;
array[40850] <= 16'b0000_0000_0000_0000;
array[40851] <= 16'b0000_0000_0000_0000;
array[40852] <= 16'b0000_0000_0000_0000;
array[40853] <= 16'b0000_0000_0000_0000;
array[40854] <= 16'b0000_0000_0000_0000;
array[40855] <= 16'b0000_0000_0000_0000;
array[40856] <= 16'b0000_0000_0000_0000;
array[40857] <= 16'b0000_0000_0000_0000;
array[40858] <= 16'b0000_0000_0000_0000;
array[40859] <= 16'b0000_0000_0000_0000;
array[40860] <= 16'b0000_0000_0000_0000;
array[40861] <= 16'b0000_0000_0000_0000;
array[40862] <= 16'b0000_0000_0000_0000;
array[40863] <= 16'b0000_0000_0000_0000;
array[40864] <= 16'b0000_0000_0000_0000;
array[40865] <= 16'b0000_0000_0000_0000;
array[40866] <= 16'b0000_0000_0000_0000;
array[40867] <= 16'b0000_0000_0000_0000;
array[40868] <= 16'b0000_0000_0000_0000;
array[40869] <= 16'b0000_0000_0000_0000;
array[40870] <= 16'b0000_0000_0000_0000;
array[40871] <= 16'b0000_0000_0000_0000;
array[40872] <= 16'b0000_0000_0000_0000;
array[40873] <= 16'b0000_0000_0000_0000;
array[40874] <= 16'b0000_0000_0000_0000;
array[40875] <= 16'b0000_0000_0000_0000;
array[40876] <= 16'b0000_0000_0000_0000;
array[40877] <= 16'b0000_0000_0000_0000;
array[40878] <= 16'b0000_0000_0000_0000;
array[40879] <= 16'b0000_0000_0000_0000;
array[40880] <= 16'b0000_0000_0000_0000;
array[40881] <= 16'b0000_0000_0000_0000;
array[40882] <= 16'b0000_0000_0000_0000;
array[40883] <= 16'b0000_0000_0000_0000;
array[40884] <= 16'b0000_0000_0000_0000;
array[40885] <= 16'b0000_0000_0000_0000;
array[40886] <= 16'b0000_0000_0000_0000;
array[40887] <= 16'b0000_0000_0000_0000;
array[40888] <= 16'b0000_0000_0000_0000;
array[40889] <= 16'b0000_0000_0000_0000;
array[40890] <= 16'b0000_0000_0000_0000;
array[40891] <= 16'b0000_0000_0000_0000;
array[40892] <= 16'b0000_0000_0000_0000;
array[40893] <= 16'b0000_0000_0000_0000;
array[40894] <= 16'b0000_0000_0000_0000;
array[40895] <= 16'b0000_0000_0000_0000;
array[40896] <= 16'b0000_0000_0000_0000;
array[40897] <= 16'b0000_0000_0000_0000;
array[40898] <= 16'b0000_0000_0000_0000;
array[40899] <= 16'b0000_0000_0000_0000;
array[40900] <= 16'b0000_0000_0000_0000;
array[40901] <= 16'b0000_0000_0000_0000;
array[40902] <= 16'b0000_0000_0000_0000;
array[40903] <= 16'b0000_0000_0000_0000;
array[40904] <= 16'b0000_0000_0000_0000;
array[40905] <= 16'b0000_0000_0000_0000;
array[40906] <= 16'b0000_0000_0000_0000;
array[40907] <= 16'b0000_0000_0000_0000;
array[40908] <= 16'b0000_0000_0000_0000;
array[40909] <= 16'b0000_0000_0000_0000;
array[40910] <= 16'b0000_0000_0000_0000;
array[40911] <= 16'b0000_0000_0000_0000;
array[40912] <= 16'b0000_0000_0000_0000;
array[40913] <= 16'b0000_0000_0000_0000;
array[40914] <= 16'b0000_0000_0000_0000;
array[40915] <= 16'b0000_0000_0000_0000;
array[40916] <= 16'b0000_0000_0000_0000;
array[40917] <= 16'b0000_0000_0000_0000;
array[40918] <= 16'b0000_0000_0000_0000;
array[40919] <= 16'b0000_0000_0000_0000;
array[40920] <= 16'b0000_0000_0000_0000;
array[40921] <= 16'b0000_0000_0000_0000;
array[40922] <= 16'b0000_0000_0000_0000;
array[40923] <= 16'b0000_0000_0000_0000;
array[40924] <= 16'b0000_0000_0000_0000;
array[40925] <= 16'b0000_0000_0000_0000;
array[40926] <= 16'b0000_0000_0000_0000;
array[40927] <= 16'b0000_0000_0000_0000;
array[40928] <= 16'b0000_0000_0000_0000;
array[40929] <= 16'b0000_0000_0000_0000;
array[40930] <= 16'b0000_0000_0000_0000;
array[40931] <= 16'b0000_0000_0000_0000;
array[40932] <= 16'b0000_0000_0000_0000;
array[40933] <= 16'b0000_0000_0000_0000;
array[40934] <= 16'b0000_0000_0000_0000;
array[40935] <= 16'b0000_0000_0000_0000;
array[40936] <= 16'b0000_0000_0000_0000;
array[40937] <= 16'b0000_0000_0000_0000;
array[40938] <= 16'b0000_0000_0000_0000;
array[40939] <= 16'b0000_0000_0000_0000;
array[40940] <= 16'b0000_0000_0000_0000;
array[40941] <= 16'b0000_0000_0000_0000;
array[40942] <= 16'b0000_0000_0000_0000;
array[40943] <= 16'b0000_0000_0000_0000;
array[40944] <= 16'b0000_0000_0000_0000;
array[40945] <= 16'b0000_0000_0000_0000;
array[40946] <= 16'b0000_0000_0000_0000;
array[40947] <= 16'b0000_0000_0000_0000;
array[40948] <= 16'b0000_0000_0000_0000;
array[40949] <= 16'b0000_0000_0000_0000;
array[40950] <= 16'b0000_0000_0000_0000;
array[40951] <= 16'b0000_0000_0000_0000;
array[40952] <= 16'b0000_0000_0000_0000;
array[40953] <= 16'b0000_0000_0000_0000;
array[40954] <= 16'b0000_0000_0000_0000;
array[40955] <= 16'b0000_0000_0000_0000;
array[40956] <= 16'b0000_0000_0000_0000;
array[40957] <= 16'b0000_0000_0000_0000;
array[40958] <= 16'b0000_0000_0000_0000;
array[40959] <= 16'b0000_0000_0000_0000;
array[40960] <= 16'b0000_0000_0000_0000;
array[40961] <= 16'b0000_0000_0000_0000;
array[40962] <= 16'b0000_0000_0000_0000;
array[40963] <= 16'b0000_0000_0000_0000;
array[40964] <= 16'b0000_0000_0000_0000;
array[40965] <= 16'b0000_0000_0000_0000;
array[40966] <= 16'b0000_0000_0000_0000;
array[40967] <= 16'b0000_0000_0000_0000;
array[40968] <= 16'b0000_0000_0000_0000;
array[40969] <= 16'b0000_0000_0000_0000;
array[40970] <= 16'b0000_0000_0000_0000;
array[40971] <= 16'b0000_0000_0000_0000;
array[40972] <= 16'b0000_0000_0000_0000;
array[40973] <= 16'b0000_0000_0000_0000;
array[40974] <= 16'b0000_0000_0000_0000;
array[40975] <= 16'b0000_0000_0000_0000;
array[40976] <= 16'b0000_0000_0000_0000;
array[40977] <= 16'b0000_0000_0000_0000;
array[40978] <= 16'b0000_0000_0000_0000;
array[40979] <= 16'b0000_0000_0000_0000;
array[40980] <= 16'b0000_0000_0000_0000;
array[40981] <= 16'b0000_0000_0000_0000;
array[40982] <= 16'b0000_0000_0000_0000;
array[40983] <= 16'b0000_0000_0000_0000;
array[40984] <= 16'b0000_0000_0000_0000;
array[40985] <= 16'b0000_0000_0000_0000;
array[40986] <= 16'b0000_0000_0000_0000;
array[40987] <= 16'b0000_0000_0000_0000;
array[40988] <= 16'b0000_0000_0000_0000;
array[40989] <= 16'b0000_0000_0000_0000;
array[40990] <= 16'b0000_0000_0000_0000;
array[40991] <= 16'b0000_0000_0000_0000;
array[40992] <= 16'b0000_0000_0000_0000;
array[40993] <= 16'b0000_0000_0000_0000;
array[40994] <= 16'b0000_0000_0000_0000;
array[40995] <= 16'b0000_0000_0000_0000;
array[40996] <= 16'b0000_0000_0000_0000;
array[40997] <= 16'b0000_0000_0000_0000;
array[40998] <= 16'b0000_0000_0000_0000;
array[40999] <= 16'b0000_0000_0000_0000;
array[41000] <= 16'b0000_0000_0000_0000;
array[41001] <= 16'b0000_0000_0000_0000;
array[41002] <= 16'b0000_0000_0000_0000;
array[41003] <= 16'b0000_0000_0000_0000;
array[41004] <= 16'b0000_0000_0000_0000;
array[41005] <= 16'b0000_0000_0000_0000;
array[41006] <= 16'b0000_0000_0000_0000;
array[41007] <= 16'b0000_0000_0000_0000;
array[41008] <= 16'b0000_0000_0000_0000;
array[41009] <= 16'b0000_0000_0000_0000;
array[41010] <= 16'b0000_0000_0000_0000;
array[41011] <= 16'b0000_0000_0000_0000;
array[41012] <= 16'b0000_0000_0000_0000;
array[41013] <= 16'b0000_0000_0000_0000;
array[41014] <= 16'b0000_0000_0000_0000;
array[41015] <= 16'b0000_0000_0000_0000;
array[41016] <= 16'b0000_0000_0000_0000;
array[41017] <= 16'b0000_0000_0000_0000;
array[41018] <= 16'b0000_0000_0000_0000;
array[41019] <= 16'b0000_0000_0000_0000;
array[41020] <= 16'b0000_0000_0000_0000;
array[41021] <= 16'b0000_0000_0000_0000;
array[41022] <= 16'b0000_0000_0000_0000;
array[41023] <= 16'b0000_0000_0000_0000;
array[41024] <= 16'b0000_0000_0000_0000;
array[41025] <= 16'b0000_0000_0000_0000;
array[41026] <= 16'b0000_0000_0000_0000;
array[41027] <= 16'b0000_0000_0000_0000;
array[41028] <= 16'b0000_0000_0000_0000;
array[41029] <= 16'b0000_0000_0000_0000;
array[41030] <= 16'b0000_0000_0000_0000;
array[41031] <= 16'b0000_0000_0000_0000;
array[41032] <= 16'b0000_0000_0000_0000;
array[41033] <= 16'b0000_0000_0000_0000;
array[41034] <= 16'b0000_0000_0000_0000;
array[41035] <= 16'b0000_0000_0000_0000;
array[41036] <= 16'b0000_0000_0000_0000;
array[41037] <= 16'b0000_0000_0000_0000;
array[41038] <= 16'b0000_0000_0000_0000;
array[41039] <= 16'b0000_0000_0000_0000;
array[41040] <= 16'b0000_0000_0000_0000;
array[41041] <= 16'b0000_0000_0000_0000;
array[41042] <= 16'b0000_0000_0000_0000;
array[41043] <= 16'b0000_0000_0000_0000;
array[41044] <= 16'b0000_0000_0000_0000;
array[41045] <= 16'b0000_0000_0000_0000;
array[41046] <= 16'b0000_0000_0000_0000;
array[41047] <= 16'b0000_0000_0000_0000;
array[41048] <= 16'b0000_0000_0000_0000;
array[41049] <= 16'b0000_0000_0000_0000;
array[41050] <= 16'b0000_0000_0000_0000;
array[41051] <= 16'b0000_0000_0000_0000;
array[41052] <= 16'b0000_0000_0000_0000;
array[41053] <= 16'b0000_0000_0000_0000;
array[41054] <= 16'b0000_0000_0000_0000;
array[41055] <= 16'b0000_0000_0000_0000;
array[41056] <= 16'b0000_0000_0000_0000;
array[41057] <= 16'b0000_0000_0000_0000;
array[41058] <= 16'b0000_0000_0000_0000;
array[41059] <= 16'b0000_0000_0000_0000;
array[41060] <= 16'b0000_0000_0000_0000;
array[41061] <= 16'b0000_0000_0000_0000;
array[41062] <= 16'b0000_0000_0000_0000;
array[41063] <= 16'b0000_0000_0000_0000;
array[41064] <= 16'b0000_0000_0000_0000;
array[41065] <= 16'b0000_0000_0000_0000;
array[41066] <= 16'b0000_0000_0000_0000;
array[41067] <= 16'b0000_0000_0000_0000;
array[41068] <= 16'b0000_0000_0000_0000;
array[41069] <= 16'b0000_0000_0000_0000;
array[41070] <= 16'b0000_0000_0000_0000;
array[41071] <= 16'b0000_0000_0000_0000;
array[41072] <= 16'b0000_0000_0000_0000;
array[41073] <= 16'b0000_0000_0000_0000;
array[41074] <= 16'b0000_0000_0000_0000;
array[41075] <= 16'b0000_0000_0000_0000;
array[41076] <= 16'b0000_0000_0000_0000;
array[41077] <= 16'b0000_0000_0000_0000;
array[41078] <= 16'b0000_0000_0000_0000;
array[41079] <= 16'b0000_0000_0000_0000;
array[41080] <= 16'b0000_0000_0000_0000;
array[41081] <= 16'b0000_0000_0000_0000;
array[41082] <= 16'b0000_0000_0000_0000;
array[41083] <= 16'b0000_0000_0000_0000;
array[41084] <= 16'b0000_0000_0000_0000;
array[41085] <= 16'b0000_0000_0000_0000;
array[41086] <= 16'b0000_0000_0000_0000;
array[41087] <= 16'b0000_0000_0000_0000;
array[41088] <= 16'b0000_0000_0000_0000;
array[41089] <= 16'b0000_0000_0000_0000;
array[41090] <= 16'b0000_0000_0000_0000;
array[41091] <= 16'b0000_0000_0000_0000;
array[41092] <= 16'b0000_0000_0000_0000;
array[41093] <= 16'b0000_0000_0000_0000;
array[41094] <= 16'b0000_0000_0000_0000;
array[41095] <= 16'b0000_0000_0000_0000;
array[41096] <= 16'b0000_0000_0000_0000;
array[41097] <= 16'b0000_0000_0000_0000;
array[41098] <= 16'b0000_0000_0000_0000;
array[41099] <= 16'b0000_0000_0000_0000;
array[41100] <= 16'b0000_0000_0000_0000;
array[41101] <= 16'b0000_0000_0000_0000;
array[41102] <= 16'b0000_0000_0000_0000;
array[41103] <= 16'b0000_0000_0000_0000;
array[41104] <= 16'b0000_0000_0000_0000;
array[41105] <= 16'b0000_0000_0000_0000;
array[41106] <= 16'b0000_0000_0000_0000;
array[41107] <= 16'b0000_0000_0000_0000;
array[41108] <= 16'b0000_0000_0000_0000;
array[41109] <= 16'b0000_0000_0000_0000;
array[41110] <= 16'b0000_0000_0000_0000;
array[41111] <= 16'b0000_0000_0000_0000;
array[41112] <= 16'b0000_0000_0000_0000;
array[41113] <= 16'b0000_0000_0000_0000;
array[41114] <= 16'b0000_0000_0000_0000;
array[41115] <= 16'b0000_0000_0000_0000;
array[41116] <= 16'b0000_0000_0000_0000;
array[41117] <= 16'b0000_0000_0000_0000;
array[41118] <= 16'b0000_0000_0000_0000;
array[41119] <= 16'b0000_0000_0000_0000;
array[41120] <= 16'b0000_0000_0000_0000;
array[41121] <= 16'b0000_0000_0000_0000;
array[41122] <= 16'b0000_0000_0000_0000;
array[41123] <= 16'b0000_0000_0000_0000;
array[41124] <= 16'b0000_0000_0000_0000;
array[41125] <= 16'b0000_0000_0000_0000;
array[41126] <= 16'b0000_0000_0000_0000;
array[41127] <= 16'b0000_0000_0000_0000;
array[41128] <= 16'b0000_0000_0000_0000;
array[41129] <= 16'b0000_0000_0000_0000;
array[41130] <= 16'b0000_0000_0000_0000;
array[41131] <= 16'b0000_0000_0000_0000;
array[41132] <= 16'b0000_0000_0000_0000;
array[41133] <= 16'b0000_0000_0000_0000;
array[41134] <= 16'b0000_0000_0000_0000;
array[41135] <= 16'b0000_0000_0000_0000;
array[41136] <= 16'b0000_0000_0000_0000;
array[41137] <= 16'b0000_0000_0000_0000;
array[41138] <= 16'b0000_0000_0000_0000;
array[41139] <= 16'b0000_0000_0000_0000;
array[41140] <= 16'b0000_0000_0000_0000;
array[41141] <= 16'b0000_0000_0000_0000;
array[41142] <= 16'b0000_0000_0000_0000;
array[41143] <= 16'b0000_0000_0000_0000;
array[41144] <= 16'b0000_0000_0000_0000;
array[41145] <= 16'b0000_0000_0000_0000;
array[41146] <= 16'b0000_0000_0000_0000;
array[41147] <= 16'b0000_0000_0000_0000;
array[41148] <= 16'b0000_0000_0000_0000;
array[41149] <= 16'b0000_0000_0000_0000;
array[41150] <= 16'b0000_0000_0000_0000;
array[41151] <= 16'b0000_0000_0000_0000;
array[41152] <= 16'b0000_0000_0000_0000;
array[41153] <= 16'b0000_0000_0000_0000;
array[41154] <= 16'b0000_0000_0000_0000;
array[41155] <= 16'b0000_0000_0000_0000;
array[41156] <= 16'b0000_0000_0000_0000;
array[41157] <= 16'b0000_0000_0000_0000;
array[41158] <= 16'b0000_0000_0000_0000;
array[41159] <= 16'b0000_0000_0000_0000;
array[41160] <= 16'b0000_0000_0000_0000;
array[41161] <= 16'b0000_0000_0000_0000;
array[41162] <= 16'b0000_0000_0000_0000;
array[41163] <= 16'b0000_0000_0000_0000;
array[41164] <= 16'b0000_0000_0000_0000;
array[41165] <= 16'b0000_0000_0000_0000;
array[41166] <= 16'b0000_0000_0000_0000;
array[41167] <= 16'b0000_0000_0000_0000;
array[41168] <= 16'b0000_0000_0000_0000;
array[41169] <= 16'b0000_0000_0000_0000;
array[41170] <= 16'b0000_0000_0000_0000;
array[41171] <= 16'b0000_0000_0000_0000;
array[41172] <= 16'b0000_0000_0000_0000;
array[41173] <= 16'b0000_0000_0000_0000;
array[41174] <= 16'b0000_0000_0000_0000;
array[41175] <= 16'b0000_0000_0000_0000;
array[41176] <= 16'b0000_0000_0000_0000;
array[41177] <= 16'b0000_0000_0000_0000;
array[41178] <= 16'b0000_0000_0000_0000;
array[41179] <= 16'b0000_0000_0000_0000;
array[41180] <= 16'b0000_0000_0000_0000;
array[41181] <= 16'b0000_0000_0000_0000;
array[41182] <= 16'b0000_0000_0000_0000;
array[41183] <= 16'b0000_0000_0000_0000;
array[41184] <= 16'b0000_0000_0000_0000;
array[41185] <= 16'b0000_0000_0000_0000;
array[41186] <= 16'b0000_0000_0000_0000;
array[41187] <= 16'b0000_0000_0000_0000;
array[41188] <= 16'b0000_0000_0000_0000;
array[41189] <= 16'b0000_0000_0000_0000;
array[41190] <= 16'b0000_0000_0000_0000;
array[41191] <= 16'b0000_0000_0000_0000;
array[41192] <= 16'b0000_0000_0000_0000;
array[41193] <= 16'b0000_0000_0000_0000;
array[41194] <= 16'b0000_0000_0000_0000;
array[41195] <= 16'b0000_0000_0000_0000;
array[41196] <= 16'b0000_0000_0000_0000;
array[41197] <= 16'b0000_0000_0000_0000;
array[41198] <= 16'b0000_0000_0000_0000;
array[41199] <= 16'b0000_0000_0000_0000;
array[41200] <= 16'b0000_0000_0000_0000;
array[41201] <= 16'b0000_0000_0000_0000;
array[41202] <= 16'b0000_0000_0000_0000;
array[41203] <= 16'b0000_0000_0000_0000;
array[41204] <= 16'b0000_0000_0000_0000;
array[41205] <= 16'b0000_0000_0000_0000;
array[41206] <= 16'b0000_0000_0000_0000;
array[41207] <= 16'b0000_0000_0000_0000;
array[41208] <= 16'b0000_0000_0000_0000;
array[41209] <= 16'b0000_0000_0000_0000;
array[41210] <= 16'b0000_0000_0000_0000;
array[41211] <= 16'b0000_0000_0000_0000;
array[41212] <= 16'b0000_0000_0000_0000;
array[41213] <= 16'b0000_0000_0000_0000;
array[41214] <= 16'b0000_0000_0000_0000;
array[41215] <= 16'b0000_0000_0000_0000;
array[41216] <= 16'b0000_0000_0000_0000;
array[41217] <= 16'b0000_0000_0000_0000;
array[41218] <= 16'b0000_0000_0000_0000;
array[41219] <= 16'b0000_0000_0000_0000;
array[41220] <= 16'b0000_0000_0000_0000;
array[41221] <= 16'b0000_0000_0000_0000;
array[41222] <= 16'b0000_0000_0000_0000;
array[41223] <= 16'b0000_0000_0000_0000;
array[41224] <= 16'b0000_0000_0000_0000;
array[41225] <= 16'b0000_0000_0000_0000;
array[41226] <= 16'b0000_0000_0000_0000;
array[41227] <= 16'b0000_0000_0000_0000;
array[41228] <= 16'b0000_0000_0000_0000;
array[41229] <= 16'b0000_0000_0000_0000;
array[41230] <= 16'b0000_0000_0000_0000;
array[41231] <= 16'b0000_0000_0000_0000;
array[41232] <= 16'b0000_0000_0000_0000;
array[41233] <= 16'b0000_0000_0000_0000;
array[41234] <= 16'b0000_0000_0000_0000;
array[41235] <= 16'b0000_0000_0000_0000;
array[41236] <= 16'b0000_0000_0000_0000;
array[41237] <= 16'b0000_0000_0000_0000;
array[41238] <= 16'b0000_0000_0000_0000;
array[41239] <= 16'b0000_0000_0000_0000;
array[41240] <= 16'b0000_0000_0000_0000;
array[41241] <= 16'b0000_0000_0000_0000;
array[41242] <= 16'b0000_0000_0000_0000;
array[41243] <= 16'b0000_0000_0000_0000;
array[41244] <= 16'b0000_0000_0000_0000;
array[41245] <= 16'b0000_0000_0000_0000;
array[41246] <= 16'b0000_0000_0000_0000;
array[41247] <= 16'b0000_0000_0000_0000;
array[41248] <= 16'b0000_0000_0000_0000;
array[41249] <= 16'b0000_0000_0000_0000;
array[41250] <= 16'b0000_0000_0000_0000;
array[41251] <= 16'b0000_0000_0000_0000;
array[41252] <= 16'b0000_0000_0000_0000;
array[41253] <= 16'b0000_0000_0000_0000;
array[41254] <= 16'b0000_0000_0000_0000;
array[41255] <= 16'b0000_0000_0000_0000;
array[41256] <= 16'b0000_0000_0000_0000;
array[41257] <= 16'b0000_0000_0000_0000;
array[41258] <= 16'b0000_0000_0000_0000;
array[41259] <= 16'b0000_0000_0000_0000;
array[41260] <= 16'b0000_0000_0000_0000;
array[41261] <= 16'b0000_0000_0000_0000;
array[41262] <= 16'b0000_0000_0000_0000;
array[41263] <= 16'b0000_0000_0000_0000;
array[41264] <= 16'b0000_0000_0000_0000;
array[41265] <= 16'b0000_0000_0000_0000;
array[41266] <= 16'b0000_0000_0000_0000;
array[41267] <= 16'b0000_0000_0000_0000;
array[41268] <= 16'b0000_0000_0000_0000;
array[41269] <= 16'b0000_0000_0000_0000;
array[41270] <= 16'b0000_0000_0000_0000;
array[41271] <= 16'b0000_0000_0000_0000;
array[41272] <= 16'b0000_0000_0000_0000;
array[41273] <= 16'b0000_0000_0000_0000;
array[41274] <= 16'b0000_0000_0000_0000;
array[41275] <= 16'b0000_0000_0000_0000;
array[41276] <= 16'b0000_0000_0000_0000;
array[41277] <= 16'b0000_0000_0000_0000;
array[41278] <= 16'b0000_0000_0000_0000;
array[41279] <= 16'b0000_0000_0000_0000;
array[41280] <= 16'b0000_0000_0000_0000;
array[41281] <= 16'b0000_0000_0000_0000;
array[41282] <= 16'b0000_0000_0000_0000;
array[41283] <= 16'b0000_0000_0000_0000;
array[41284] <= 16'b0000_0000_0000_0000;
array[41285] <= 16'b0000_0000_0000_0000;
array[41286] <= 16'b0000_0000_0000_0000;
array[41287] <= 16'b0000_0000_0000_0000;
array[41288] <= 16'b0000_0000_0000_0000;
array[41289] <= 16'b0000_0000_0000_0000;
array[41290] <= 16'b0000_0000_0000_0000;
array[41291] <= 16'b0000_0000_0000_0000;
array[41292] <= 16'b0000_0000_0000_0000;
array[41293] <= 16'b0000_0000_0000_0000;
array[41294] <= 16'b0000_0000_0000_0000;
array[41295] <= 16'b0000_0000_0000_0000;
array[41296] <= 16'b0000_0000_0000_0000;
array[41297] <= 16'b0000_0000_0000_0000;
array[41298] <= 16'b0000_0000_0000_0000;
array[41299] <= 16'b0000_0000_0000_0000;
array[41300] <= 16'b0000_0000_0000_0000;
array[41301] <= 16'b0000_0000_0000_0000;
array[41302] <= 16'b0000_0000_0000_0000;
array[41303] <= 16'b0000_0000_0000_0000;
array[41304] <= 16'b0000_0000_0000_0000;
array[41305] <= 16'b0000_0000_0000_0000;
array[41306] <= 16'b0000_0000_0000_0000;
array[41307] <= 16'b0000_0000_0000_0000;
array[41308] <= 16'b0000_0000_0000_0000;
array[41309] <= 16'b0000_0000_0000_0000;
array[41310] <= 16'b0000_0000_0000_0000;
array[41311] <= 16'b0000_0000_0000_0000;
array[41312] <= 16'b0000_0000_0000_0000;
array[41313] <= 16'b0000_0000_0000_0000;
array[41314] <= 16'b0000_0000_0000_0000;
array[41315] <= 16'b0000_0000_0000_0000;
array[41316] <= 16'b0000_0000_0000_0000;
array[41317] <= 16'b0000_0000_0000_0000;
array[41318] <= 16'b0000_0000_0000_0000;
array[41319] <= 16'b0000_0000_0000_0000;
array[41320] <= 16'b0000_0000_0000_0000;
array[41321] <= 16'b0000_0000_0000_0000;
array[41322] <= 16'b0000_0000_0000_0000;
array[41323] <= 16'b0000_0000_0000_0000;
array[41324] <= 16'b0000_0000_0000_0000;
array[41325] <= 16'b0000_0000_0000_0000;
array[41326] <= 16'b0000_0000_0000_0000;
array[41327] <= 16'b0000_0000_0000_0000;
array[41328] <= 16'b0000_0000_0000_0000;
array[41329] <= 16'b0000_0000_0000_0000;
array[41330] <= 16'b0000_0000_0000_0000;
array[41331] <= 16'b0000_0000_0000_0000;
array[41332] <= 16'b0000_0000_0000_0000;
array[41333] <= 16'b0000_0000_0000_0000;
array[41334] <= 16'b0000_0000_0000_0000;
array[41335] <= 16'b0000_0000_0000_0000;
array[41336] <= 16'b0000_0000_0000_0000;
array[41337] <= 16'b0000_0000_0000_0000;
array[41338] <= 16'b0000_0000_0000_0000;
array[41339] <= 16'b0000_0000_0000_0000;
array[41340] <= 16'b0000_0000_0000_0000;
array[41341] <= 16'b0000_0000_0000_0000;
array[41342] <= 16'b0000_0000_0000_0000;
array[41343] <= 16'b0000_0000_0000_0000;
array[41344] <= 16'b0000_0000_0000_0000;
array[41345] <= 16'b0000_0000_0000_0000;
array[41346] <= 16'b0000_0000_0000_0000;
array[41347] <= 16'b0000_0000_0000_0000;
array[41348] <= 16'b0000_0000_0000_0000;
array[41349] <= 16'b0000_0000_0000_0000;
array[41350] <= 16'b0000_0000_0000_0000;
array[41351] <= 16'b0000_0000_0000_0000;
array[41352] <= 16'b0000_0000_0000_0000;
array[41353] <= 16'b0000_0000_0000_0000;
array[41354] <= 16'b0000_0000_0000_0000;
array[41355] <= 16'b0000_0000_0000_0000;
array[41356] <= 16'b0000_0000_0000_0000;
array[41357] <= 16'b0000_0000_0000_0000;
array[41358] <= 16'b0000_0000_0000_0000;
array[41359] <= 16'b0000_0000_0000_0000;
array[41360] <= 16'b0000_0000_0000_0000;
array[41361] <= 16'b0000_0000_0000_0000;
array[41362] <= 16'b0000_0000_0000_0000;
array[41363] <= 16'b0000_0000_0000_0000;
array[41364] <= 16'b0000_0000_0000_0000;
array[41365] <= 16'b0000_0000_0000_0000;
array[41366] <= 16'b0000_0000_0000_0000;
array[41367] <= 16'b0000_0000_0000_0000;
array[41368] <= 16'b0000_0000_0000_0000;
array[41369] <= 16'b0000_0000_0000_0000;
array[41370] <= 16'b0000_0000_0000_0000;
array[41371] <= 16'b0000_0000_0000_0000;
array[41372] <= 16'b0000_0000_0000_0000;
array[41373] <= 16'b0000_0000_0000_0000;
array[41374] <= 16'b0000_0000_0000_0000;
array[41375] <= 16'b0000_0000_0000_0000;
array[41376] <= 16'b0000_0000_0000_0000;
array[41377] <= 16'b0000_0000_0000_0000;
array[41378] <= 16'b0000_0000_0000_0000;
array[41379] <= 16'b0000_0000_0000_0000;
array[41380] <= 16'b0000_0000_0000_0000;
array[41381] <= 16'b0000_0000_0000_0000;
array[41382] <= 16'b0000_0000_0000_0000;
array[41383] <= 16'b0000_0000_0000_0000;
array[41384] <= 16'b0000_0000_0000_0000;
array[41385] <= 16'b0000_0000_0000_0000;
array[41386] <= 16'b0000_0000_0000_0000;
array[41387] <= 16'b0000_0000_0000_0000;
array[41388] <= 16'b0000_0000_0000_0000;
array[41389] <= 16'b0000_0000_0000_0000;
array[41390] <= 16'b0000_0000_0000_0000;
array[41391] <= 16'b0000_0000_0000_0000;
array[41392] <= 16'b0000_0000_0000_0000;
array[41393] <= 16'b0000_0000_0000_0000;
array[41394] <= 16'b0000_0000_0000_0000;
array[41395] <= 16'b0000_0000_0000_0000;
array[41396] <= 16'b0000_0000_0000_0000;
array[41397] <= 16'b0000_0000_0000_0000;
array[41398] <= 16'b0000_0000_0000_0000;
array[41399] <= 16'b0000_0000_0000_0000;
array[41400] <= 16'b0000_0000_0000_0000;
array[41401] <= 16'b0000_0000_0000_0000;
array[41402] <= 16'b0000_0000_0000_0000;
array[41403] <= 16'b0000_0000_0000_0000;
array[41404] <= 16'b0000_0000_0000_0000;
array[41405] <= 16'b0000_0000_0000_0000;
array[41406] <= 16'b0000_0000_0000_0000;
array[41407] <= 16'b0000_0000_0000_0000;
array[41408] <= 16'b0000_0000_0000_0000;
array[41409] <= 16'b0000_0000_0000_0000;
array[41410] <= 16'b0000_0000_0000_0000;
array[41411] <= 16'b0000_0000_0000_0000;
array[41412] <= 16'b0000_0000_0000_0000;
array[41413] <= 16'b0000_0000_0000_0000;
array[41414] <= 16'b0000_0000_0000_0000;
array[41415] <= 16'b0000_0000_0000_0000;
array[41416] <= 16'b0000_0000_0000_0000;
array[41417] <= 16'b0000_0000_0000_0000;
array[41418] <= 16'b0000_0000_0000_0000;
array[41419] <= 16'b0000_0000_0000_0000;
array[41420] <= 16'b0000_0000_0000_0000;
array[41421] <= 16'b0000_0000_0000_0000;
array[41422] <= 16'b0000_0000_0000_0000;
array[41423] <= 16'b0000_0000_0000_0000;
array[41424] <= 16'b0000_0000_0000_0000;
array[41425] <= 16'b0000_0000_0000_0000;
array[41426] <= 16'b0000_0000_0000_0000;
array[41427] <= 16'b0000_0000_0000_0000;
array[41428] <= 16'b0000_0000_0000_0000;
array[41429] <= 16'b0000_0000_0000_0000;
array[41430] <= 16'b0000_0000_0000_0000;
array[41431] <= 16'b0000_0000_0000_0000;
array[41432] <= 16'b0000_0000_0000_0000;
array[41433] <= 16'b0000_0000_0000_0000;
array[41434] <= 16'b0000_0000_0000_0000;
array[41435] <= 16'b0000_0000_0000_0000;
array[41436] <= 16'b0000_0000_0000_0000;
array[41437] <= 16'b0000_0000_0000_0000;
array[41438] <= 16'b0000_0000_0000_0000;
array[41439] <= 16'b0000_0000_0000_0000;
array[41440] <= 16'b0000_0000_0000_0000;
array[41441] <= 16'b0000_0000_0000_0000;
array[41442] <= 16'b0000_0000_0000_0000;
array[41443] <= 16'b0000_0000_0000_0000;
array[41444] <= 16'b0000_0000_0000_0000;
array[41445] <= 16'b0000_0000_0000_0000;
array[41446] <= 16'b0000_0000_0000_0000;
array[41447] <= 16'b0000_0000_0000_0000;
array[41448] <= 16'b0000_0000_0000_0000;
array[41449] <= 16'b0000_0000_0000_0000;
array[41450] <= 16'b0000_0000_0000_0000;
array[41451] <= 16'b0000_0000_0000_0000;
array[41452] <= 16'b0000_0000_0000_0000;
array[41453] <= 16'b0000_0000_0000_0000;
array[41454] <= 16'b0000_0000_0000_0000;
array[41455] <= 16'b0000_0000_0000_0000;
array[41456] <= 16'b0000_0000_0000_0000;
array[41457] <= 16'b0000_0000_0000_0000;
array[41458] <= 16'b0000_0000_0000_0000;
array[41459] <= 16'b0000_0000_0000_0000;
array[41460] <= 16'b0000_0000_0000_0000;
array[41461] <= 16'b0000_0000_0000_0000;
array[41462] <= 16'b0000_0000_0000_0000;
array[41463] <= 16'b0000_0000_0000_0000;
array[41464] <= 16'b0000_0000_0000_0000;
array[41465] <= 16'b0000_0000_0000_0000;
array[41466] <= 16'b0000_0000_0000_0000;
array[41467] <= 16'b0000_0000_0000_0000;
array[41468] <= 16'b0000_0000_0000_0000;
array[41469] <= 16'b0000_0000_0000_0000;
array[41470] <= 16'b0000_0000_0000_0000;
array[41471] <= 16'b0000_0000_0000_0000;
array[41472] <= 16'b0000_0000_0000_0000;
array[41473] <= 16'b0000_0000_0000_0000;
array[41474] <= 16'b0000_0000_0000_0000;
array[41475] <= 16'b0000_0000_0000_0000;
array[41476] <= 16'b0000_0000_0000_0000;
array[41477] <= 16'b0000_0000_0000_0000;
array[41478] <= 16'b0000_0000_0000_0000;
array[41479] <= 16'b0000_0000_0000_0000;
array[41480] <= 16'b0000_0000_0000_0000;
array[41481] <= 16'b0000_0000_0000_0000;
array[41482] <= 16'b0000_0000_0000_0000;
array[41483] <= 16'b0000_0000_0000_0000;
array[41484] <= 16'b0000_0000_0000_0000;
array[41485] <= 16'b0000_0000_0000_0000;
array[41486] <= 16'b0000_0000_0000_0000;
array[41487] <= 16'b0000_0000_0000_0000;
array[41488] <= 16'b0000_0000_0000_0000;
array[41489] <= 16'b0000_0000_0000_0000;
array[41490] <= 16'b0000_0000_0000_0000;
array[41491] <= 16'b0000_0000_0000_0000;
array[41492] <= 16'b0000_0000_0000_0000;
array[41493] <= 16'b0000_0000_0000_0000;
array[41494] <= 16'b0000_0000_0000_0000;
array[41495] <= 16'b0000_0000_0000_0000;
array[41496] <= 16'b0000_0000_0000_0000;
array[41497] <= 16'b0000_0000_0000_0000;
array[41498] <= 16'b0000_0000_0000_0000;
array[41499] <= 16'b0000_0000_0000_0000;
array[41500] <= 16'b0000_0000_0000_0000;
array[41501] <= 16'b0000_0000_0000_0000;
array[41502] <= 16'b0000_0000_0000_0000;
array[41503] <= 16'b0000_0000_0000_0000;
array[41504] <= 16'b0000_0000_0000_0000;
array[41505] <= 16'b0000_0000_0000_0000;
array[41506] <= 16'b0000_0000_0000_0000;
array[41507] <= 16'b0000_0000_0000_0000;
array[41508] <= 16'b0000_0000_0000_0000;
array[41509] <= 16'b0000_0000_0000_0000;
array[41510] <= 16'b0000_0000_0000_0000;
array[41511] <= 16'b0000_0000_0000_0000;
array[41512] <= 16'b0000_0000_0000_0000;
array[41513] <= 16'b0000_0000_0000_0000;
array[41514] <= 16'b0000_0000_0000_0000;
array[41515] <= 16'b0000_0000_0000_0000;
array[41516] <= 16'b0000_0000_0000_0000;
array[41517] <= 16'b0000_0000_0000_0000;
array[41518] <= 16'b0000_0000_0000_0000;
array[41519] <= 16'b0000_0000_0000_0000;
array[41520] <= 16'b0000_0000_0000_0000;
array[41521] <= 16'b0000_0000_0000_0000;
array[41522] <= 16'b0000_0000_0000_0000;
array[41523] <= 16'b0000_0000_0000_0000;
array[41524] <= 16'b0000_0000_0000_0000;
array[41525] <= 16'b0000_0000_0000_0000;
array[41526] <= 16'b0000_0000_0000_0000;
array[41527] <= 16'b0000_0000_0000_0000;
array[41528] <= 16'b0000_0000_0000_0000;
array[41529] <= 16'b0000_0000_0000_0000;
array[41530] <= 16'b0000_0000_0000_0000;
array[41531] <= 16'b0000_0000_0000_0000;
array[41532] <= 16'b0000_0000_0000_0000;
array[41533] <= 16'b0000_0000_0000_0000;
array[41534] <= 16'b0000_0000_0000_0000;
array[41535] <= 16'b0000_0000_0000_0000;
array[41536] <= 16'b0000_0000_0000_0000;
array[41537] <= 16'b0000_0000_0000_0000;
array[41538] <= 16'b0000_0000_0000_0000;
array[41539] <= 16'b0000_0000_0000_0000;
array[41540] <= 16'b0000_0000_0000_0000;
array[41541] <= 16'b0000_0000_0000_0000;
array[41542] <= 16'b0000_0000_0000_0000;
array[41543] <= 16'b0000_0000_0000_0000;
array[41544] <= 16'b0000_0000_0000_0000;
array[41545] <= 16'b0000_0000_0000_0000;
array[41546] <= 16'b0000_0000_0000_0000;
array[41547] <= 16'b0000_0000_0000_0000;
array[41548] <= 16'b0000_0000_0000_0000;
array[41549] <= 16'b0000_0000_0000_0000;
array[41550] <= 16'b0000_0000_0000_0000;
array[41551] <= 16'b0000_0000_0000_0000;
array[41552] <= 16'b0000_0000_0000_0000;
array[41553] <= 16'b0000_0000_0000_0000;
array[41554] <= 16'b0000_0000_0000_0000;
array[41555] <= 16'b0000_0000_0000_0000;
array[41556] <= 16'b0000_0000_0000_0000;
array[41557] <= 16'b0000_0000_0000_0000;
array[41558] <= 16'b0000_0000_0000_0000;
array[41559] <= 16'b0000_0000_0000_0000;
array[41560] <= 16'b0000_0000_0000_0000;
array[41561] <= 16'b0000_0000_0000_0000;
array[41562] <= 16'b0000_0000_0000_0000;
array[41563] <= 16'b0000_0000_0000_0000;
array[41564] <= 16'b0000_0000_0000_0000;
array[41565] <= 16'b0000_0000_0000_0000;
array[41566] <= 16'b0000_0000_0000_0000;
array[41567] <= 16'b0000_0000_0000_0000;
array[41568] <= 16'b0000_0000_0000_0000;
array[41569] <= 16'b0000_0000_0000_0000;
array[41570] <= 16'b0000_0000_0000_0000;
array[41571] <= 16'b0000_0000_0000_0000;
array[41572] <= 16'b0000_0000_0000_0000;
array[41573] <= 16'b0000_0000_0000_0000;
array[41574] <= 16'b0000_0000_0000_0000;
array[41575] <= 16'b0000_0000_0000_0000;
array[41576] <= 16'b0000_0000_0000_0000;
array[41577] <= 16'b0000_0000_0000_0000;
array[41578] <= 16'b0000_0000_0000_0000;
array[41579] <= 16'b0000_0000_0000_0000;
array[41580] <= 16'b0000_0000_0000_0000;
array[41581] <= 16'b0000_0000_0000_0000;
array[41582] <= 16'b0000_0000_0000_0000;
array[41583] <= 16'b0000_0000_0000_0000;
array[41584] <= 16'b0000_0000_0000_0000;
array[41585] <= 16'b0000_0000_0000_0000;
array[41586] <= 16'b0000_0000_0000_0000;
array[41587] <= 16'b0000_0000_0000_0000;
array[41588] <= 16'b0000_0000_0000_0000;
array[41589] <= 16'b0000_0000_0000_0000;
array[41590] <= 16'b0000_0000_0000_0000;
array[41591] <= 16'b0000_0000_0000_0000;
array[41592] <= 16'b0000_0000_0000_0000;
array[41593] <= 16'b0000_0000_0000_0000;
array[41594] <= 16'b0000_0000_0000_0000;
array[41595] <= 16'b0000_0000_0000_0000;
array[41596] <= 16'b0000_0000_0000_0000;
array[41597] <= 16'b0000_0000_0000_0000;
array[41598] <= 16'b0000_0000_0000_0000;
array[41599] <= 16'b0000_0000_0000_0000;
array[41600] <= 16'b0000_0000_0000_0000;
array[41601] <= 16'b0000_0000_0000_0000;
array[41602] <= 16'b0000_0000_0000_0000;
array[41603] <= 16'b0000_0000_0000_0000;
array[41604] <= 16'b0000_0000_0000_0000;
array[41605] <= 16'b0000_0000_0000_0000;
array[41606] <= 16'b0000_0000_0000_0000;
array[41607] <= 16'b0000_0000_0000_0000;
array[41608] <= 16'b0000_0000_0000_0000;
array[41609] <= 16'b0000_0000_0000_0000;
array[41610] <= 16'b0000_0000_0000_0000;
array[41611] <= 16'b0000_0000_0000_0000;
array[41612] <= 16'b0000_0000_0000_0000;
array[41613] <= 16'b0000_0000_0000_0000;
array[41614] <= 16'b0000_0000_0000_0000;
array[41615] <= 16'b0000_0000_0000_0000;
array[41616] <= 16'b0000_0000_0000_0000;
array[41617] <= 16'b0000_0000_0000_0000;
array[41618] <= 16'b0000_0000_0000_0000;
array[41619] <= 16'b0000_0000_0000_0000;
array[41620] <= 16'b0000_0000_0000_0000;
array[41621] <= 16'b0000_0000_0000_0000;
array[41622] <= 16'b0000_0000_0000_0000;
array[41623] <= 16'b0000_0000_0000_0000;
array[41624] <= 16'b0000_0000_0000_0000;
array[41625] <= 16'b0000_0000_0000_0000;
array[41626] <= 16'b0000_0000_0000_0000;
array[41627] <= 16'b0000_0000_0000_0000;
array[41628] <= 16'b0000_0000_0000_0000;
array[41629] <= 16'b0000_0000_0000_0000;
array[41630] <= 16'b0000_0000_0000_0000;
array[41631] <= 16'b0000_0000_0000_0000;
array[41632] <= 16'b0000_0000_0000_0000;
array[41633] <= 16'b0000_0000_0000_0000;
array[41634] <= 16'b0000_0000_0000_0000;
array[41635] <= 16'b0000_0000_0000_0000;
array[41636] <= 16'b0000_0000_0000_0000;
array[41637] <= 16'b0000_0000_0000_0000;
array[41638] <= 16'b0000_0000_0000_0000;
array[41639] <= 16'b0000_0000_0000_0000;
array[41640] <= 16'b0000_0000_0000_0000;
array[41641] <= 16'b0000_0000_0000_0000;
array[41642] <= 16'b0000_0000_0000_0000;
array[41643] <= 16'b0000_0000_0000_0000;
array[41644] <= 16'b0000_0000_0000_0000;
array[41645] <= 16'b0000_0000_0000_0000;
array[41646] <= 16'b0000_0000_0000_0000;
array[41647] <= 16'b0000_0000_0000_0000;
array[41648] <= 16'b0000_0000_0000_0000;
array[41649] <= 16'b0000_0000_0000_0000;
array[41650] <= 16'b0000_0000_0000_0000;
array[41651] <= 16'b0000_0000_0000_0000;
array[41652] <= 16'b0000_0000_0000_0000;
array[41653] <= 16'b0000_0000_0000_0000;
array[41654] <= 16'b0000_0000_0000_0000;
array[41655] <= 16'b0000_0000_0000_0000;
array[41656] <= 16'b0000_0000_0000_0000;
array[41657] <= 16'b0000_0000_0000_0000;
array[41658] <= 16'b0000_0000_0000_0000;
array[41659] <= 16'b0000_0000_0000_0000;
array[41660] <= 16'b0000_0000_0000_0000;
array[41661] <= 16'b0000_0000_0000_0000;
array[41662] <= 16'b0000_0000_0000_0000;
array[41663] <= 16'b0000_0000_0000_0000;
array[41664] <= 16'b0000_0000_0000_0000;
array[41665] <= 16'b0000_0000_0000_0000;
array[41666] <= 16'b0000_0000_0000_0000;
array[41667] <= 16'b0000_0000_0000_0000;
array[41668] <= 16'b0000_0000_0000_0000;
array[41669] <= 16'b0000_0000_0000_0000;
array[41670] <= 16'b0000_0000_0000_0000;
array[41671] <= 16'b0000_0000_0000_0000;
array[41672] <= 16'b0000_0000_0000_0000;
array[41673] <= 16'b0000_0000_0000_0000;
array[41674] <= 16'b0000_0000_0000_0000;
array[41675] <= 16'b0000_0000_0000_0000;
array[41676] <= 16'b0000_0000_0000_0000;
array[41677] <= 16'b0000_0000_0000_0000;
array[41678] <= 16'b0000_0000_0000_0000;
array[41679] <= 16'b0000_0000_0000_0000;
array[41680] <= 16'b0000_0000_0000_0000;
array[41681] <= 16'b0000_0000_0000_0000;
array[41682] <= 16'b0000_0000_0000_0000;
array[41683] <= 16'b0000_0000_0000_0000;
array[41684] <= 16'b0000_0000_0000_0000;
array[41685] <= 16'b0000_0000_0000_0000;
array[41686] <= 16'b0000_0000_0000_0000;
array[41687] <= 16'b0000_0000_0000_0000;
array[41688] <= 16'b0000_0000_0000_0000;
array[41689] <= 16'b0000_0000_0000_0000;
array[41690] <= 16'b0000_0000_0000_0000;
array[41691] <= 16'b0000_0000_0000_0000;
array[41692] <= 16'b0000_0000_0000_0000;
array[41693] <= 16'b0000_0000_0000_0000;
array[41694] <= 16'b0000_0000_0000_0000;
array[41695] <= 16'b0000_0000_0000_0000;
array[41696] <= 16'b0000_0000_0000_0000;
array[41697] <= 16'b0000_0000_0000_0000;
array[41698] <= 16'b0000_0000_0000_0000;
array[41699] <= 16'b0000_0000_0000_0000;
array[41700] <= 16'b0000_0000_0000_0000;
array[41701] <= 16'b0000_0000_0000_0000;
array[41702] <= 16'b0000_0000_0000_0000;
array[41703] <= 16'b0000_0000_0000_0000;
array[41704] <= 16'b0000_0000_0000_0000;
array[41705] <= 16'b0000_0000_0000_0000;
array[41706] <= 16'b0000_0000_0000_0000;
array[41707] <= 16'b0000_0000_0000_0000;
array[41708] <= 16'b0000_0000_0000_0000;
array[41709] <= 16'b0000_0000_0000_0000;
array[41710] <= 16'b0000_0000_0000_0000;
array[41711] <= 16'b0000_0000_0000_0000;
array[41712] <= 16'b0000_0000_0000_0000;
array[41713] <= 16'b0000_0000_0000_0000;
array[41714] <= 16'b0000_0000_0000_0000;
array[41715] <= 16'b0000_0000_0000_0000;
array[41716] <= 16'b0000_0000_0000_0000;
array[41717] <= 16'b0000_0000_0000_0000;
array[41718] <= 16'b0000_0000_0000_0000;
array[41719] <= 16'b0000_0000_0000_0000;
array[41720] <= 16'b0000_0000_0000_0000;
array[41721] <= 16'b0000_0000_0000_0000;
array[41722] <= 16'b0000_0000_0000_0000;
array[41723] <= 16'b0000_0000_0000_0000;
array[41724] <= 16'b0000_0000_0000_0000;
array[41725] <= 16'b0000_0000_0000_0000;
array[41726] <= 16'b0000_0000_0000_0000;
array[41727] <= 16'b0000_0000_0000_0000;
array[41728] <= 16'b0000_0000_0000_0000;
array[41729] <= 16'b0000_0000_0000_0000;
array[41730] <= 16'b0000_0000_0000_0000;
array[41731] <= 16'b0000_0000_0000_0000;
array[41732] <= 16'b0000_0000_0000_0000;
array[41733] <= 16'b0000_0000_0000_0000;
array[41734] <= 16'b0000_0000_0000_0000;
array[41735] <= 16'b0000_0000_0000_0000;
array[41736] <= 16'b0000_0000_0000_0000;
array[41737] <= 16'b0000_0000_0000_0000;
array[41738] <= 16'b0000_0000_0000_0000;
array[41739] <= 16'b0000_0000_0000_0000;
array[41740] <= 16'b0000_0000_0000_0000;
array[41741] <= 16'b0000_0000_0000_0000;
array[41742] <= 16'b0000_0000_0000_0000;
array[41743] <= 16'b0000_0000_0000_0000;
array[41744] <= 16'b0000_0000_0000_0000;
array[41745] <= 16'b0000_0000_0000_0000;
array[41746] <= 16'b0000_0000_0000_0000;
array[41747] <= 16'b0000_0000_0000_0000;
array[41748] <= 16'b0000_0000_0000_0000;
array[41749] <= 16'b0000_0000_0000_0000;
array[41750] <= 16'b0000_0000_0000_0000;
array[41751] <= 16'b0000_0000_0000_0000;
array[41752] <= 16'b0000_0000_0000_0000;
array[41753] <= 16'b0000_0000_0000_0000;
array[41754] <= 16'b0000_0000_0000_0000;
array[41755] <= 16'b0000_0000_0000_0000;
array[41756] <= 16'b0000_0000_0000_0000;
array[41757] <= 16'b0000_0000_0000_0000;
array[41758] <= 16'b0000_0000_0000_0000;
array[41759] <= 16'b0000_0000_0000_0000;
array[41760] <= 16'b0000_0000_0000_0000;
array[41761] <= 16'b0000_0000_0000_0000;
array[41762] <= 16'b0000_0000_0000_0000;
array[41763] <= 16'b0000_0000_0000_0000;
array[41764] <= 16'b0000_0000_0000_0000;
array[41765] <= 16'b0000_0000_0000_0000;
array[41766] <= 16'b0000_0000_0000_0000;
array[41767] <= 16'b0000_0000_0000_0000;
array[41768] <= 16'b0000_0000_0000_0000;
array[41769] <= 16'b0000_0000_0000_0000;
array[41770] <= 16'b0000_0000_0000_0000;
array[41771] <= 16'b0000_0000_0000_0000;
array[41772] <= 16'b0000_0000_0000_0000;
array[41773] <= 16'b0000_0000_0000_0000;
array[41774] <= 16'b0000_0000_0000_0000;
array[41775] <= 16'b0000_0000_0000_0000;
array[41776] <= 16'b0000_0000_0000_0000;
array[41777] <= 16'b0000_0000_0000_0000;
array[41778] <= 16'b0000_0000_0000_0000;
array[41779] <= 16'b0000_0000_0000_0000;
array[41780] <= 16'b0000_0000_0000_0000;
array[41781] <= 16'b0000_0000_0000_0000;
array[41782] <= 16'b0000_0000_0000_0000;
array[41783] <= 16'b0000_0000_0000_0000;
array[41784] <= 16'b0000_0000_0000_0000;
array[41785] <= 16'b0000_0000_0000_0000;
array[41786] <= 16'b0000_0000_0000_0000;
array[41787] <= 16'b0000_0000_0000_0000;
array[41788] <= 16'b0000_0000_0000_0000;
array[41789] <= 16'b0000_0000_0000_0000;
array[41790] <= 16'b0000_0000_0000_0000;
array[41791] <= 16'b0000_0000_0000_0000;
array[41792] <= 16'b0000_0000_0000_0000;
array[41793] <= 16'b0000_0000_0000_0000;
array[41794] <= 16'b0000_0000_0000_0000;
array[41795] <= 16'b0000_0000_0000_0000;
array[41796] <= 16'b0000_0000_0000_0000;
array[41797] <= 16'b0000_0000_0000_0000;
array[41798] <= 16'b0000_0000_0000_0000;
array[41799] <= 16'b0000_0000_0000_0000;
array[41800] <= 16'b0000_0000_0000_0000;
array[41801] <= 16'b0000_0000_0000_0000;
array[41802] <= 16'b0000_0000_0000_0000;
array[41803] <= 16'b0000_0000_0000_0000;
array[41804] <= 16'b0000_0000_0000_0000;
array[41805] <= 16'b0000_0000_0000_0000;
array[41806] <= 16'b0000_0000_0000_0000;
array[41807] <= 16'b0000_0000_0000_0000;
array[41808] <= 16'b0000_0000_0000_0000;
array[41809] <= 16'b0000_0000_0000_0000;
array[41810] <= 16'b0000_0000_0000_0000;
array[41811] <= 16'b0000_0000_0000_0000;
array[41812] <= 16'b0000_0000_0000_0000;
array[41813] <= 16'b0000_0000_0000_0000;
array[41814] <= 16'b0000_0000_0000_0000;
array[41815] <= 16'b0000_0000_0000_0000;
array[41816] <= 16'b0000_0000_0000_0000;
array[41817] <= 16'b0000_0000_0000_0000;
array[41818] <= 16'b0000_0000_0000_0000;
array[41819] <= 16'b0000_0000_0000_0000;
array[41820] <= 16'b0000_0000_0000_0000;
array[41821] <= 16'b0000_0000_0000_0000;
array[41822] <= 16'b0000_0000_0000_0000;
array[41823] <= 16'b0000_0000_0000_0000;
array[41824] <= 16'b0000_0000_0000_0000;
array[41825] <= 16'b0000_0000_0000_0000;
array[41826] <= 16'b0000_0000_0000_0000;
array[41827] <= 16'b0000_0000_0000_0000;
array[41828] <= 16'b0000_0000_0000_0000;
array[41829] <= 16'b0000_0000_0000_0000;
array[41830] <= 16'b0000_0000_0000_0000;
array[41831] <= 16'b0000_0000_0000_0000;
array[41832] <= 16'b0000_0000_0000_0000;
array[41833] <= 16'b0000_0000_0000_0000;
array[41834] <= 16'b0000_0000_0000_0000;
array[41835] <= 16'b0000_0000_0000_0000;
array[41836] <= 16'b0000_0000_0000_0000;
array[41837] <= 16'b0000_0000_0000_0000;
array[41838] <= 16'b0000_0000_0000_0000;
array[41839] <= 16'b0000_0000_0000_0000;
array[41840] <= 16'b0000_0000_0000_0000;
array[41841] <= 16'b0000_0000_0000_0000;
array[41842] <= 16'b0000_0000_0000_0000;
array[41843] <= 16'b0000_0000_0000_0000;
array[41844] <= 16'b0000_0000_0000_0000;
array[41845] <= 16'b0000_0000_0000_0000;
array[41846] <= 16'b0000_0000_0000_0000;
array[41847] <= 16'b0000_0000_0000_0000;
array[41848] <= 16'b0000_0000_0000_0000;
array[41849] <= 16'b0000_0000_0000_0000;
array[41850] <= 16'b0000_0000_0000_0000;
array[41851] <= 16'b0000_0000_0000_0000;
array[41852] <= 16'b0000_0000_0000_0000;
array[41853] <= 16'b0000_0000_0000_0000;
array[41854] <= 16'b0000_0000_0000_0000;
array[41855] <= 16'b0000_0000_0000_0000;
array[41856] <= 16'b0000_0000_0000_0000;
array[41857] <= 16'b0000_0000_0000_0000;
array[41858] <= 16'b0000_0000_0000_0000;
array[41859] <= 16'b0000_0000_0000_0000;
array[41860] <= 16'b0000_0000_0000_0000;
array[41861] <= 16'b0000_0000_0000_0000;
array[41862] <= 16'b0000_0000_0000_0000;
array[41863] <= 16'b0000_0000_0000_0000;
array[41864] <= 16'b0000_0000_0000_0000;
array[41865] <= 16'b0000_0000_0000_0000;
array[41866] <= 16'b0000_0000_0000_0000;
array[41867] <= 16'b0000_0000_0000_0000;
array[41868] <= 16'b0000_0000_0000_0000;
array[41869] <= 16'b0000_0000_0000_0000;
array[41870] <= 16'b0000_0000_0000_0000;
array[41871] <= 16'b0000_0000_0000_0000;
array[41872] <= 16'b0000_0000_0000_0000;
array[41873] <= 16'b0000_0000_0000_0000;
array[41874] <= 16'b0000_0000_0000_0000;
array[41875] <= 16'b0000_0000_0000_0000;
array[41876] <= 16'b0000_0000_0000_0000;
array[41877] <= 16'b0000_0000_0000_0000;
array[41878] <= 16'b0000_0000_0000_0000;
array[41879] <= 16'b0000_0000_0000_0000;
array[41880] <= 16'b0000_0000_0000_0000;
array[41881] <= 16'b0000_0000_0000_0000;
array[41882] <= 16'b0000_0000_0000_0000;
array[41883] <= 16'b0000_0000_0000_0000;
array[41884] <= 16'b0000_0000_0000_0000;
array[41885] <= 16'b0000_0000_0000_0000;
array[41886] <= 16'b0000_0000_0000_0000;
array[41887] <= 16'b0000_0000_0000_0000;
array[41888] <= 16'b0000_0000_0000_0000;
array[41889] <= 16'b0000_0000_0000_0000;
array[41890] <= 16'b0000_0000_0000_0000;
array[41891] <= 16'b0000_0000_0000_0000;
array[41892] <= 16'b0000_0000_0000_0000;
array[41893] <= 16'b0000_0000_0000_0000;
array[41894] <= 16'b0000_0000_0000_0000;
array[41895] <= 16'b0000_0000_0000_0000;
array[41896] <= 16'b0000_0000_0000_0000;
array[41897] <= 16'b0000_0000_0000_0000;
array[41898] <= 16'b0000_0000_0000_0000;
array[41899] <= 16'b0000_0000_0000_0000;
array[41900] <= 16'b0000_0000_0000_0000;
array[41901] <= 16'b0000_0000_0000_0000;
array[41902] <= 16'b0000_0000_0000_0000;
array[41903] <= 16'b0000_0000_0000_0000;
array[41904] <= 16'b0000_0000_0000_0000;
array[41905] <= 16'b0000_0000_0000_0000;
array[41906] <= 16'b0000_0000_0000_0000;
array[41907] <= 16'b0000_0000_0000_0000;
array[41908] <= 16'b0000_0000_0000_0000;
array[41909] <= 16'b0000_0000_0000_0000;
array[41910] <= 16'b0000_0000_0000_0000;
array[41911] <= 16'b0000_0000_0000_0000;
array[41912] <= 16'b0000_0000_0000_0000;
array[41913] <= 16'b0000_0000_0000_0000;
array[41914] <= 16'b0000_0000_0000_0000;
array[41915] <= 16'b0000_0000_0000_0000;
array[41916] <= 16'b0000_0000_0000_0000;
array[41917] <= 16'b0000_0000_0000_0000;
array[41918] <= 16'b0000_0000_0000_0000;
array[41919] <= 16'b0000_0000_0000_0000;
array[41920] <= 16'b0000_0000_0000_0000;
array[41921] <= 16'b0000_0000_0000_0000;
array[41922] <= 16'b0000_0000_0000_0000;
array[41923] <= 16'b0000_0000_0000_0000;
array[41924] <= 16'b0000_0000_0000_0000;
array[41925] <= 16'b0000_0000_0000_0000;
array[41926] <= 16'b0000_0000_0000_0000;
array[41927] <= 16'b0000_0000_0000_0000;
array[41928] <= 16'b0000_0000_0000_0000;
array[41929] <= 16'b0000_0000_0000_0000;
array[41930] <= 16'b0000_0000_0000_0000;
array[41931] <= 16'b0000_0000_0000_0000;
array[41932] <= 16'b0000_0000_0000_0000;
array[41933] <= 16'b0000_0000_0000_0000;
array[41934] <= 16'b0000_0000_0000_0000;
array[41935] <= 16'b0000_0000_0000_0000;
array[41936] <= 16'b0000_0000_0000_0000;
array[41937] <= 16'b0000_0000_0000_0000;
array[41938] <= 16'b0000_0000_0000_0000;
array[41939] <= 16'b0000_0000_0000_0000;
array[41940] <= 16'b0000_0000_0000_0000;
array[41941] <= 16'b0000_0000_0000_0000;
array[41942] <= 16'b0000_0000_0000_0000;
array[41943] <= 16'b0000_0000_0000_0000;
array[41944] <= 16'b0000_0000_0000_0000;
array[41945] <= 16'b0000_0000_0000_0000;
array[41946] <= 16'b0000_0000_0000_0000;
array[41947] <= 16'b0000_0000_0000_0000;
array[41948] <= 16'b0000_0000_0000_0000;
array[41949] <= 16'b0000_0000_0000_0000;
array[41950] <= 16'b0000_0000_0000_0000;
array[41951] <= 16'b0000_0000_0000_0000;
array[41952] <= 16'b0000_0000_0000_0000;
array[41953] <= 16'b0000_0000_0000_0000;
array[41954] <= 16'b0000_0000_0000_0000;
array[41955] <= 16'b0000_0000_0000_0000;
array[41956] <= 16'b0000_0000_0000_0000;
array[41957] <= 16'b0000_0000_0000_0000;
array[41958] <= 16'b0000_0000_0000_0000;
array[41959] <= 16'b0000_0000_0000_0000;
array[41960] <= 16'b0000_0000_0000_0000;
array[41961] <= 16'b0000_0000_0000_0000;
array[41962] <= 16'b0000_0000_0000_0000;
array[41963] <= 16'b0000_0000_0000_0000;
array[41964] <= 16'b0000_0000_0000_0000;
array[41965] <= 16'b0000_0000_0000_0000;
array[41966] <= 16'b0000_0000_0000_0000;
array[41967] <= 16'b0000_0000_0000_0000;
array[41968] <= 16'b0000_0000_0000_0000;
array[41969] <= 16'b0000_0000_0000_0000;
array[41970] <= 16'b0000_0000_0000_0000;
array[41971] <= 16'b0000_0000_0000_0000;
array[41972] <= 16'b0000_0000_0000_0000;
array[41973] <= 16'b0000_0000_0000_0000;
array[41974] <= 16'b0000_0000_0000_0000;
array[41975] <= 16'b0000_0000_0000_0000;
array[41976] <= 16'b0000_0000_0000_0000;
array[41977] <= 16'b0000_0000_0000_0000;
array[41978] <= 16'b0000_0000_0000_0000;
array[41979] <= 16'b0000_0000_0000_0000;
array[41980] <= 16'b0000_0000_0000_0000;
array[41981] <= 16'b0000_0000_0000_0000;
array[41982] <= 16'b0000_0000_0000_0000;
array[41983] <= 16'b0000_0000_0000_0000;
array[41984] <= 16'b0000_0000_0000_0000;
array[41985] <= 16'b0000_0000_0000_0000;
array[41986] <= 16'b0000_0000_0000_0000;
array[41987] <= 16'b0000_0000_0000_0000;
array[41988] <= 16'b0000_0000_0000_0000;
array[41989] <= 16'b0000_0000_0000_0000;
array[41990] <= 16'b0000_0000_0000_0000;
array[41991] <= 16'b0000_0000_0000_0000;
array[41992] <= 16'b0000_0000_0000_0000;
array[41993] <= 16'b0000_0000_0000_0000;
array[41994] <= 16'b0000_0000_0000_0000;
array[41995] <= 16'b0000_0000_0000_0000;
array[41996] <= 16'b0000_0000_0000_0000;
array[41997] <= 16'b0000_0000_0000_0000;
array[41998] <= 16'b0000_0000_0000_0000;
array[41999] <= 16'b0000_0000_0000_0000;
array[42000] <= 16'b0000_0000_0000_0000;
array[42001] <= 16'b0000_0000_0000_0000;
array[42002] <= 16'b0000_0000_0000_0000;
array[42003] <= 16'b0000_0000_0000_0000;
array[42004] <= 16'b0000_0000_0000_0000;
array[42005] <= 16'b0000_0000_0000_0000;
array[42006] <= 16'b0000_0000_0000_0000;
array[42007] <= 16'b0000_0000_0000_0000;
array[42008] <= 16'b0000_0000_0000_0000;
array[42009] <= 16'b0000_0000_0000_0000;
array[42010] <= 16'b0000_0000_0000_0000;
array[42011] <= 16'b0000_0000_0000_0000;
array[42012] <= 16'b0000_0000_0000_0000;
array[42013] <= 16'b0000_0000_0000_0000;
array[42014] <= 16'b0000_0000_0000_0000;
array[42015] <= 16'b0000_0000_0000_0000;
array[42016] <= 16'b0000_0000_0000_0000;
array[42017] <= 16'b0000_0000_0000_0000;
array[42018] <= 16'b0000_0000_0000_0000;
array[42019] <= 16'b0000_0000_0000_0000;
array[42020] <= 16'b0000_0000_0000_0000;
array[42021] <= 16'b0000_0000_0000_0000;
array[42022] <= 16'b0000_0000_0000_0000;
array[42023] <= 16'b0000_0000_0000_0000;
array[42024] <= 16'b0000_0000_0000_0000;
array[42025] <= 16'b0000_0000_0000_0000;
array[42026] <= 16'b0000_0000_0000_0000;
array[42027] <= 16'b0000_0000_0000_0000;
array[42028] <= 16'b0000_0000_0000_0000;
array[42029] <= 16'b0000_0000_0000_0000;
array[42030] <= 16'b0000_0000_0000_0000;
array[42031] <= 16'b0000_0000_0000_0000;
array[42032] <= 16'b0000_0000_0000_0000;
array[42033] <= 16'b0000_0000_0000_0000;
array[42034] <= 16'b0000_0000_0000_0000;
array[42035] <= 16'b0000_0000_0000_0000;
array[42036] <= 16'b0000_0000_0000_0000;
array[42037] <= 16'b0000_0000_0000_0000;
array[42038] <= 16'b0000_0000_0000_0000;
array[42039] <= 16'b0000_0000_0000_0000;
array[42040] <= 16'b0000_0000_0000_0000;
array[42041] <= 16'b0000_0000_0000_0000;
array[42042] <= 16'b0000_0000_0000_0000;
array[42043] <= 16'b0000_0000_0000_0000;
array[42044] <= 16'b0000_0000_0000_0000;
array[42045] <= 16'b0000_0000_0000_0000;
array[42046] <= 16'b0000_0000_0000_0000;
array[42047] <= 16'b0000_0000_0000_0000;
array[42048] <= 16'b0000_0000_0000_0000;
array[42049] <= 16'b0000_0000_0000_0000;
array[42050] <= 16'b0000_0000_0000_0000;
array[42051] <= 16'b0000_0000_0000_0000;
array[42052] <= 16'b0000_0000_0000_0000;
array[42053] <= 16'b0000_0000_0000_0000;
array[42054] <= 16'b0000_0000_0000_0000;
array[42055] <= 16'b0000_0000_0000_0000;
array[42056] <= 16'b0000_0000_0000_0000;
array[42057] <= 16'b0000_0000_0000_0000;
array[42058] <= 16'b0000_0000_0000_0000;
array[42059] <= 16'b0000_0000_0000_0000;
array[42060] <= 16'b0000_0000_0000_0000;
array[42061] <= 16'b0000_0000_0000_0000;
array[42062] <= 16'b0000_0000_0000_0000;
array[42063] <= 16'b0000_0000_0000_0000;
array[42064] <= 16'b0000_0000_0000_0000;
array[42065] <= 16'b0000_0000_0000_0000;
array[42066] <= 16'b0000_0000_0000_0000;
array[42067] <= 16'b0000_0000_0000_0000;
array[42068] <= 16'b0000_0000_0000_0000;
array[42069] <= 16'b0000_0000_0000_0000;
array[42070] <= 16'b0000_0000_0000_0000;
array[42071] <= 16'b0000_0000_0000_0000;
array[42072] <= 16'b0000_0000_0000_0000;
array[42073] <= 16'b0000_0000_0000_0000;
array[42074] <= 16'b0000_0000_0000_0000;
array[42075] <= 16'b0000_0000_0000_0000;
array[42076] <= 16'b0000_0000_0000_0000;
array[42077] <= 16'b0000_0000_0000_0000;
array[42078] <= 16'b0000_0000_0000_0000;
array[42079] <= 16'b0000_0000_0000_0000;
array[42080] <= 16'b0000_0000_0000_0000;
array[42081] <= 16'b0000_0000_0000_0000;
array[42082] <= 16'b0000_0000_0000_0000;
array[42083] <= 16'b0000_0000_0000_0000;
array[42084] <= 16'b0000_0000_0000_0000;
array[42085] <= 16'b0000_0000_0000_0000;
array[42086] <= 16'b0000_0000_0000_0000;
array[42087] <= 16'b0000_0000_0000_0000;
array[42088] <= 16'b0000_0000_0000_0000;
array[42089] <= 16'b0000_0000_0000_0000;
array[42090] <= 16'b0000_0000_0000_0000;
array[42091] <= 16'b0000_0000_0000_0000;
array[42092] <= 16'b0000_0000_0000_0000;
array[42093] <= 16'b0000_0000_0000_0000;
array[42094] <= 16'b0000_0000_0000_0000;
array[42095] <= 16'b0000_0000_0000_0000;
array[42096] <= 16'b0000_0000_0000_0000;
array[42097] <= 16'b0000_0000_0000_0000;
array[42098] <= 16'b0000_0000_0000_0000;
array[42099] <= 16'b0000_0000_0000_0000;
array[42100] <= 16'b0000_0000_0000_0000;
array[42101] <= 16'b0000_0000_0000_0000;
array[42102] <= 16'b0000_0000_0000_0000;
array[42103] <= 16'b0000_0000_0000_0000;
array[42104] <= 16'b0000_0000_0000_0000;
array[42105] <= 16'b0000_0000_0000_0000;
array[42106] <= 16'b0000_0000_0000_0000;
array[42107] <= 16'b0000_0000_0000_0000;
array[42108] <= 16'b0000_0000_0000_0000;
array[42109] <= 16'b0000_0000_0000_0000;
array[42110] <= 16'b0000_0000_0000_0000;
array[42111] <= 16'b0000_0000_0000_0000;
array[42112] <= 16'b0000_0000_0000_0000;
array[42113] <= 16'b0000_0000_0000_0000;
array[42114] <= 16'b0000_0000_0000_0000;
array[42115] <= 16'b0000_0000_0000_0000;
array[42116] <= 16'b0000_0000_0000_0000;
array[42117] <= 16'b0000_0000_0000_0000;
array[42118] <= 16'b0000_0000_0000_0000;
array[42119] <= 16'b0000_0000_0000_0000;
array[42120] <= 16'b0000_0000_0000_0000;
array[42121] <= 16'b0000_0000_0000_0000;
array[42122] <= 16'b0000_0000_0000_0000;
array[42123] <= 16'b0000_0000_0000_0000;
array[42124] <= 16'b0000_0000_0000_0000;
array[42125] <= 16'b0000_0000_0000_0000;
array[42126] <= 16'b0000_0000_0000_0000;
array[42127] <= 16'b0000_0000_0000_0000;
array[42128] <= 16'b0000_0000_0000_0000;
array[42129] <= 16'b0000_0000_0000_0000;
array[42130] <= 16'b0000_0000_0000_0000;
array[42131] <= 16'b0000_0000_0000_0000;
array[42132] <= 16'b0000_0000_0000_0000;
array[42133] <= 16'b0000_0000_0000_0000;
array[42134] <= 16'b0000_0000_0000_0000;
array[42135] <= 16'b0000_0000_0000_0000;
array[42136] <= 16'b0000_0000_0000_0000;
array[42137] <= 16'b0000_0000_0000_0000;
array[42138] <= 16'b0000_0000_0000_0000;
array[42139] <= 16'b0000_0000_0000_0000;
array[42140] <= 16'b0000_0000_0000_0000;
array[42141] <= 16'b0000_0000_0000_0000;
array[42142] <= 16'b0000_0000_0000_0000;
array[42143] <= 16'b0000_0000_0000_0000;
array[42144] <= 16'b0000_0000_0000_0000;
array[42145] <= 16'b0000_0000_0000_0000;
array[42146] <= 16'b0000_0000_0000_0000;
array[42147] <= 16'b0000_0000_0000_0000;
array[42148] <= 16'b0000_0000_0000_0000;
array[42149] <= 16'b0000_0000_0000_0000;
array[42150] <= 16'b0000_0000_0000_0000;
array[42151] <= 16'b0000_0000_0000_0000;
array[42152] <= 16'b0000_0000_0000_0000;
array[42153] <= 16'b0000_0000_0000_0000;
array[42154] <= 16'b0000_0000_0000_0000;
array[42155] <= 16'b0000_0000_0000_0000;
array[42156] <= 16'b0000_0000_0000_0000;
array[42157] <= 16'b0000_0000_0000_0000;
array[42158] <= 16'b0000_0000_0000_0000;
array[42159] <= 16'b0000_0000_0000_0000;
array[42160] <= 16'b0000_0000_0000_0000;
array[42161] <= 16'b0000_0000_0000_0000;
array[42162] <= 16'b0000_0000_0000_0000;
array[42163] <= 16'b0000_0000_0000_0000;
array[42164] <= 16'b0000_0000_0000_0000;
array[42165] <= 16'b0000_0000_0000_0000;
array[42166] <= 16'b0000_0000_0000_0000;
array[42167] <= 16'b0000_0000_0000_0000;
array[42168] <= 16'b0000_0000_0000_0000;
array[42169] <= 16'b0000_0000_0000_0000;
array[42170] <= 16'b0000_0000_0000_0000;
array[42171] <= 16'b0000_0000_0000_0000;
array[42172] <= 16'b0000_0000_0000_0000;
array[42173] <= 16'b0000_0000_0000_0000;
array[42174] <= 16'b0000_0000_0000_0000;
array[42175] <= 16'b0000_0000_0000_0000;
array[42176] <= 16'b0000_0000_0000_0000;
array[42177] <= 16'b0000_0000_0000_0000;
array[42178] <= 16'b0000_0000_0000_0000;
array[42179] <= 16'b0000_0000_0000_0000;
array[42180] <= 16'b0000_0000_0000_0000;
array[42181] <= 16'b0000_0000_0000_0000;
array[42182] <= 16'b0000_0000_0000_0000;
array[42183] <= 16'b0000_0000_0000_0000;
array[42184] <= 16'b0000_0000_0000_0000;
array[42185] <= 16'b0000_0000_0000_0000;
array[42186] <= 16'b0000_0000_0000_0000;
array[42187] <= 16'b0000_0000_0000_0000;
array[42188] <= 16'b0000_0000_0000_0000;
array[42189] <= 16'b0000_0000_0000_0000;
array[42190] <= 16'b0000_0000_0000_0000;
array[42191] <= 16'b0000_0000_0000_0000;
array[42192] <= 16'b0000_0000_0000_0000;
array[42193] <= 16'b0000_0000_0000_0000;
array[42194] <= 16'b0000_0000_0000_0000;
array[42195] <= 16'b0000_0000_0000_0000;
array[42196] <= 16'b0000_0000_0000_0000;
array[42197] <= 16'b0000_0000_0000_0000;
array[42198] <= 16'b0000_0000_0000_0000;
array[42199] <= 16'b0000_0000_0000_0000;
array[42200] <= 16'b0000_0000_0000_0000;
array[42201] <= 16'b0000_0000_0000_0000;
array[42202] <= 16'b0000_0000_0000_0000;
array[42203] <= 16'b0000_0000_0000_0000;
array[42204] <= 16'b0000_0000_0000_0000;
array[42205] <= 16'b0000_0000_0000_0000;
array[42206] <= 16'b0000_0000_0000_0000;
array[42207] <= 16'b0000_0000_0000_0000;
array[42208] <= 16'b0000_0000_0000_0000;
array[42209] <= 16'b0000_0000_0000_0000;
array[42210] <= 16'b0000_0000_0000_0000;
array[42211] <= 16'b0000_0000_0000_0000;
array[42212] <= 16'b0000_0000_0000_0000;
array[42213] <= 16'b0000_0000_0000_0000;
array[42214] <= 16'b0000_0000_0000_0000;
array[42215] <= 16'b0000_0000_0000_0000;
array[42216] <= 16'b0000_0000_0000_0000;
array[42217] <= 16'b0000_0000_0000_0000;
array[42218] <= 16'b0000_0000_0000_0000;
array[42219] <= 16'b0000_0000_0000_0000;
array[42220] <= 16'b0000_0000_0000_0000;
array[42221] <= 16'b0000_0000_0000_0000;
array[42222] <= 16'b0000_0000_0000_0000;
array[42223] <= 16'b0000_0000_0000_0000;
array[42224] <= 16'b0000_0000_0000_0000;
array[42225] <= 16'b0000_0000_0000_0000;
array[42226] <= 16'b0000_0000_0000_0000;
array[42227] <= 16'b0000_0000_0000_0000;
array[42228] <= 16'b0000_0000_0000_0000;
array[42229] <= 16'b0000_0000_0000_0000;
array[42230] <= 16'b0000_0000_0000_0000;
array[42231] <= 16'b0000_0000_0000_0000;
array[42232] <= 16'b0000_0000_0000_0000;
array[42233] <= 16'b0000_0000_0000_0000;
array[42234] <= 16'b0000_0000_0000_0000;
array[42235] <= 16'b0000_0000_0000_0000;
array[42236] <= 16'b0000_0000_0000_0000;
array[42237] <= 16'b0000_0000_0000_0000;
array[42238] <= 16'b0000_0000_0000_0000;
array[42239] <= 16'b0000_0000_0000_0000;
array[42240] <= 16'b0000_0000_0000_0000;
array[42241] <= 16'b0000_0000_0000_0000;
array[42242] <= 16'b0000_0000_0000_0000;
array[42243] <= 16'b0000_0000_0000_0000;
array[42244] <= 16'b0000_0000_0000_0000;
array[42245] <= 16'b0000_0000_0000_0000;
array[42246] <= 16'b0000_0000_0000_0000;
array[42247] <= 16'b0000_0000_0000_0000;
array[42248] <= 16'b0000_0000_0000_0000;
array[42249] <= 16'b0000_0000_0000_0000;
array[42250] <= 16'b0000_0000_0000_0000;
array[42251] <= 16'b0000_0000_0000_0000;
array[42252] <= 16'b0000_0000_0000_0000;
array[42253] <= 16'b0000_0000_0000_0000;
array[42254] <= 16'b0000_0000_0000_0000;
array[42255] <= 16'b0000_0000_0000_0000;
array[42256] <= 16'b0000_0000_0000_0000;
array[42257] <= 16'b0000_0000_0000_0000;
array[42258] <= 16'b0000_0000_0000_0000;
array[42259] <= 16'b0000_0000_0000_0000;
array[42260] <= 16'b0000_0000_0000_0000;
array[42261] <= 16'b0000_0000_0000_0000;
array[42262] <= 16'b0000_0000_0000_0000;
array[42263] <= 16'b0000_0000_0000_0000;
array[42264] <= 16'b0000_0000_0000_0000;
array[42265] <= 16'b0000_0000_0000_0000;
array[42266] <= 16'b0000_0000_0000_0000;
array[42267] <= 16'b0000_0000_0000_0000;
array[42268] <= 16'b0000_0000_0000_0000;
array[42269] <= 16'b0000_0000_0000_0000;
array[42270] <= 16'b0000_0000_0000_0000;
array[42271] <= 16'b0000_0000_0000_0000;
array[42272] <= 16'b0000_0000_0000_0000;
array[42273] <= 16'b0000_0000_0000_0000;
array[42274] <= 16'b0000_0000_0000_0000;
array[42275] <= 16'b0000_0000_0000_0000;
array[42276] <= 16'b0000_0000_0000_0000;
array[42277] <= 16'b0000_0000_0000_0000;
array[42278] <= 16'b0000_0000_0000_0000;
array[42279] <= 16'b0000_0000_0000_0000;
array[42280] <= 16'b0000_0000_0000_0000;
array[42281] <= 16'b0000_0000_0000_0000;
array[42282] <= 16'b0000_0000_0000_0000;
array[42283] <= 16'b0000_0000_0000_0000;
array[42284] <= 16'b0000_0000_0000_0000;
array[42285] <= 16'b0000_0000_0000_0000;
array[42286] <= 16'b0000_0000_0000_0000;
array[42287] <= 16'b0000_0000_0000_0000;
array[42288] <= 16'b0000_0000_0000_0000;
array[42289] <= 16'b0000_0000_0000_0000;
array[42290] <= 16'b0000_0000_0000_0000;
array[42291] <= 16'b0000_0000_0000_0000;
array[42292] <= 16'b0000_0000_0000_0000;
array[42293] <= 16'b0000_0000_0000_0000;
array[42294] <= 16'b0000_0000_0000_0000;
array[42295] <= 16'b0000_0000_0000_0000;
array[42296] <= 16'b0000_0000_0000_0000;
array[42297] <= 16'b0000_0000_0000_0000;
array[42298] <= 16'b0000_0000_0000_0000;
array[42299] <= 16'b0000_0000_0000_0000;
array[42300] <= 16'b0000_0000_0000_0000;
array[42301] <= 16'b0000_0000_0000_0000;
array[42302] <= 16'b0000_0000_0000_0000;
array[42303] <= 16'b0000_0000_0000_0000;
array[42304] <= 16'b0000_0000_0000_0000;
array[42305] <= 16'b0000_0000_0000_0000;
array[42306] <= 16'b0000_0000_0000_0000;
array[42307] <= 16'b0000_0000_0000_0000;
array[42308] <= 16'b0000_0000_0000_0000;
array[42309] <= 16'b0000_0000_0000_0000;
array[42310] <= 16'b0000_0000_0000_0000;
array[42311] <= 16'b0000_0000_0000_0000;
array[42312] <= 16'b0000_0000_0000_0000;
array[42313] <= 16'b0000_0000_0000_0000;
array[42314] <= 16'b0000_0000_0000_0000;
array[42315] <= 16'b0000_0000_0000_0000;
array[42316] <= 16'b0000_0000_0000_0000;
array[42317] <= 16'b0000_0000_0000_0000;
array[42318] <= 16'b0000_0000_0000_0000;
array[42319] <= 16'b0000_0000_0000_0000;
array[42320] <= 16'b0000_0000_0000_0000;
array[42321] <= 16'b0000_0000_0000_0000;
array[42322] <= 16'b0000_0000_0000_0000;
array[42323] <= 16'b0000_0000_0000_0000;
array[42324] <= 16'b0000_0000_0000_0000;
array[42325] <= 16'b0000_0000_0000_0000;
array[42326] <= 16'b0000_0000_0000_0000;
array[42327] <= 16'b0000_0000_0000_0000;
array[42328] <= 16'b0000_0000_0000_0000;
array[42329] <= 16'b0000_0000_0000_0000;
array[42330] <= 16'b0000_0000_0000_0000;
array[42331] <= 16'b0000_0000_0000_0000;
array[42332] <= 16'b0000_0000_0000_0000;
array[42333] <= 16'b0000_0000_0000_0000;
array[42334] <= 16'b0000_0000_0000_0000;
array[42335] <= 16'b0000_0000_0000_0000;
array[42336] <= 16'b0000_0000_0000_0000;
array[42337] <= 16'b0000_0000_0000_0000;
array[42338] <= 16'b0000_0000_0000_0000;
array[42339] <= 16'b0000_0000_0000_0000;
array[42340] <= 16'b0000_0000_0000_0000;
array[42341] <= 16'b0000_0000_0000_0000;
array[42342] <= 16'b0000_0000_0000_0000;
array[42343] <= 16'b0000_0000_0000_0000;
array[42344] <= 16'b0000_0000_0000_0000;
array[42345] <= 16'b0000_0000_0000_0000;
array[42346] <= 16'b0000_0000_0000_0000;
array[42347] <= 16'b0000_0000_0000_0000;
array[42348] <= 16'b0000_0000_0000_0000;
array[42349] <= 16'b0000_0000_0000_0000;
array[42350] <= 16'b0000_0000_0000_0000;
array[42351] <= 16'b0000_0000_0000_0000;
array[42352] <= 16'b0000_0000_0000_0000;
array[42353] <= 16'b0000_0000_0000_0000;
array[42354] <= 16'b0000_0000_0000_0000;
array[42355] <= 16'b0000_0000_0000_0000;
array[42356] <= 16'b0000_0000_0000_0000;
array[42357] <= 16'b0000_0000_0000_0000;
array[42358] <= 16'b0000_0000_0000_0000;
array[42359] <= 16'b0000_0000_0000_0000;
array[42360] <= 16'b0000_0000_0000_0000;
array[42361] <= 16'b0000_0000_0000_0000;
array[42362] <= 16'b0000_0000_0000_0000;
array[42363] <= 16'b0000_0000_0000_0000;
array[42364] <= 16'b0000_0000_0000_0000;
array[42365] <= 16'b0000_0000_0000_0000;
array[42366] <= 16'b0000_0000_0000_0000;
array[42367] <= 16'b0000_0000_0000_0000;
array[42368] <= 16'b0000_0000_0000_0000;
array[42369] <= 16'b0000_0000_0000_0000;
array[42370] <= 16'b0000_0000_0000_0000;
array[42371] <= 16'b0000_0000_0000_0000;
array[42372] <= 16'b0000_0000_0000_0000;
array[42373] <= 16'b0000_0000_0000_0000;
array[42374] <= 16'b0000_0000_0000_0000;
array[42375] <= 16'b0000_0000_0000_0000;
array[42376] <= 16'b0000_0000_0000_0000;
array[42377] <= 16'b0000_0000_0000_0000;
array[42378] <= 16'b0000_0000_0000_0000;
array[42379] <= 16'b0000_0000_0000_0000;
array[42380] <= 16'b0000_0000_0000_0000;
array[42381] <= 16'b0000_0000_0000_0000;
array[42382] <= 16'b0000_0000_0000_0000;
array[42383] <= 16'b0000_0000_0000_0000;
array[42384] <= 16'b0000_0000_0000_0000;
array[42385] <= 16'b0000_0000_0000_0000;
array[42386] <= 16'b0000_0000_0000_0000;
array[42387] <= 16'b0000_0000_0000_0000;
array[42388] <= 16'b0000_0000_0000_0000;
array[42389] <= 16'b0000_0000_0000_0000;
array[42390] <= 16'b0000_0000_0000_0000;
array[42391] <= 16'b0000_0000_0000_0000;
array[42392] <= 16'b0000_0000_0000_0000;
array[42393] <= 16'b0000_0000_0000_0000;
array[42394] <= 16'b0000_0000_0000_0000;
array[42395] <= 16'b0000_0000_0000_0000;
array[42396] <= 16'b0000_0000_0000_0000;
array[42397] <= 16'b0000_0000_0000_0000;
array[42398] <= 16'b0000_0000_0000_0000;
array[42399] <= 16'b0000_0000_0000_0000;
array[42400] <= 16'b0000_0000_0000_0000;
array[42401] <= 16'b0000_0000_0000_0000;
array[42402] <= 16'b0000_0000_0000_0000;
array[42403] <= 16'b0000_0000_0000_0000;
array[42404] <= 16'b0000_0000_0000_0000;
array[42405] <= 16'b0000_0000_0000_0000;
array[42406] <= 16'b0000_0000_0000_0000;
array[42407] <= 16'b0000_0000_0000_0000;
array[42408] <= 16'b0000_0000_0000_0000;
array[42409] <= 16'b0000_0000_0000_0000;
array[42410] <= 16'b0000_0000_0000_0000;
array[42411] <= 16'b0000_0000_0000_0000;
array[42412] <= 16'b0000_0000_0000_0000;
array[42413] <= 16'b0000_0000_0000_0000;
array[42414] <= 16'b0000_0000_0000_0000;
array[42415] <= 16'b0000_0000_0000_0000;
array[42416] <= 16'b0000_0000_0000_0000;
array[42417] <= 16'b0000_0000_0000_0000;
array[42418] <= 16'b0000_0000_0000_0000;
array[42419] <= 16'b0000_0000_0000_0000;
array[42420] <= 16'b0000_0000_0000_0000;
array[42421] <= 16'b0000_0000_0000_0000;
array[42422] <= 16'b0000_0000_0000_0000;
array[42423] <= 16'b0000_0000_0000_0000;
array[42424] <= 16'b0000_0000_0000_0000;
array[42425] <= 16'b0000_0000_0000_0000;
array[42426] <= 16'b0000_0000_0000_0000;
array[42427] <= 16'b0000_0000_0000_0000;
array[42428] <= 16'b0000_0000_0000_0000;
array[42429] <= 16'b0000_0000_0000_0000;
array[42430] <= 16'b0000_0000_0000_0000;
array[42431] <= 16'b0000_0000_0000_0000;
array[42432] <= 16'b0000_0000_0000_0000;
array[42433] <= 16'b0000_0000_0000_0000;
array[42434] <= 16'b0000_0000_0000_0000;
array[42435] <= 16'b0000_0000_0000_0000;
array[42436] <= 16'b0000_0000_0000_0000;
array[42437] <= 16'b0000_0000_0000_0000;
array[42438] <= 16'b0000_0000_0000_0000;
array[42439] <= 16'b0000_0000_0000_0000;
array[42440] <= 16'b0000_0000_0000_0000;
array[42441] <= 16'b0000_0000_0000_0000;
array[42442] <= 16'b0000_0000_0000_0000;
array[42443] <= 16'b0000_0000_0000_0000;
array[42444] <= 16'b0000_0000_0000_0000;
array[42445] <= 16'b0000_0000_0000_0000;
array[42446] <= 16'b0000_0000_0000_0000;
array[42447] <= 16'b0000_0000_0000_0000;
array[42448] <= 16'b0000_0000_0000_0000;
array[42449] <= 16'b0000_0000_0000_0000;
array[42450] <= 16'b0000_0000_0000_0000;
array[42451] <= 16'b0000_0000_0000_0000;
array[42452] <= 16'b0000_0000_0000_0000;
array[42453] <= 16'b0000_0000_0000_0000;
array[42454] <= 16'b0000_0000_0000_0000;
array[42455] <= 16'b0000_0000_0000_0000;
array[42456] <= 16'b0000_0000_0000_0000;
array[42457] <= 16'b0000_0000_0000_0000;
array[42458] <= 16'b0000_0000_0000_0000;
array[42459] <= 16'b0000_0000_0000_0000;
array[42460] <= 16'b0000_0000_0000_0000;
array[42461] <= 16'b0000_0000_0000_0000;
array[42462] <= 16'b0000_0000_0000_0000;
array[42463] <= 16'b0000_0000_0000_0000;
array[42464] <= 16'b0000_0000_0000_0000;
array[42465] <= 16'b0000_0000_0000_0000;
array[42466] <= 16'b0000_0000_0000_0000;
array[42467] <= 16'b0000_0000_0000_0000;
array[42468] <= 16'b0000_0000_0000_0000;
array[42469] <= 16'b0000_0000_0000_0000;
array[42470] <= 16'b0000_0000_0000_0000;
array[42471] <= 16'b0000_0000_0000_0000;
array[42472] <= 16'b0000_0000_0000_0000;
array[42473] <= 16'b0000_0000_0000_0000;
array[42474] <= 16'b0000_0000_0000_0000;
array[42475] <= 16'b0000_0000_0000_0000;
array[42476] <= 16'b0000_0000_0000_0000;
array[42477] <= 16'b0000_0000_0000_0000;
array[42478] <= 16'b0000_0000_0000_0000;
array[42479] <= 16'b0000_0000_0000_0000;
array[42480] <= 16'b0000_0000_0000_0000;
array[42481] <= 16'b0000_0000_0000_0000;
array[42482] <= 16'b0000_0000_0000_0000;
array[42483] <= 16'b0000_0000_0000_0000;
array[42484] <= 16'b0000_0000_0000_0000;
array[42485] <= 16'b0000_0000_0000_0000;
array[42486] <= 16'b0000_0000_0000_0000;
array[42487] <= 16'b0000_0000_0000_0000;
array[42488] <= 16'b0000_0000_0000_0000;
array[42489] <= 16'b0000_0000_0000_0000;
array[42490] <= 16'b0000_0000_0000_0000;
array[42491] <= 16'b0000_0000_0000_0000;
array[42492] <= 16'b0000_0000_0000_0000;
array[42493] <= 16'b0000_0000_0000_0000;
array[42494] <= 16'b0000_0000_0000_0000;
array[42495] <= 16'b0000_0000_0000_0000;
array[42496] <= 16'b0000_0000_0000_0000;
array[42497] <= 16'b0000_0000_0000_0000;
array[42498] <= 16'b0000_0000_0000_0000;
array[42499] <= 16'b0000_0000_0000_0000;
array[42500] <= 16'b0000_0000_0000_0000;
array[42501] <= 16'b0000_0000_0000_0000;
array[42502] <= 16'b0000_0000_0000_0000;
array[42503] <= 16'b0000_0000_0000_0000;
array[42504] <= 16'b0000_0000_0000_0000;
array[42505] <= 16'b0000_0000_0000_0000;
array[42506] <= 16'b0000_0000_0000_0000;
array[42507] <= 16'b0000_0000_0000_0000;
array[42508] <= 16'b0000_0000_0000_0000;
array[42509] <= 16'b0000_0000_0000_0000;
array[42510] <= 16'b0000_0000_0000_0000;
array[42511] <= 16'b0000_0000_0000_0000;
array[42512] <= 16'b0000_0000_0000_0000;
array[42513] <= 16'b0000_0000_0000_0000;
array[42514] <= 16'b0000_0000_0000_0000;
array[42515] <= 16'b0000_0000_0000_0000;
array[42516] <= 16'b0000_0000_0000_0000;
array[42517] <= 16'b0000_0000_0000_0000;
array[42518] <= 16'b0000_0000_0000_0000;
array[42519] <= 16'b0000_0000_0000_0000;
array[42520] <= 16'b0000_0000_0000_0000;
array[42521] <= 16'b0000_0000_0000_0000;
array[42522] <= 16'b0000_0000_0000_0000;
array[42523] <= 16'b0000_0000_0000_0000;
array[42524] <= 16'b0000_0000_0000_0000;
array[42525] <= 16'b0000_0000_0000_0000;
array[42526] <= 16'b0000_0000_0000_0000;
array[42527] <= 16'b0000_0000_0000_0000;
array[42528] <= 16'b0000_0000_0000_0000;
array[42529] <= 16'b0000_0000_0000_0000;
array[42530] <= 16'b0000_0000_0000_0000;
array[42531] <= 16'b0000_0000_0000_0000;
array[42532] <= 16'b0000_0000_0000_0000;
array[42533] <= 16'b0000_0000_0000_0000;
array[42534] <= 16'b0000_0000_0000_0000;
array[42535] <= 16'b0000_0000_0000_0000;
array[42536] <= 16'b0000_0000_0000_0000;
array[42537] <= 16'b0000_0000_0000_0000;
array[42538] <= 16'b0000_0000_0000_0000;
array[42539] <= 16'b0000_0000_0000_0000;
array[42540] <= 16'b0000_0000_0000_0000;
array[42541] <= 16'b0000_0000_0000_0000;
array[42542] <= 16'b0000_0000_0000_0000;
array[42543] <= 16'b0000_0000_0000_0000;
array[42544] <= 16'b0000_0000_0000_0000;
array[42545] <= 16'b0000_0000_0000_0000;
array[42546] <= 16'b0000_0000_0000_0000;
array[42547] <= 16'b0000_0000_0000_0000;
array[42548] <= 16'b0000_0000_0000_0000;
array[42549] <= 16'b0000_0000_0000_0000;
array[42550] <= 16'b0000_0000_0000_0000;
array[42551] <= 16'b0000_0000_0000_0000;
array[42552] <= 16'b0000_0000_0000_0000;
array[42553] <= 16'b0000_0000_0000_0000;
array[42554] <= 16'b0000_0000_0000_0000;
array[42555] <= 16'b0000_0000_0000_0000;
array[42556] <= 16'b0000_0000_0000_0000;
array[42557] <= 16'b0000_0000_0000_0000;
array[42558] <= 16'b0000_0000_0000_0000;
array[42559] <= 16'b0000_0000_0000_0000;
array[42560] <= 16'b0000_0000_0000_0000;
array[42561] <= 16'b0000_0000_0000_0000;
array[42562] <= 16'b0000_0000_0000_0000;
array[42563] <= 16'b0000_0000_0000_0000;
array[42564] <= 16'b0000_0000_0000_0000;
array[42565] <= 16'b0000_0000_0000_0000;
array[42566] <= 16'b0000_0000_0000_0000;
array[42567] <= 16'b0000_0000_0000_0000;
array[42568] <= 16'b0000_0000_0000_0000;
array[42569] <= 16'b0000_0000_0000_0000;
array[42570] <= 16'b0000_0000_0000_0000;
array[42571] <= 16'b0000_0000_0000_0000;
array[42572] <= 16'b0000_0000_0000_0000;
array[42573] <= 16'b0000_0000_0000_0000;
array[42574] <= 16'b0000_0000_0000_0000;
array[42575] <= 16'b0000_0000_0000_0000;
array[42576] <= 16'b0000_0000_0000_0000;
array[42577] <= 16'b0000_0000_0000_0000;
array[42578] <= 16'b0000_0000_0000_0000;
array[42579] <= 16'b0000_0000_0000_0000;
array[42580] <= 16'b0000_0000_0000_0000;
array[42581] <= 16'b0000_0000_0000_0000;
array[42582] <= 16'b0000_0000_0000_0000;
array[42583] <= 16'b0000_0000_0000_0000;
array[42584] <= 16'b0000_0000_0000_0000;
array[42585] <= 16'b0000_0000_0000_0000;
array[42586] <= 16'b0000_0000_0000_0000;
array[42587] <= 16'b0000_0000_0000_0000;
array[42588] <= 16'b0000_0000_0000_0000;
array[42589] <= 16'b0000_0000_0000_0000;
array[42590] <= 16'b0000_0000_0000_0000;
array[42591] <= 16'b0000_0000_0000_0000;
array[42592] <= 16'b0000_0000_0000_0000;
array[42593] <= 16'b0000_0000_0000_0000;
array[42594] <= 16'b0000_0000_0000_0000;
array[42595] <= 16'b0000_0000_0000_0000;
array[42596] <= 16'b0000_0000_0000_0000;
array[42597] <= 16'b0000_0000_0000_0000;
array[42598] <= 16'b0000_0000_0000_0000;
array[42599] <= 16'b0000_0000_0000_0000;
array[42600] <= 16'b0000_0000_0000_0000;
array[42601] <= 16'b0000_0000_0000_0000;
array[42602] <= 16'b0000_0000_0000_0000;
array[42603] <= 16'b0000_0000_0000_0000;
array[42604] <= 16'b0000_0000_0000_0000;
array[42605] <= 16'b0000_0000_0000_0000;
array[42606] <= 16'b0000_0000_0000_0000;
array[42607] <= 16'b0000_0000_0000_0000;
array[42608] <= 16'b0000_0000_0000_0000;
array[42609] <= 16'b0000_0000_0000_0000;
array[42610] <= 16'b0000_0000_0000_0000;
array[42611] <= 16'b0000_0000_0000_0000;
array[42612] <= 16'b0000_0000_0000_0000;
array[42613] <= 16'b0000_0000_0000_0000;
array[42614] <= 16'b0000_0000_0000_0000;
array[42615] <= 16'b0000_0000_0000_0000;
array[42616] <= 16'b0000_0000_0000_0000;
array[42617] <= 16'b0000_0000_0000_0000;
array[42618] <= 16'b0000_0000_0000_0000;
array[42619] <= 16'b0000_0000_0000_0000;
array[42620] <= 16'b0000_0000_0000_0000;
array[42621] <= 16'b0000_0000_0000_0000;
array[42622] <= 16'b0000_0000_0000_0000;
array[42623] <= 16'b0000_0000_0000_0000;
array[42624] <= 16'b0000_0000_0000_0000;
array[42625] <= 16'b0000_0000_0000_0000;
array[42626] <= 16'b0000_0000_0000_0000;
array[42627] <= 16'b0000_0000_0000_0000;
array[42628] <= 16'b0000_0000_0000_0000;
array[42629] <= 16'b0000_0000_0000_0000;
array[42630] <= 16'b0000_0000_0000_0000;
array[42631] <= 16'b0000_0000_0000_0000;
array[42632] <= 16'b0000_0000_0000_0000;
array[42633] <= 16'b0000_0000_0000_0000;
array[42634] <= 16'b0000_0000_0000_0000;
array[42635] <= 16'b0000_0000_0000_0000;
array[42636] <= 16'b0000_0000_0000_0000;
array[42637] <= 16'b0000_0000_0000_0000;
array[42638] <= 16'b0000_0000_0000_0000;
array[42639] <= 16'b0000_0000_0000_0000;
array[42640] <= 16'b0000_0000_0000_0000;
array[42641] <= 16'b0000_0000_0000_0000;
array[42642] <= 16'b0000_0000_0000_0000;
array[42643] <= 16'b0000_0000_0000_0000;
array[42644] <= 16'b0000_0000_0000_0000;
array[42645] <= 16'b0000_0000_0000_0000;
array[42646] <= 16'b0000_0000_0000_0000;
array[42647] <= 16'b0000_0000_0000_0000;
array[42648] <= 16'b0000_0000_0000_0000;
array[42649] <= 16'b0000_0000_0000_0000;
array[42650] <= 16'b0000_0000_0000_0000;
array[42651] <= 16'b0000_0000_0000_0000;
array[42652] <= 16'b0000_0000_0000_0000;
array[42653] <= 16'b0000_0000_0000_0000;
array[42654] <= 16'b0000_0000_0000_0000;
array[42655] <= 16'b0000_0000_0000_0000;
array[42656] <= 16'b0000_0000_0000_0000;
array[42657] <= 16'b0000_0000_0000_0000;
array[42658] <= 16'b0000_0000_0000_0000;
array[42659] <= 16'b0000_0000_0000_0000;
array[42660] <= 16'b0000_0000_0000_0000;
array[42661] <= 16'b0000_0000_0000_0000;
array[42662] <= 16'b0000_0000_0000_0000;
array[42663] <= 16'b0000_0000_0000_0000;
array[42664] <= 16'b0000_0000_0000_0000;
array[42665] <= 16'b0000_0000_0000_0000;
array[42666] <= 16'b0000_0000_0000_0000;
array[42667] <= 16'b0000_0000_0000_0000;
array[42668] <= 16'b0000_0000_0000_0000;
array[42669] <= 16'b0000_0000_0000_0000;
array[42670] <= 16'b0000_0000_0000_0000;
array[42671] <= 16'b0000_0000_0000_0000;
array[42672] <= 16'b0000_0000_0000_0000;
array[42673] <= 16'b0000_0000_0000_0000;
array[42674] <= 16'b0000_0000_0000_0000;
array[42675] <= 16'b0000_0000_0000_0000;
array[42676] <= 16'b0000_0000_0000_0000;
array[42677] <= 16'b0000_0000_0000_0000;
array[42678] <= 16'b0000_0000_0000_0000;
array[42679] <= 16'b0000_0000_0000_0000;
array[42680] <= 16'b0000_0000_0000_0000;
array[42681] <= 16'b0000_0000_0000_0000;
array[42682] <= 16'b0000_0000_0000_0000;
array[42683] <= 16'b0000_0000_0000_0000;
array[42684] <= 16'b0000_0000_0000_0000;
array[42685] <= 16'b0000_0000_0000_0000;
array[42686] <= 16'b0000_0000_0000_0000;
array[42687] <= 16'b0000_0000_0000_0000;
array[42688] <= 16'b0000_0000_0000_0000;
array[42689] <= 16'b0000_0000_0000_0000;
array[42690] <= 16'b0000_0000_0000_0000;
array[42691] <= 16'b0000_0000_0000_0000;
array[42692] <= 16'b0000_0000_0000_0000;
array[42693] <= 16'b0000_0000_0000_0000;
array[42694] <= 16'b0000_0000_0000_0000;
array[42695] <= 16'b0000_0000_0000_0000;
array[42696] <= 16'b0000_0000_0000_0000;
array[42697] <= 16'b0000_0000_0000_0000;
array[42698] <= 16'b0000_0000_0000_0000;
array[42699] <= 16'b0000_0000_0000_0000;
array[42700] <= 16'b0000_0000_0000_0000;
array[42701] <= 16'b0000_0000_0000_0000;
array[42702] <= 16'b0000_0000_0000_0000;
array[42703] <= 16'b0000_0000_0000_0000;
array[42704] <= 16'b0000_0000_0000_0000;
array[42705] <= 16'b0000_0000_0000_0000;
array[42706] <= 16'b0000_0000_0000_0000;
array[42707] <= 16'b0000_0000_0000_0000;
array[42708] <= 16'b0000_0000_0000_0000;
array[42709] <= 16'b0000_0000_0000_0000;
array[42710] <= 16'b0000_0000_0000_0000;
array[42711] <= 16'b0000_0000_0000_0000;
array[42712] <= 16'b0000_0000_0000_0000;
array[42713] <= 16'b0000_0000_0000_0000;
array[42714] <= 16'b0000_0000_0000_0000;
array[42715] <= 16'b0000_0000_0000_0000;
array[42716] <= 16'b0000_0000_0000_0000;
array[42717] <= 16'b0000_0000_0000_0000;
array[42718] <= 16'b0000_0000_0000_0000;
array[42719] <= 16'b0000_0000_0000_0000;
array[42720] <= 16'b0000_0000_0000_0000;
array[42721] <= 16'b0000_0000_0000_0000;
array[42722] <= 16'b0000_0000_0000_0000;
array[42723] <= 16'b0000_0000_0000_0000;
array[42724] <= 16'b0000_0000_0000_0000;
array[42725] <= 16'b0000_0000_0000_0000;
array[42726] <= 16'b0000_0000_0000_0000;
array[42727] <= 16'b0000_0000_0000_0000;
array[42728] <= 16'b0000_0000_0000_0000;
array[42729] <= 16'b0000_0000_0000_0000;
array[42730] <= 16'b0000_0000_0000_0000;
array[42731] <= 16'b0000_0000_0000_0000;
array[42732] <= 16'b0000_0000_0000_0000;
array[42733] <= 16'b0000_0000_0000_0000;
array[42734] <= 16'b0000_0000_0000_0000;
array[42735] <= 16'b0000_0000_0000_0000;
array[42736] <= 16'b0000_0000_0000_0000;
array[42737] <= 16'b0000_0000_0000_0000;
array[42738] <= 16'b0000_0000_0000_0000;
array[42739] <= 16'b0000_0000_0000_0000;
array[42740] <= 16'b0000_0000_0000_0000;
array[42741] <= 16'b0000_0000_0000_0000;
array[42742] <= 16'b0000_0000_0000_0000;
array[42743] <= 16'b0000_0000_0000_0000;
array[42744] <= 16'b0000_0000_0000_0000;
array[42745] <= 16'b0000_0000_0000_0000;
array[42746] <= 16'b0000_0000_0000_0000;
array[42747] <= 16'b0000_0000_0000_0000;
array[42748] <= 16'b0000_0000_0000_0000;
array[42749] <= 16'b0000_0000_0000_0000;
array[42750] <= 16'b0000_0000_0000_0000;
array[42751] <= 16'b0000_0000_0000_0000;
array[42752] <= 16'b0000_0000_0000_0000;
array[42753] <= 16'b0000_0000_0000_0000;
array[42754] <= 16'b0000_0000_0000_0000;
array[42755] <= 16'b0000_0000_0000_0000;
array[42756] <= 16'b0000_0000_0000_0000;
array[42757] <= 16'b0000_0000_0000_0000;
array[42758] <= 16'b0000_0000_0000_0000;
array[42759] <= 16'b0000_0000_0000_0000;
array[42760] <= 16'b0000_0000_0000_0000;
array[42761] <= 16'b0000_0000_0000_0000;
array[42762] <= 16'b0000_0000_0000_0000;
array[42763] <= 16'b0000_0000_0000_0000;
array[42764] <= 16'b0000_0000_0000_0000;
array[42765] <= 16'b0000_0000_0000_0000;
array[42766] <= 16'b0000_0000_0000_0000;
array[42767] <= 16'b0000_0000_0000_0000;
array[42768] <= 16'b0000_0000_0000_0000;
array[42769] <= 16'b0000_0000_0000_0000;
array[42770] <= 16'b0000_0000_0000_0000;
array[42771] <= 16'b0000_0000_0000_0000;
array[42772] <= 16'b0000_0000_0000_0000;
array[42773] <= 16'b0000_0000_0000_0000;
array[42774] <= 16'b0000_0000_0000_0000;
array[42775] <= 16'b0000_0000_0000_0000;
array[42776] <= 16'b0000_0000_0000_0000;
array[42777] <= 16'b0000_0000_0000_0000;
array[42778] <= 16'b0000_0000_0000_0000;
array[42779] <= 16'b0000_0000_0000_0000;
array[42780] <= 16'b0000_0000_0000_0000;
array[42781] <= 16'b0000_0000_0000_0000;
array[42782] <= 16'b0000_0000_0000_0000;
array[42783] <= 16'b0000_0000_0000_0000;
array[42784] <= 16'b0000_0000_0000_0000;
array[42785] <= 16'b0000_0000_0000_0000;
array[42786] <= 16'b0000_0000_0000_0000;
array[42787] <= 16'b0000_0000_0000_0000;
array[42788] <= 16'b0000_0000_0000_0000;
array[42789] <= 16'b0000_0000_0000_0000;
array[42790] <= 16'b0000_0000_0000_0000;
array[42791] <= 16'b0000_0000_0000_0000;
array[42792] <= 16'b0000_0000_0000_0000;
array[42793] <= 16'b0000_0000_0000_0000;
array[42794] <= 16'b0000_0000_0000_0000;
array[42795] <= 16'b0000_0000_0000_0000;
array[42796] <= 16'b0000_0000_0000_0000;
array[42797] <= 16'b0000_0000_0000_0000;
array[42798] <= 16'b0000_0000_0000_0000;
array[42799] <= 16'b0000_0000_0000_0000;
array[42800] <= 16'b0000_0000_0000_0000;
array[42801] <= 16'b0000_0000_0000_0000;
array[42802] <= 16'b0000_0000_0000_0000;
array[42803] <= 16'b0000_0000_0000_0000;
array[42804] <= 16'b0000_0000_0000_0000;
array[42805] <= 16'b0000_0000_0000_0000;
array[42806] <= 16'b0000_0000_0000_0000;
array[42807] <= 16'b0000_0000_0000_0000;
array[42808] <= 16'b0000_0000_0000_0000;
array[42809] <= 16'b0000_0000_0000_0000;
array[42810] <= 16'b0000_0000_0000_0000;
array[42811] <= 16'b0000_0000_0000_0000;
array[42812] <= 16'b0000_0000_0000_0000;
array[42813] <= 16'b0000_0000_0000_0000;
array[42814] <= 16'b0000_0000_0000_0000;
array[42815] <= 16'b0000_0000_0000_0000;
array[42816] <= 16'b0000_0000_0000_0000;
array[42817] <= 16'b0000_0000_0000_0000;
array[42818] <= 16'b0000_0000_0000_0000;
array[42819] <= 16'b0000_0000_0000_0000;
array[42820] <= 16'b0000_0000_0000_0000;
array[42821] <= 16'b0000_0000_0000_0000;
array[42822] <= 16'b0000_0000_0000_0000;
array[42823] <= 16'b0000_0000_0000_0000;
array[42824] <= 16'b0000_0000_0000_0000;
array[42825] <= 16'b0000_0000_0000_0000;
array[42826] <= 16'b0000_0000_0000_0000;
array[42827] <= 16'b0000_0000_0000_0000;
array[42828] <= 16'b0000_0000_0000_0000;
array[42829] <= 16'b0000_0000_0000_0000;
array[42830] <= 16'b0000_0000_0000_0000;
array[42831] <= 16'b0000_0000_0000_0000;
array[42832] <= 16'b0000_0000_0000_0000;
array[42833] <= 16'b0000_0000_0000_0000;
array[42834] <= 16'b0000_0000_0000_0000;
array[42835] <= 16'b0000_0000_0000_0000;
array[42836] <= 16'b0000_0000_0000_0000;
array[42837] <= 16'b0000_0000_0000_0000;
array[42838] <= 16'b0000_0000_0000_0000;
array[42839] <= 16'b0000_0000_0000_0000;
array[42840] <= 16'b0000_0000_0000_0000;
array[42841] <= 16'b0000_0000_0000_0000;
array[42842] <= 16'b0000_0000_0000_0000;
array[42843] <= 16'b0000_0000_0000_0000;
array[42844] <= 16'b0000_0000_0000_0000;
array[42845] <= 16'b0000_0000_0000_0000;
array[42846] <= 16'b0000_0000_0000_0000;
array[42847] <= 16'b0000_0000_0000_0000;
array[42848] <= 16'b0000_0000_0000_0000;
array[42849] <= 16'b0000_0000_0000_0000;
array[42850] <= 16'b0000_0000_0000_0000;
array[42851] <= 16'b0000_0000_0000_0000;
array[42852] <= 16'b0000_0000_0000_0000;
array[42853] <= 16'b0000_0000_0000_0000;
array[42854] <= 16'b0000_0000_0000_0000;
array[42855] <= 16'b0000_0000_0000_0000;
array[42856] <= 16'b0000_0000_0000_0000;
array[42857] <= 16'b0000_0000_0000_0000;
array[42858] <= 16'b0000_0000_0000_0000;
array[42859] <= 16'b0000_0000_0000_0000;
array[42860] <= 16'b0000_0000_0000_0000;
array[42861] <= 16'b0000_0000_0000_0000;
array[42862] <= 16'b0000_0000_0000_0000;
array[42863] <= 16'b0000_0000_0000_0000;
array[42864] <= 16'b0000_0000_0000_0000;
array[42865] <= 16'b0000_0000_0000_0000;
array[42866] <= 16'b0000_0000_0000_0000;
array[42867] <= 16'b0000_0000_0000_0000;
array[42868] <= 16'b0000_0000_0000_0000;
array[42869] <= 16'b0000_0000_0000_0000;
array[42870] <= 16'b0000_0000_0000_0000;
array[42871] <= 16'b0000_0000_0000_0000;
array[42872] <= 16'b0000_0000_0000_0000;
array[42873] <= 16'b0000_0000_0000_0000;
array[42874] <= 16'b0000_0000_0000_0000;
array[42875] <= 16'b0000_0000_0000_0000;
array[42876] <= 16'b0000_0000_0000_0000;
array[42877] <= 16'b0000_0000_0000_0000;
array[42878] <= 16'b0000_0000_0000_0000;
array[42879] <= 16'b0000_0000_0000_0000;
array[42880] <= 16'b0000_0000_0000_0000;
array[42881] <= 16'b0000_0000_0000_0000;
array[42882] <= 16'b0000_0000_0000_0000;
array[42883] <= 16'b0000_0000_0000_0000;
array[42884] <= 16'b0000_0000_0000_0000;
array[42885] <= 16'b0000_0000_0000_0000;
array[42886] <= 16'b0000_0000_0000_0000;
array[42887] <= 16'b0000_0000_0000_0000;
array[42888] <= 16'b0000_0000_0000_0000;
array[42889] <= 16'b0000_0000_0000_0000;
array[42890] <= 16'b0000_0000_0000_0000;
array[42891] <= 16'b0000_0000_0000_0000;
array[42892] <= 16'b0000_0000_0000_0000;
array[42893] <= 16'b0000_0000_0000_0000;
array[42894] <= 16'b0000_0000_0000_0000;
array[42895] <= 16'b0000_0000_0000_0000;
array[42896] <= 16'b0000_0000_0000_0000;
array[42897] <= 16'b0000_0000_0000_0000;
array[42898] <= 16'b0000_0000_0000_0000;
array[42899] <= 16'b0000_0000_0000_0000;
array[42900] <= 16'b0000_0000_0000_0000;
array[42901] <= 16'b0000_0000_0000_0000;
array[42902] <= 16'b0000_0000_0000_0000;
array[42903] <= 16'b0000_0000_0000_0000;
array[42904] <= 16'b0000_0000_0000_0000;
array[42905] <= 16'b0000_0000_0000_0000;
array[42906] <= 16'b0000_0000_0000_0000;
array[42907] <= 16'b0000_0000_0000_0000;
array[42908] <= 16'b0000_0000_0000_0000;
array[42909] <= 16'b0000_0000_0000_0000;
array[42910] <= 16'b0000_0000_0000_0000;
array[42911] <= 16'b0000_0000_0000_0000;
array[42912] <= 16'b0000_0000_0000_0000;
array[42913] <= 16'b0000_0000_0000_0000;
array[42914] <= 16'b0000_0000_0000_0000;
array[42915] <= 16'b0000_0000_0000_0000;
array[42916] <= 16'b0000_0000_0000_0000;
array[42917] <= 16'b0000_0000_0000_0000;
array[42918] <= 16'b0000_0000_0000_0000;
array[42919] <= 16'b0000_0000_0000_0000;
array[42920] <= 16'b0000_0000_0000_0000;
array[42921] <= 16'b0000_0000_0000_0000;
array[42922] <= 16'b0000_0000_0000_0000;
array[42923] <= 16'b0000_0000_0000_0000;
array[42924] <= 16'b0000_0000_0000_0000;
array[42925] <= 16'b0000_0000_0000_0000;
array[42926] <= 16'b0000_0000_0000_0000;
array[42927] <= 16'b0000_0000_0000_0000;
array[42928] <= 16'b0000_0000_0000_0000;
array[42929] <= 16'b0000_0000_0000_0000;
array[42930] <= 16'b0000_0000_0000_0000;
array[42931] <= 16'b0000_0000_0000_0000;
array[42932] <= 16'b0000_0000_0000_0000;
array[42933] <= 16'b0000_0000_0000_0000;
array[42934] <= 16'b0000_0000_0000_0000;
array[42935] <= 16'b0000_0000_0000_0000;
array[42936] <= 16'b0000_0000_0000_0000;
array[42937] <= 16'b0000_0000_0000_0000;
array[42938] <= 16'b0000_0000_0000_0000;
array[42939] <= 16'b0000_0000_0000_0000;
array[42940] <= 16'b0000_0000_0000_0000;
array[42941] <= 16'b0000_0000_0000_0000;
array[42942] <= 16'b0000_0000_0000_0000;
array[42943] <= 16'b0000_0000_0000_0000;
array[42944] <= 16'b0000_0000_0000_0000;
array[42945] <= 16'b0000_0000_0000_0000;
array[42946] <= 16'b0000_0000_0000_0000;
array[42947] <= 16'b0000_0000_0000_0000;
array[42948] <= 16'b0000_0000_0000_0000;
array[42949] <= 16'b0000_0000_0000_0000;
array[42950] <= 16'b0000_0000_0000_0000;
array[42951] <= 16'b0000_0000_0000_0000;
array[42952] <= 16'b0000_0000_0000_0000;
array[42953] <= 16'b0000_0000_0000_0000;
array[42954] <= 16'b0000_0000_0000_0000;
array[42955] <= 16'b0000_0000_0000_0000;
array[42956] <= 16'b0000_0000_0000_0000;
array[42957] <= 16'b0000_0000_0000_0000;
array[42958] <= 16'b0000_0000_0000_0000;
array[42959] <= 16'b0000_0000_0000_0000;
array[42960] <= 16'b0000_0000_0000_0000;
array[42961] <= 16'b0000_0000_0000_0000;
array[42962] <= 16'b0000_0000_0000_0000;
array[42963] <= 16'b0000_0000_0000_0000;
array[42964] <= 16'b0000_0000_0000_0000;
array[42965] <= 16'b0000_0000_0000_0000;
array[42966] <= 16'b0000_0000_0000_0000;
array[42967] <= 16'b0000_0000_0000_0000;
array[42968] <= 16'b0000_0000_0000_0000;
array[42969] <= 16'b0000_0000_0000_0000;
array[42970] <= 16'b0000_0000_0000_0000;
array[42971] <= 16'b0000_0000_0000_0000;
array[42972] <= 16'b0000_0000_0000_0000;
array[42973] <= 16'b0000_0000_0000_0000;
array[42974] <= 16'b0000_0000_0000_0000;
array[42975] <= 16'b0000_0000_0000_0000;
array[42976] <= 16'b0000_0000_0000_0000;
array[42977] <= 16'b0000_0000_0000_0000;
array[42978] <= 16'b0000_0000_0000_0000;
array[42979] <= 16'b0000_0000_0000_0000;
array[42980] <= 16'b0000_0000_0000_0000;
array[42981] <= 16'b0000_0000_0000_0000;
array[42982] <= 16'b0000_0000_0000_0000;
array[42983] <= 16'b0000_0000_0000_0000;
array[42984] <= 16'b0000_0000_0000_0000;
array[42985] <= 16'b0000_0000_0000_0000;
array[42986] <= 16'b0000_0000_0000_0000;
array[42987] <= 16'b0000_0000_0000_0000;
array[42988] <= 16'b0000_0000_0000_0000;
array[42989] <= 16'b0000_0000_0000_0000;
array[42990] <= 16'b0000_0000_0000_0000;
array[42991] <= 16'b0000_0000_0000_0000;
array[42992] <= 16'b0000_0000_0000_0000;
array[42993] <= 16'b0000_0000_0000_0000;
array[42994] <= 16'b0000_0000_0000_0000;
array[42995] <= 16'b0000_0000_0000_0000;
array[42996] <= 16'b0000_0000_0000_0000;
array[42997] <= 16'b0000_0000_0000_0000;
array[42998] <= 16'b0000_0000_0000_0000;
array[42999] <= 16'b0000_0000_0000_0000;
array[43000] <= 16'b0000_0000_0000_0000;
array[43001] <= 16'b0000_0000_0000_0000;
array[43002] <= 16'b0000_0000_0000_0000;
array[43003] <= 16'b0000_0000_0000_0000;
array[43004] <= 16'b0000_0000_0000_0000;
array[43005] <= 16'b0000_0000_0000_0000;
array[43006] <= 16'b0000_0000_0000_0000;
array[43007] <= 16'b0000_0000_0000_0000;
array[43008] <= 16'b0000_0000_0000_0000;
array[43009] <= 16'b0000_0000_0000_0000;
array[43010] <= 16'b0000_0000_0000_0000;
array[43011] <= 16'b0000_0000_0000_0000;
array[43012] <= 16'b0000_0000_0000_0000;
array[43013] <= 16'b0000_0000_0000_0000;
array[43014] <= 16'b0000_0000_0000_0000;
array[43015] <= 16'b0000_0000_0000_0000;
array[43016] <= 16'b0000_0000_0000_0000;
array[43017] <= 16'b0000_0000_0000_0000;
array[43018] <= 16'b0000_0000_0000_0000;
array[43019] <= 16'b0000_0000_0000_0000;
array[43020] <= 16'b0000_0000_0000_0000;
array[43021] <= 16'b0000_0000_0000_0000;
array[43022] <= 16'b0000_0000_0000_0000;
array[43023] <= 16'b0000_0000_0000_0000;
array[43024] <= 16'b0000_0000_0000_0000;
array[43025] <= 16'b0000_0000_0000_0000;
array[43026] <= 16'b0000_0000_0000_0000;
array[43027] <= 16'b0000_0000_0000_0000;
array[43028] <= 16'b0000_0000_0000_0000;
array[43029] <= 16'b0000_0000_0000_0000;
array[43030] <= 16'b0000_0000_0000_0000;
array[43031] <= 16'b0000_0000_0000_0000;
array[43032] <= 16'b0000_0000_0000_0000;
array[43033] <= 16'b0000_0000_0000_0000;
array[43034] <= 16'b0000_0000_0000_0000;
array[43035] <= 16'b0000_0000_0000_0000;
array[43036] <= 16'b0000_0000_0000_0000;
array[43037] <= 16'b0000_0000_0000_0000;
array[43038] <= 16'b0000_0000_0000_0000;
array[43039] <= 16'b0000_0000_0000_0000;
array[43040] <= 16'b0000_0000_0000_0000;
array[43041] <= 16'b0000_0000_0000_0000;
array[43042] <= 16'b0000_0000_0000_0000;
array[43043] <= 16'b0000_0000_0000_0000;
array[43044] <= 16'b0000_0000_0000_0000;
array[43045] <= 16'b0000_0000_0000_0000;
array[43046] <= 16'b0000_0000_0000_0000;
array[43047] <= 16'b0000_0000_0000_0000;
array[43048] <= 16'b0000_0000_0000_0000;
array[43049] <= 16'b0000_0000_0000_0000;
array[43050] <= 16'b0000_0000_0000_0000;
array[43051] <= 16'b0000_0000_0000_0000;
array[43052] <= 16'b0000_0000_0000_0000;
array[43053] <= 16'b0000_0000_0000_0000;
array[43054] <= 16'b0000_0000_0000_0000;
array[43055] <= 16'b0000_0000_0000_0000;
array[43056] <= 16'b0000_0000_0000_0000;
array[43057] <= 16'b0000_0000_0000_0000;
array[43058] <= 16'b0000_0000_0000_0000;
array[43059] <= 16'b0000_0000_0000_0000;
array[43060] <= 16'b0000_0000_0000_0000;
array[43061] <= 16'b0000_0000_0000_0000;
array[43062] <= 16'b0000_0000_0000_0000;
array[43063] <= 16'b0000_0000_0000_0000;
array[43064] <= 16'b0000_0000_0000_0000;
array[43065] <= 16'b0000_0000_0000_0000;
array[43066] <= 16'b0000_0000_0000_0000;
array[43067] <= 16'b0000_0000_0000_0000;
array[43068] <= 16'b0000_0000_0000_0000;
array[43069] <= 16'b0000_0000_0000_0000;
array[43070] <= 16'b0000_0000_0000_0000;
array[43071] <= 16'b0000_0000_0000_0000;
array[43072] <= 16'b0000_0000_0000_0000;
array[43073] <= 16'b0000_0000_0000_0000;
array[43074] <= 16'b0000_0000_0000_0000;
array[43075] <= 16'b0000_0000_0000_0000;
array[43076] <= 16'b0000_0000_0000_0000;
array[43077] <= 16'b0000_0000_0000_0000;
array[43078] <= 16'b0000_0000_0000_0000;
array[43079] <= 16'b0000_0000_0000_0000;
array[43080] <= 16'b0000_0000_0000_0000;
array[43081] <= 16'b0000_0000_0000_0000;
array[43082] <= 16'b0000_0000_0000_0000;
array[43083] <= 16'b0000_0000_0000_0000;
array[43084] <= 16'b0000_0000_0000_0000;
array[43085] <= 16'b0000_0000_0000_0000;
array[43086] <= 16'b0000_0000_0000_0000;
array[43087] <= 16'b0000_0000_0000_0000;
array[43088] <= 16'b0000_0000_0000_0000;
array[43089] <= 16'b0000_0000_0000_0000;
array[43090] <= 16'b0000_0000_0000_0000;
array[43091] <= 16'b0000_0000_0000_0000;
array[43092] <= 16'b0000_0000_0000_0000;
array[43093] <= 16'b0000_0000_0000_0000;
array[43094] <= 16'b0000_0000_0000_0000;
array[43095] <= 16'b0000_0000_0000_0000;
array[43096] <= 16'b0000_0000_0000_0000;
array[43097] <= 16'b0000_0000_0000_0000;
array[43098] <= 16'b0000_0000_0000_0000;
array[43099] <= 16'b0000_0000_0000_0000;
array[43100] <= 16'b0000_0000_0000_0000;
array[43101] <= 16'b0000_0000_0000_0000;
array[43102] <= 16'b0000_0000_0000_0000;
array[43103] <= 16'b0000_0000_0000_0000;
array[43104] <= 16'b0000_0000_0000_0000;
array[43105] <= 16'b0000_0000_0000_0000;
array[43106] <= 16'b0000_0000_0000_0000;
array[43107] <= 16'b0000_0000_0000_0000;
array[43108] <= 16'b0000_0000_0000_0000;
array[43109] <= 16'b0000_0000_0000_0000;
array[43110] <= 16'b0000_0000_0000_0000;
array[43111] <= 16'b0000_0000_0000_0000;
array[43112] <= 16'b0000_0000_0000_0000;
array[43113] <= 16'b0000_0000_0000_0000;
array[43114] <= 16'b0000_0000_0000_0000;
array[43115] <= 16'b0000_0000_0000_0000;
array[43116] <= 16'b0000_0000_0000_0000;
array[43117] <= 16'b0000_0000_0000_0000;
array[43118] <= 16'b0000_0000_0000_0000;
array[43119] <= 16'b0000_0000_0000_0000;
array[43120] <= 16'b0000_0000_0000_0000;
array[43121] <= 16'b0000_0000_0000_0000;
array[43122] <= 16'b0000_0000_0000_0000;
array[43123] <= 16'b0000_0000_0000_0000;
array[43124] <= 16'b0000_0000_0000_0000;
array[43125] <= 16'b0000_0000_0000_0000;
array[43126] <= 16'b0000_0000_0000_0000;
array[43127] <= 16'b0000_0000_0000_0000;
array[43128] <= 16'b0000_0000_0000_0000;
array[43129] <= 16'b0000_0000_0000_0000;
array[43130] <= 16'b0000_0000_0000_0000;
array[43131] <= 16'b0000_0000_0000_0000;
array[43132] <= 16'b0000_0000_0000_0000;
array[43133] <= 16'b0000_0000_0000_0000;
array[43134] <= 16'b0000_0000_0000_0000;
array[43135] <= 16'b0000_0000_0000_0000;
array[43136] <= 16'b0000_0000_0000_0000;
array[43137] <= 16'b0000_0000_0000_0000;
array[43138] <= 16'b0000_0000_0000_0000;
array[43139] <= 16'b0000_0000_0000_0000;
array[43140] <= 16'b0000_0000_0000_0000;
array[43141] <= 16'b0000_0000_0000_0000;
array[43142] <= 16'b0000_0000_0000_0000;
array[43143] <= 16'b0000_0000_0000_0000;
array[43144] <= 16'b0000_0000_0000_0000;
array[43145] <= 16'b0000_0000_0000_0000;
array[43146] <= 16'b0000_0000_0000_0000;
array[43147] <= 16'b0000_0000_0000_0000;
array[43148] <= 16'b0000_0000_0000_0000;
array[43149] <= 16'b0000_0000_0000_0000;
array[43150] <= 16'b0000_0000_0000_0000;
array[43151] <= 16'b0000_0000_0000_0000;
array[43152] <= 16'b0000_0000_0000_0000;
array[43153] <= 16'b0000_0000_0000_0000;
array[43154] <= 16'b0000_0000_0000_0000;
array[43155] <= 16'b0000_0000_0000_0000;
array[43156] <= 16'b0000_0000_0000_0000;
array[43157] <= 16'b0000_0000_0000_0000;
array[43158] <= 16'b0000_0000_0000_0000;
array[43159] <= 16'b0000_0000_0000_0000;
array[43160] <= 16'b0000_0000_0000_0000;
array[43161] <= 16'b0000_0000_0000_0000;
array[43162] <= 16'b0000_0000_0000_0000;
array[43163] <= 16'b0000_0000_0000_0000;
array[43164] <= 16'b0000_0000_0000_0000;
array[43165] <= 16'b0000_0000_0000_0000;
array[43166] <= 16'b0000_0000_0000_0000;
array[43167] <= 16'b0000_0000_0000_0000;
array[43168] <= 16'b0000_0000_0000_0000;
array[43169] <= 16'b0000_0000_0000_0000;
array[43170] <= 16'b0000_0000_0000_0000;
array[43171] <= 16'b0000_0000_0000_0000;
array[43172] <= 16'b0000_0000_0000_0000;
array[43173] <= 16'b0000_0000_0000_0000;
array[43174] <= 16'b0000_0000_0000_0000;
array[43175] <= 16'b0000_0000_0000_0000;
array[43176] <= 16'b0000_0000_0000_0000;
array[43177] <= 16'b0000_0000_0000_0000;
array[43178] <= 16'b0000_0000_0000_0000;
array[43179] <= 16'b0000_0000_0000_0000;
array[43180] <= 16'b0000_0000_0000_0000;
array[43181] <= 16'b0000_0000_0000_0000;
array[43182] <= 16'b0000_0000_0000_0000;
array[43183] <= 16'b0000_0000_0000_0000;
array[43184] <= 16'b0000_0000_0000_0000;
array[43185] <= 16'b0000_0000_0000_0000;
array[43186] <= 16'b0000_0000_0000_0000;
array[43187] <= 16'b0000_0000_0000_0000;
array[43188] <= 16'b0000_0000_0000_0000;
array[43189] <= 16'b0000_0000_0000_0000;
array[43190] <= 16'b0000_0000_0000_0000;
array[43191] <= 16'b0000_0000_0000_0000;
array[43192] <= 16'b0000_0000_0000_0000;
array[43193] <= 16'b0000_0000_0000_0000;
array[43194] <= 16'b0000_0000_0000_0000;
array[43195] <= 16'b0000_0000_0000_0000;
array[43196] <= 16'b0000_0000_0000_0000;
array[43197] <= 16'b0000_0000_0000_0000;
array[43198] <= 16'b0000_0000_0000_0000;
array[43199] <= 16'b0000_0000_0000_0000;
array[43200] <= 16'b0000_0000_0000_0000;
array[43201] <= 16'b0000_0000_0000_0000;
array[43202] <= 16'b0000_0000_0000_0000;
array[43203] <= 16'b0000_0000_0000_0000;
array[43204] <= 16'b0000_0000_0000_0000;
array[43205] <= 16'b0000_0000_0000_0000;
array[43206] <= 16'b0000_0000_0000_0000;
array[43207] <= 16'b0000_0000_0000_0000;
array[43208] <= 16'b0000_0000_0000_0000;
array[43209] <= 16'b0000_0000_0000_0000;
array[43210] <= 16'b0000_0000_0000_0000;
array[43211] <= 16'b0000_0000_0000_0000;
array[43212] <= 16'b0000_0000_0000_0000;
array[43213] <= 16'b0000_0000_0000_0000;
array[43214] <= 16'b0000_0000_0000_0000;
array[43215] <= 16'b0000_0000_0000_0000;
array[43216] <= 16'b0000_0000_0000_0000;
array[43217] <= 16'b0000_0000_0000_0000;
array[43218] <= 16'b0000_0000_0000_0000;
array[43219] <= 16'b0000_0000_0000_0000;
array[43220] <= 16'b0000_0000_0000_0000;
array[43221] <= 16'b0000_0000_0000_0000;
array[43222] <= 16'b0000_0000_0000_0000;
array[43223] <= 16'b0000_0000_0000_0000;
array[43224] <= 16'b0000_0000_0000_0000;
array[43225] <= 16'b0000_0000_0000_0000;
array[43226] <= 16'b0000_0000_0000_0000;
array[43227] <= 16'b0000_0000_0000_0000;
array[43228] <= 16'b0000_0000_0000_0000;
array[43229] <= 16'b0000_0000_0000_0000;
array[43230] <= 16'b0000_0000_0000_0000;
array[43231] <= 16'b0000_0000_0000_0000;
array[43232] <= 16'b0000_0000_0000_0000;
array[43233] <= 16'b0000_0000_0000_0000;
array[43234] <= 16'b0000_0000_0000_0000;
array[43235] <= 16'b0000_0000_0000_0000;
array[43236] <= 16'b0000_0000_0000_0000;
array[43237] <= 16'b0000_0000_0000_0000;
array[43238] <= 16'b0000_0000_0000_0000;
array[43239] <= 16'b0000_0000_0000_0000;
array[43240] <= 16'b0000_0000_0000_0000;
array[43241] <= 16'b0000_0000_0000_0000;
array[43242] <= 16'b0000_0000_0000_0000;
array[43243] <= 16'b0000_0000_0000_0000;
array[43244] <= 16'b0000_0000_0000_0000;
array[43245] <= 16'b0000_0000_0000_0000;
array[43246] <= 16'b0000_0000_0000_0000;
array[43247] <= 16'b0000_0000_0000_0000;
array[43248] <= 16'b0000_0000_0000_0000;
array[43249] <= 16'b0000_0000_0000_0000;
array[43250] <= 16'b0000_0000_0000_0000;
array[43251] <= 16'b0000_0000_0000_0000;
array[43252] <= 16'b0000_0000_0000_0000;
array[43253] <= 16'b0000_0000_0000_0000;
array[43254] <= 16'b0000_0000_0000_0000;
array[43255] <= 16'b0000_0000_0000_0000;
array[43256] <= 16'b0000_0000_0000_0000;
array[43257] <= 16'b0000_0000_0000_0000;
array[43258] <= 16'b0000_0000_0000_0000;
array[43259] <= 16'b0000_0000_0000_0000;
array[43260] <= 16'b0000_0000_0000_0000;
array[43261] <= 16'b0000_0000_0000_0000;
array[43262] <= 16'b0000_0000_0000_0000;
array[43263] <= 16'b0000_0000_0000_0000;
array[43264] <= 16'b0000_0000_0000_0000;
array[43265] <= 16'b0000_0000_0000_0000;
array[43266] <= 16'b0000_0000_0000_0000;
array[43267] <= 16'b0000_0000_0000_0000;
array[43268] <= 16'b0000_0000_0000_0000;
array[43269] <= 16'b0000_0000_0000_0000;
array[43270] <= 16'b0000_0000_0000_0000;
array[43271] <= 16'b0000_0000_0000_0000;
array[43272] <= 16'b0000_0000_0000_0000;
array[43273] <= 16'b0000_0000_0000_0000;
array[43274] <= 16'b0000_0000_0000_0000;
array[43275] <= 16'b0000_0000_0000_0000;
array[43276] <= 16'b0000_0000_0000_0000;
array[43277] <= 16'b0000_0000_0000_0000;
array[43278] <= 16'b0000_0000_0000_0000;
array[43279] <= 16'b0000_0000_0000_0000;
array[43280] <= 16'b0000_0000_0000_0000;
array[43281] <= 16'b0000_0000_0000_0000;
array[43282] <= 16'b0000_0000_0000_0000;
array[43283] <= 16'b0000_0000_0000_0000;
array[43284] <= 16'b0000_0000_0000_0000;
array[43285] <= 16'b0000_0000_0000_0000;
array[43286] <= 16'b0000_0000_0000_0000;
array[43287] <= 16'b0000_0000_0000_0000;
array[43288] <= 16'b0000_0000_0000_0000;
array[43289] <= 16'b0000_0000_0000_0000;
array[43290] <= 16'b0000_0000_0000_0000;
array[43291] <= 16'b0000_0000_0000_0000;
array[43292] <= 16'b0000_0000_0000_0000;
array[43293] <= 16'b0000_0000_0000_0000;
array[43294] <= 16'b0000_0000_0000_0000;
array[43295] <= 16'b0000_0000_0000_0000;
array[43296] <= 16'b0000_0000_0000_0000;
array[43297] <= 16'b0000_0000_0000_0000;
array[43298] <= 16'b0000_0000_0000_0000;
array[43299] <= 16'b0000_0000_0000_0000;
array[43300] <= 16'b0000_0000_0000_0000;
array[43301] <= 16'b0000_0000_0000_0000;
array[43302] <= 16'b0000_0000_0000_0000;
array[43303] <= 16'b0000_0000_0000_0000;
array[43304] <= 16'b0000_0000_0000_0000;
array[43305] <= 16'b0000_0000_0000_0000;
array[43306] <= 16'b0000_0000_0000_0000;
array[43307] <= 16'b0000_0000_0000_0000;
array[43308] <= 16'b0000_0000_0000_0000;
array[43309] <= 16'b0000_0000_0000_0000;
array[43310] <= 16'b0000_0000_0000_0000;
array[43311] <= 16'b0000_0000_0000_0000;
array[43312] <= 16'b0000_0000_0000_0000;
array[43313] <= 16'b0000_0000_0000_0000;
array[43314] <= 16'b0000_0000_0000_0000;
array[43315] <= 16'b0000_0000_0000_0000;
array[43316] <= 16'b0000_0000_0000_0000;
array[43317] <= 16'b0000_0000_0000_0000;
array[43318] <= 16'b0000_0000_0000_0000;
array[43319] <= 16'b0000_0000_0000_0000;
array[43320] <= 16'b0000_0000_0000_0000;
array[43321] <= 16'b0000_0000_0000_0000;
array[43322] <= 16'b0000_0000_0000_0000;
array[43323] <= 16'b0000_0000_0000_0000;
array[43324] <= 16'b0000_0000_0000_0000;
array[43325] <= 16'b0000_0000_0000_0000;
array[43326] <= 16'b0000_0000_0000_0000;
array[43327] <= 16'b0000_0000_0000_0000;
array[43328] <= 16'b0000_0000_0000_0000;
array[43329] <= 16'b0000_0000_0000_0000;
array[43330] <= 16'b0000_0000_0000_0000;
array[43331] <= 16'b0000_0000_0000_0000;
array[43332] <= 16'b0000_0000_0000_0000;
array[43333] <= 16'b0000_0000_0000_0000;
array[43334] <= 16'b0000_0000_0000_0000;
array[43335] <= 16'b0000_0000_0000_0000;
array[43336] <= 16'b0000_0000_0000_0000;
array[43337] <= 16'b0000_0000_0000_0000;
array[43338] <= 16'b0000_0000_0000_0000;
array[43339] <= 16'b0000_0000_0000_0000;
array[43340] <= 16'b0000_0000_0000_0000;
array[43341] <= 16'b0000_0000_0000_0000;
array[43342] <= 16'b0000_0000_0000_0000;
array[43343] <= 16'b0000_0000_0000_0000;
array[43344] <= 16'b0000_0000_0000_0000;
array[43345] <= 16'b0000_0000_0000_0000;
array[43346] <= 16'b0000_0000_0000_0000;
array[43347] <= 16'b0000_0000_0000_0000;
array[43348] <= 16'b0000_0000_0000_0000;
array[43349] <= 16'b0000_0000_0000_0000;
array[43350] <= 16'b0000_0000_0000_0000;
array[43351] <= 16'b0000_0000_0000_0000;
array[43352] <= 16'b0000_0000_0000_0000;
array[43353] <= 16'b0000_0000_0000_0000;
array[43354] <= 16'b0000_0000_0000_0000;
array[43355] <= 16'b0000_0000_0000_0000;
array[43356] <= 16'b0000_0000_0000_0000;
array[43357] <= 16'b0000_0000_0000_0000;
array[43358] <= 16'b0000_0000_0000_0000;
array[43359] <= 16'b0000_0000_0000_0000;
array[43360] <= 16'b0000_0000_0000_0000;
array[43361] <= 16'b0000_0000_0000_0000;
array[43362] <= 16'b0000_0000_0000_0000;
array[43363] <= 16'b0000_0000_0000_0000;
array[43364] <= 16'b0000_0000_0000_0000;
array[43365] <= 16'b0000_0000_0000_0000;
array[43366] <= 16'b0000_0000_0000_0000;
array[43367] <= 16'b0000_0000_0000_0000;
array[43368] <= 16'b0000_0000_0000_0000;
array[43369] <= 16'b0000_0000_0000_0000;
array[43370] <= 16'b0000_0000_0000_0000;
array[43371] <= 16'b0000_0000_0000_0000;
array[43372] <= 16'b0000_0000_0000_0000;
array[43373] <= 16'b0000_0000_0000_0000;
array[43374] <= 16'b0000_0000_0000_0000;
array[43375] <= 16'b0000_0000_0000_0000;
array[43376] <= 16'b0000_0000_0000_0000;
array[43377] <= 16'b0000_0000_0000_0000;
array[43378] <= 16'b0000_0000_0000_0000;
array[43379] <= 16'b0000_0000_0000_0000;
array[43380] <= 16'b0000_0000_0000_0000;
array[43381] <= 16'b0000_0000_0000_0000;
array[43382] <= 16'b0000_0000_0000_0000;
array[43383] <= 16'b0000_0000_0000_0000;
array[43384] <= 16'b0000_0000_0000_0000;
array[43385] <= 16'b0000_0000_0000_0000;
array[43386] <= 16'b0000_0000_0000_0000;
array[43387] <= 16'b0000_0000_0000_0000;
array[43388] <= 16'b0000_0000_0000_0000;
array[43389] <= 16'b0000_0000_0000_0000;
array[43390] <= 16'b0000_0000_0000_0000;
array[43391] <= 16'b0000_0000_0000_0000;
array[43392] <= 16'b0000_0000_0000_0000;
array[43393] <= 16'b0000_0000_0000_0000;
array[43394] <= 16'b0000_0000_0000_0000;
array[43395] <= 16'b0000_0000_0000_0000;
array[43396] <= 16'b0000_0000_0000_0000;
array[43397] <= 16'b0000_0000_0000_0000;
array[43398] <= 16'b0000_0000_0000_0000;
array[43399] <= 16'b0000_0000_0000_0000;
array[43400] <= 16'b0000_0000_0000_0000;
array[43401] <= 16'b0000_0000_0000_0000;
array[43402] <= 16'b0000_0000_0000_0000;
array[43403] <= 16'b0000_0000_0000_0000;
array[43404] <= 16'b0000_0000_0000_0000;
array[43405] <= 16'b0000_0000_0000_0000;
array[43406] <= 16'b0000_0000_0000_0000;
array[43407] <= 16'b0000_0000_0000_0000;
array[43408] <= 16'b0000_0000_0000_0000;
array[43409] <= 16'b0000_0000_0000_0000;
array[43410] <= 16'b0000_0000_0000_0000;
array[43411] <= 16'b0000_0000_0000_0000;
array[43412] <= 16'b0000_0000_0000_0000;
array[43413] <= 16'b0000_0000_0000_0000;
array[43414] <= 16'b0000_0000_0000_0000;
array[43415] <= 16'b0000_0000_0000_0000;
array[43416] <= 16'b0000_0000_0000_0000;
array[43417] <= 16'b0000_0000_0000_0000;
array[43418] <= 16'b0000_0000_0000_0000;
array[43419] <= 16'b0000_0000_0000_0000;
array[43420] <= 16'b0000_0000_0000_0000;
array[43421] <= 16'b0000_0000_0000_0000;
array[43422] <= 16'b0000_0000_0000_0000;
array[43423] <= 16'b0000_0000_0000_0000;
array[43424] <= 16'b0000_0000_0000_0000;
array[43425] <= 16'b0000_0000_0000_0000;
array[43426] <= 16'b0000_0000_0000_0000;
array[43427] <= 16'b0000_0000_0000_0000;
array[43428] <= 16'b0000_0000_0000_0000;
array[43429] <= 16'b0000_0000_0000_0000;
array[43430] <= 16'b0000_0000_0000_0000;
array[43431] <= 16'b0000_0000_0000_0000;
array[43432] <= 16'b0000_0000_0000_0000;
array[43433] <= 16'b0000_0000_0000_0000;
array[43434] <= 16'b0000_0000_0000_0000;
array[43435] <= 16'b0000_0000_0000_0000;
array[43436] <= 16'b0000_0000_0000_0000;
array[43437] <= 16'b0000_0000_0000_0000;
array[43438] <= 16'b0000_0000_0000_0000;
array[43439] <= 16'b0000_0000_0000_0000;
array[43440] <= 16'b0000_0000_0000_0000;
array[43441] <= 16'b0000_0000_0000_0000;
array[43442] <= 16'b0000_0000_0000_0000;
array[43443] <= 16'b0000_0000_0000_0000;
array[43444] <= 16'b0000_0000_0000_0000;
array[43445] <= 16'b0000_0000_0000_0000;
array[43446] <= 16'b0000_0000_0000_0000;
array[43447] <= 16'b0000_0000_0000_0000;
array[43448] <= 16'b0000_0000_0000_0000;
array[43449] <= 16'b0000_0000_0000_0000;
array[43450] <= 16'b0000_0000_0000_0000;
array[43451] <= 16'b0000_0000_0000_0000;
array[43452] <= 16'b0000_0000_0000_0000;
array[43453] <= 16'b0000_0000_0000_0000;
array[43454] <= 16'b0000_0000_0000_0000;
array[43455] <= 16'b0000_0000_0000_0000;
array[43456] <= 16'b0000_0000_0000_0000;
array[43457] <= 16'b0000_0000_0000_0000;
array[43458] <= 16'b0000_0000_0000_0000;
array[43459] <= 16'b0000_0000_0000_0000;
array[43460] <= 16'b0000_0000_0000_0000;
array[43461] <= 16'b0000_0000_0000_0000;
array[43462] <= 16'b0000_0000_0000_0000;
array[43463] <= 16'b0000_0000_0000_0000;
array[43464] <= 16'b0000_0000_0000_0000;
array[43465] <= 16'b0000_0000_0000_0000;
array[43466] <= 16'b0000_0000_0000_0000;
array[43467] <= 16'b0000_0000_0000_0000;
array[43468] <= 16'b0000_0000_0000_0000;
array[43469] <= 16'b0000_0000_0000_0000;
array[43470] <= 16'b0000_0000_0000_0000;
array[43471] <= 16'b0000_0000_0000_0000;
array[43472] <= 16'b0000_0000_0000_0000;
array[43473] <= 16'b0000_0000_0000_0000;
array[43474] <= 16'b0000_0000_0000_0000;
array[43475] <= 16'b0000_0000_0000_0000;
array[43476] <= 16'b0000_0000_0000_0000;
array[43477] <= 16'b0000_0000_0000_0000;
array[43478] <= 16'b0000_0000_0000_0000;
array[43479] <= 16'b0000_0000_0000_0000;
array[43480] <= 16'b0000_0000_0000_0000;
array[43481] <= 16'b0000_0000_0000_0000;
array[43482] <= 16'b0000_0000_0000_0000;
array[43483] <= 16'b0000_0000_0000_0000;
array[43484] <= 16'b0000_0000_0000_0000;
array[43485] <= 16'b0000_0000_0000_0000;
array[43486] <= 16'b0000_0000_0000_0000;
array[43487] <= 16'b0000_0000_0000_0000;
array[43488] <= 16'b0000_0000_0000_0000;
array[43489] <= 16'b0000_0000_0000_0000;
array[43490] <= 16'b0000_0000_0000_0000;
array[43491] <= 16'b0000_0000_0000_0000;
array[43492] <= 16'b0000_0000_0000_0000;
array[43493] <= 16'b0000_0000_0000_0000;
array[43494] <= 16'b0000_0000_0000_0000;
array[43495] <= 16'b0000_0000_0000_0000;
array[43496] <= 16'b0000_0000_0000_0000;
array[43497] <= 16'b0000_0000_0000_0000;
array[43498] <= 16'b0000_0000_0000_0000;
array[43499] <= 16'b0000_0000_0000_0000;
array[43500] <= 16'b0000_0000_0000_0000;
array[43501] <= 16'b0000_0000_0000_0000;
array[43502] <= 16'b0000_0000_0000_0000;
array[43503] <= 16'b0000_0000_0000_0000;
array[43504] <= 16'b0000_0000_0000_0000;
array[43505] <= 16'b0000_0000_0000_0000;
array[43506] <= 16'b0000_0000_0000_0000;
array[43507] <= 16'b0000_0000_0000_0000;
array[43508] <= 16'b0000_0000_0000_0000;
array[43509] <= 16'b0000_0000_0000_0000;
array[43510] <= 16'b0000_0000_0000_0000;
array[43511] <= 16'b0000_0000_0000_0000;
array[43512] <= 16'b0000_0000_0000_0000;
array[43513] <= 16'b0000_0000_0000_0000;
array[43514] <= 16'b0000_0000_0000_0000;
array[43515] <= 16'b0000_0000_0000_0000;
array[43516] <= 16'b0000_0000_0000_0000;
array[43517] <= 16'b0000_0000_0000_0000;
array[43518] <= 16'b0000_0000_0000_0000;
array[43519] <= 16'b0000_0000_0000_0000;
array[43520] <= 16'b0000_0000_0000_0000;
array[43521] <= 16'b0000_0000_0000_0000;
array[43522] <= 16'b0000_0000_0000_0000;
array[43523] <= 16'b0000_0000_0000_0000;
array[43524] <= 16'b0000_0000_0000_0000;
array[43525] <= 16'b0000_0000_0000_0000;
array[43526] <= 16'b0000_0000_0000_0000;
array[43527] <= 16'b0000_0000_0000_0000;
array[43528] <= 16'b0000_0000_0000_0000;
array[43529] <= 16'b0000_0000_0000_0000;
array[43530] <= 16'b0000_0000_0000_0000;
array[43531] <= 16'b0000_0000_0000_0000;
array[43532] <= 16'b0000_0000_0000_0000;
array[43533] <= 16'b0000_0000_0000_0000;
array[43534] <= 16'b0000_0000_0000_0000;
array[43535] <= 16'b0000_0000_0000_0000;
array[43536] <= 16'b0000_0000_0000_0000;
array[43537] <= 16'b0000_0000_0000_0000;
array[43538] <= 16'b0000_0000_0000_0000;
array[43539] <= 16'b0000_0000_0000_0000;
array[43540] <= 16'b0000_0000_0000_0000;
array[43541] <= 16'b0000_0000_0000_0000;
array[43542] <= 16'b0000_0000_0000_0000;
array[43543] <= 16'b0000_0000_0000_0000;
array[43544] <= 16'b0000_0000_0000_0000;
array[43545] <= 16'b0000_0000_0000_0000;
array[43546] <= 16'b0000_0000_0000_0000;
array[43547] <= 16'b0000_0000_0000_0000;
array[43548] <= 16'b0000_0000_0000_0000;
array[43549] <= 16'b0000_0000_0000_0000;
array[43550] <= 16'b0000_0000_0000_0000;
array[43551] <= 16'b0000_0000_0000_0000;
array[43552] <= 16'b0000_0000_0000_0000;
array[43553] <= 16'b0000_0000_0000_0000;
array[43554] <= 16'b0000_0000_0000_0000;
array[43555] <= 16'b0000_0000_0000_0000;
array[43556] <= 16'b0000_0000_0000_0000;
array[43557] <= 16'b0000_0000_0000_0000;
array[43558] <= 16'b0000_0000_0000_0000;
array[43559] <= 16'b0000_0000_0000_0000;
array[43560] <= 16'b0000_0000_0000_0000;
array[43561] <= 16'b0000_0000_0000_0000;
array[43562] <= 16'b0000_0000_0000_0000;
array[43563] <= 16'b0000_0000_0000_0000;
array[43564] <= 16'b0000_0000_0000_0000;
array[43565] <= 16'b0000_0000_0000_0000;
array[43566] <= 16'b0000_0000_0000_0000;
array[43567] <= 16'b0000_0000_0000_0000;
array[43568] <= 16'b0000_0000_0000_0000;
array[43569] <= 16'b0000_0000_0000_0000;
array[43570] <= 16'b0000_0000_0000_0000;
array[43571] <= 16'b0000_0000_0000_0000;
array[43572] <= 16'b0000_0000_0000_0000;
array[43573] <= 16'b0000_0000_0000_0000;
array[43574] <= 16'b0000_0000_0000_0000;
array[43575] <= 16'b0000_0000_0000_0000;
array[43576] <= 16'b0000_0000_0000_0000;
array[43577] <= 16'b0000_0000_0000_0000;
array[43578] <= 16'b0000_0000_0000_0000;
array[43579] <= 16'b0000_0000_0000_0000;
array[43580] <= 16'b0000_0000_0000_0000;
array[43581] <= 16'b0000_0000_0000_0000;
array[43582] <= 16'b0000_0000_0000_0000;
array[43583] <= 16'b0000_0000_0000_0000;
array[43584] <= 16'b0000_0000_0000_0000;
array[43585] <= 16'b0000_0000_0000_0000;
array[43586] <= 16'b0000_0000_0000_0000;
array[43587] <= 16'b0000_0000_0000_0000;
array[43588] <= 16'b0000_0000_0000_0000;
array[43589] <= 16'b0000_0000_0000_0000;
array[43590] <= 16'b0000_0000_0000_0000;
array[43591] <= 16'b0000_0000_0000_0000;
array[43592] <= 16'b0000_0000_0000_0000;
array[43593] <= 16'b0000_0000_0000_0000;
array[43594] <= 16'b0000_0000_0000_0000;
array[43595] <= 16'b0000_0000_0000_0000;
array[43596] <= 16'b0000_0000_0000_0000;
array[43597] <= 16'b0000_0000_0000_0000;
array[43598] <= 16'b0000_0000_0000_0000;
array[43599] <= 16'b0000_0000_0000_0000;
array[43600] <= 16'b0000_0000_0000_0000;
array[43601] <= 16'b0000_0000_0000_0000;
array[43602] <= 16'b0000_0000_0000_0000;
array[43603] <= 16'b0000_0000_0000_0000;
array[43604] <= 16'b0000_0000_0000_0000;
array[43605] <= 16'b0000_0000_0000_0000;
array[43606] <= 16'b0000_0000_0000_0000;
array[43607] <= 16'b0000_0000_0000_0000;
array[43608] <= 16'b0000_0000_0000_0000;
array[43609] <= 16'b0000_0000_0000_0000;
array[43610] <= 16'b0000_0000_0000_0000;
array[43611] <= 16'b0000_0000_0000_0000;
array[43612] <= 16'b0000_0000_0000_0000;
array[43613] <= 16'b0000_0000_0000_0000;
array[43614] <= 16'b0000_0000_0000_0000;
array[43615] <= 16'b0000_0000_0000_0000;
array[43616] <= 16'b0000_0000_0000_0000;
array[43617] <= 16'b0000_0000_0000_0000;
array[43618] <= 16'b0000_0000_0000_0000;
array[43619] <= 16'b0000_0000_0000_0000;
array[43620] <= 16'b0000_0000_0000_0000;
array[43621] <= 16'b0000_0000_0000_0000;
array[43622] <= 16'b0000_0000_0000_0000;
array[43623] <= 16'b0000_0000_0000_0000;
array[43624] <= 16'b0000_0000_0000_0000;
array[43625] <= 16'b0000_0000_0000_0000;
array[43626] <= 16'b0000_0000_0000_0000;
array[43627] <= 16'b0000_0000_0000_0000;
array[43628] <= 16'b0000_0000_0000_0000;
array[43629] <= 16'b0000_0000_0000_0000;
array[43630] <= 16'b0000_0000_0000_0000;
array[43631] <= 16'b0000_0000_0000_0000;
array[43632] <= 16'b0000_0000_0000_0000;
array[43633] <= 16'b0000_0000_0000_0000;
array[43634] <= 16'b0000_0000_0000_0000;
array[43635] <= 16'b0000_0000_0000_0000;
array[43636] <= 16'b0000_0000_0000_0000;
array[43637] <= 16'b0000_0000_0000_0000;
array[43638] <= 16'b0000_0000_0000_0000;
array[43639] <= 16'b0000_0000_0000_0000;
array[43640] <= 16'b0000_0000_0000_0000;
array[43641] <= 16'b0000_0000_0000_0000;
array[43642] <= 16'b0000_0000_0000_0000;
array[43643] <= 16'b0000_0000_0000_0000;
array[43644] <= 16'b0000_0000_0000_0000;
array[43645] <= 16'b0000_0000_0000_0000;
array[43646] <= 16'b0000_0000_0000_0000;
array[43647] <= 16'b0000_0000_0000_0000;
array[43648] <= 16'b0000_0000_0000_0000;
array[43649] <= 16'b0000_0000_0000_0000;
array[43650] <= 16'b0000_0000_0000_0000;
array[43651] <= 16'b0000_0000_0000_0000;
array[43652] <= 16'b0000_0000_0000_0000;
array[43653] <= 16'b0000_0000_0000_0000;
array[43654] <= 16'b0000_0000_0000_0000;
array[43655] <= 16'b0000_0000_0000_0000;
array[43656] <= 16'b0000_0000_0000_0000;
array[43657] <= 16'b0000_0000_0000_0000;
array[43658] <= 16'b0000_0000_0000_0000;
array[43659] <= 16'b0000_0000_0000_0000;
array[43660] <= 16'b0000_0000_0000_0000;
array[43661] <= 16'b0000_0000_0000_0000;
array[43662] <= 16'b0000_0000_0000_0000;
array[43663] <= 16'b0000_0000_0000_0000;
array[43664] <= 16'b0000_0000_0000_0000;
array[43665] <= 16'b0000_0000_0000_0000;
array[43666] <= 16'b0000_0000_0000_0000;
array[43667] <= 16'b0000_0000_0000_0000;
array[43668] <= 16'b0000_0000_0000_0000;
array[43669] <= 16'b0000_0000_0000_0000;
array[43670] <= 16'b0000_0000_0000_0000;
array[43671] <= 16'b0000_0000_0000_0000;
array[43672] <= 16'b0000_0000_0000_0000;
array[43673] <= 16'b0000_0000_0000_0000;
array[43674] <= 16'b0000_0000_0000_0000;
array[43675] <= 16'b0000_0000_0000_0000;
array[43676] <= 16'b0000_0000_0000_0000;
array[43677] <= 16'b0000_0000_0000_0000;
array[43678] <= 16'b0000_0000_0000_0000;
array[43679] <= 16'b0000_0000_0000_0000;
array[43680] <= 16'b0000_0000_0000_0000;
array[43681] <= 16'b0000_0000_0000_0000;
array[43682] <= 16'b0000_0000_0000_0000;
array[43683] <= 16'b0000_0000_0000_0000;
array[43684] <= 16'b0000_0000_0000_0000;
array[43685] <= 16'b0000_0000_0000_0000;
array[43686] <= 16'b0000_0000_0000_0000;
array[43687] <= 16'b0000_0000_0000_0000;
array[43688] <= 16'b0000_0000_0000_0000;
array[43689] <= 16'b0000_0000_0000_0000;
array[43690] <= 16'b0000_0000_0000_0000;
array[43691] <= 16'b0000_0000_0000_0000;
array[43692] <= 16'b0000_0000_0000_0000;
array[43693] <= 16'b0000_0000_0000_0000;
array[43694] <= 16'b0000_0000_0000_0000;
array[43695] <= 16'b0000_0000_0000_0000;
array[43696] <= 16'b0000_0000_0000_0000;
array[43697] <= 16'b0000_0000_0000_0000;
array[43698] <= 16'b0000_0000_0000_0000;
array[43699] <= 16'b0000_0000_0000_0000;
array[43700] <= 16'b0000_0000_0000_0000;
array[43701] <= 16'b0000_0000_0000_0000;
array[43702] <= 16'b0000_0000_0000_0000;
array[43703] <= 16'b0000_0000_0000_0000;
array[43704] <= 16'b0000_0000_0000_0000;
array[43705] <= 16'b0000_0000_0000_0000;
array[43706] <= 16'b0000_0000_0000_0000;
array[43707] <= 16'b0000_0000_0000_0000;
array[43708] <= 16'b0000_0000_0000_0000;
array[43709] <= 16'b0000_0000_0000_0000;
array[43710] <= 16'b0000_0000_0000_0000;
array[43711] <= 16'b0000_0000_0000_0000;
array[43712] <= 16'b0000_0000_0000_0000;
array[43713] <= 16'b0000_0000_0000_0000;
array[43714] <= 16'b0000_0000_0000_0000;
array[43715] <= 16'b0000_0000_0000_0000;
array[43716] <= 16'b0000_0000_0000_0000;
array[43717] <= 16'b0000_0000_0000_0000;
array[43718] <= 16'b0000_0000_0000_0000;
array[43719] <= 16'b0000_0000_0000_0000;
array[43720] <= 16'b0000_0000_0000_0000;
array[43721] <= 16'b0000_0000_0000_0000;
array[43722] <= 16'b0000_0000_0000_0000;
array[43723] <= 16'b0000_0000_0000_0000;
array[43724] <= 16'b0000_0000_0000_0000;
array[43725] <= 16'b0000_0000_0000_0000;
array[43726] <= 16'b0000_0000_0000_0000;
array[43727] <= 16'b0000_0000_0000_0000;
array[43728] <= 16'b0000_0000_0000_0000;
array[43729] <= 16'b0000_0000_0000_0000;
array[43730] <= 16'b0000_0000_0000_0000;
array[43731] <= 16'b0000_0000_0000_0000;
array[43732] <= 16'b0000_0000_0000_0000;
array[43733] <= 16'b0000_0000_0000_0000;
array[43734] <= 16'b0000_0000_0000_0000;
array[43735] <= 16'b0000_0000_0000_0000;
array[43736] <= 16'b0000_0000_0000_0000;
array[43737] <= 16'b0000_0000_0000_0000;
array[43738] <= 16'b0000_0000_0000_0000;
array[43739] <= 16'b0000_0000_0000_0000;
array[43740] <= 16'b0000_0000_0000_0000;
array[43741] <= 16'b0000_0000_0000_0000;
array[43742] <= 16'b0000_0000_0000_0000;
array[43743] <= 16'b0000_0000_0000_0000;
array[43744] <= 16'b0000_0000_0000_0000;
array[43745] <= 16'b0000_0000_0000_0000;
array[43746] <= 16'b0000_0000_0000_0000;
array[43747] <= 16'b0000_0000_0000_0000;
array[43748] <= 16'b0000_0000_0000_0000;
array[43749] <= 16'b0000_0000_0000_0000;
array[43750] <= 16'b0000_0000_0000_0000;
array[43751] <= 16'b0000_0000_0000_0000;
array[43752] <= 16'b0000_0000_0000_0000;
array[43753] <= 16'b0000_0000_0000_0000;
array[43754] <= 16'b0000_0000_0000_0000;
array[43755] <= 16'b0000_0000_0000_0000;
array[43756] <= 16'b0000_0000_0000_0000;
array[43757] <= 16'b0000_0000_0000_0000;
array[43758] <= 16'b0000_0000_0000_0000;
array[43759] <= 16'b0000_0000_0000_0000;
array[43760] <= 16'b0000_0000_0000_0000;
array[43761] <= 16'b0000_0000_0000_0000;
array[43762] <= 16'b0000_0000_0000_0000;
array[43763] <= 16'b0000_0000_0000_0000;
array[43764] <= 16'b0000_0000_0000_0000;
array[43765] <= 16'b0000_0000_0000_0000;
array[43766] <= 16'b0000_0000_0000_0000;
array[43767] <= 16'b0000_0000_0000_0000;
array[43768] <= 16'b0000_0000_0000_0000;
array[43769] <= 16'b0000_0000_0000_0000;
array[43770] <= 16'b0000_0000_0000_0000;
array[43771] <= 16'b0000_0000_0000_0000;
array[43772] <= 16'b0000_0000_0000_0000;
array[43773] <= 16'b0000_0000_0000_0000;
array[43774] <= 16'b0000_0000_0000_0000;
array[43775] <= 16'b0000_0000_0000_0000;
array[43776] <= 16'b0000_0000_0000_0000;
array[43777] <= 16'b0000_0000_0000_0000;
array[43778] <= 16'b0000_0000_0000_0000;
array[43779] <= 16'b0000_0000_0000_0000;
array[43780] <= 16'b0000_0000_0000_0000;
array[43781] <= 16'b0000_0000_0000_0000;
array[43782] <= 16'b0000_0000_0000_0000;
array[43783] <= 16'b0000_0000_0000_0000;
array[43784] <= 16'b0000_0000_0000_0000;
array[43785] <= 16'b0000_0000_0000_0000;
array[43786] <= 16'b0000_0000_0000_0000;
array[43787] <= 16'b0000_0000_0000_0000;
array[43788] <= 16'b0000_0000_0000_0000;
array[43789] <= 16'b0000_0000_0000_0000;
array[43790] <= 16'b0000_0000_0000_0000;
array[43791] <= 16'b0000_0000_0000_0000;
array[43792] <= 16'b0000_0000_0000_0000;
array[43793] <= 16'b0000_0000_0000_0000;
array[43794] <= 16'b0000_0000_0000_0000;
array[43795] <= 16'b0000_0000_0000_0000;
array[43796] <= 16'b0000_0000_0000_0000;
array[43797] <= 16'b0000_0000_0000_0000;
array[43798] <= 16'b0000_0000_0000_0000;
array[43799] <= 16'b0000_0000_0000_0000;
array[43800] <= 16'b0000_0000_0000_0000;
array[43801] <= 16'b0000_0000_0000_0000;
array[43802] <= 16'b0000_0000_0000_0000;
array[43803] <= 16'b0000_0000_0000_0000;
array[43804] <= 16'b0000_0000_0000_0000;
array[43805] <= 16'b0000_0000_0000_0000;
array[43806] <= 16'b0000_0000_0000_0000;
array[43807] <= 16'b0000_0000_0000_0000;
array[43808] <= 16'b0000_0000_0000_0000;
array[43809] <= 16'b0000_0000_0000_0000;
array[43810] <= 16'b0000_0000_0000_0000;
array[43811] <= 16'b0000_0000_0000_0000;
array[43812] <= 16'b0000_0000_0000_0000;
array[43813] <= 16'b0000_0000_0000_0000;
array[43814] <= 16'b0000_0000_0000_0000;
array[43815] <= 16'b0000_0000_0000_0000;
array[43816] <= 16'b0000_0000_0000_0000;
array[43817] <= 16'b0000_0000_0000_0000;
array[43818] <= 16'b0000_0000_0000_0000;
array[43819] <= 16'b0000_0000_0000_0000;
array[43820] <= 16'b0000_0000_0000_0000;
array[43821] <= 16'b0000_0000_0000_0000;
array[43822] <= 16'b0000_0000_0000_0000;
array[43823] <= 16'b0000_0000_0000_0000;
array[43824] <= 16'b0000_0000_0000_0000;
array[43825] <= 16'b0000_0000_0000_0000;
array[43826] <= 16'b0000_0000_0000_0000;
array[43827] <= 16'b0000_0000_0000_0000;
array[43828] <= 16'b0000_0000_0000_0000;
array[43829] <= 16'b0000_0000_0000_0000;
array[43830] <= 16'b0000_0000_0000_0000;
array[43831] <= 16'b0000_0000_0000_0000;
array[43832] <= 16'b0000_0000_0000_0000;
array[43833] <= 16'b0000_0000_0000_0000;
array[43834] <= 16'b0000_0000_0000_0000;
array[43835] <= 16'b0000_0000_0000_0000;
array[43836] <= 16'b0000_0000_0000_0000;
array[43837] <= 16'b0000_0000_0000_0000;
array[43838] <= 16'b0000_0000_0000_0000;
array[43839] <= 16'b0000_0000_0000_0000;
array[43840] <= 16'b0000_0000_0000_0000;
array[43841] <= 16'b0000_0000_0000_0000;
array[43842] <= 16'b0000_0000_0000_0000;
array[43843] <= 16'b0000_0000_0000_0000;
array[43844] <= 16'b0000_0000_0000_0000;
array[43845] <= 16'b0000_0000_0000_0000;
array[43846] <= 16'b0000_0000_0000_0000;
array[43847] <= 16'b0000_0000_0000_0000;
array[43848] <= 16'b0000_0000_0000_0000;
array[43849] <= 16'b0000_0000_0000_0000;
array[43850] <= 16'b0000_0000_0000_0000;
array[43851] <= 16'b0000_0000_0000_0000;
array[43852] <= 16'b0000_0000_0000_0000;
array[43853] <= 16'b0000_0000_0000_0000;
array[43854] <= 16'b0000_0000_0000_0000;
array[43855] <= 16'b0000_0000_0000_0000;
array[43856] <= 16'b0000_0000_0000_0000;
array[43857] <= 16'b0000_0000_0000_0000;
array[43858] <= 16'b0000_0000_0000_0000;
array[43859] <= 16'b0000_0000_0000_0000;
array[43860] <= 16'b0000_0000_0000_0000;
array[43861] <= 16'b0000_0000_0000_0000;
array[43862] <= 16'b0000_0000_0000_0000;
array[43863] <= 16'b0000_0000_0000_0000;
array[43864] <= 16'b0000_0000_0000_0000;
array[43865] <= 16'b0000_0000_0000_0000;
array[43866] <= 16'b0000_0000_0000_0000;
array[43867] <= 16'b0000_0000_0000_0000;
array[43868] <= 16'b0000_0000_0000_0000;
array[43869] <= 16'b0000_0000_0000_0000;
array[43870] <= 16'b0000_0000_0000_0000;
array[43871] <= 16'b0000_0000_0000_0000;
array[43872] <= 16'b0000_0000_0000_0000;
array[43873] <= 16'b0000_0000_0000_0000;
array[43874] <= 16'b0000_0000_0000_0000;
array[43875] <= 16'b0000_0000_0000_0000;
array[43876] <= 16'b0000_0000_0000_0000;
array[43877] <= 16'b0000_0000_0000_0000;
array[43878] <= 16'b0000_0000_0000_0000;
array[43879] <= 16'b0000_0000_0000_0000;
array[43880] <= 16'b0000_0000_0000_0000;
array[43881] <= 16'b0000_0000_0000_0000;
array[43882] <= 16'b0000_0000_0000_0000;
array[43883] <= 16'b0000_0000_0000_0000;
array[43884] <= 16'b0000_0000_0000_0000;
array[43885] <= 16'b0000_0000_0000_0000;
array[43886] <= 16'b0000_0000_0000_0000;
array[43887] <= 16'b0000_0000_0000_0000;
array[43888] <= 16'b0000_0000_0000_0000;
array[43889] <= 16'b0000_0000_0000_0000;
array[43890] <= 16'b0000_0000_0000_0000;
array[43891] <= 16'b0000_0000_0000_0000;
array[43892] <= 16'b0000_0000_0000_0000;
array[43893] <= 16'b0000_0000_0000_0000;
array[43894] <= 16'b0000_0000_0000_0000;
array[43895] <= 16'b0000_0000_0000_0000;
array[43896] <= 16'b0000_0000_0000_0000;
array[43897] <= 16'b0000_0000_0000_0000;
array[43898] <= 16'b0000_0000_0000_0000;
array[43899] <= 16'b0000_0000_0000_0000;
array[43900] <= 16'b0000_0000_0000_0000;
array[43901] <= 16'b0000_0000_0000_0000;
array[43902] <= 16'b0000_0000_0000_0000;
array[43903] <= 16'b0000_0000_0000_0000;
array[43904] <= 16'b0000_0000_0000_0000;
array[43905] <= 16'b0000_0000_0000_0000;
array[43906] <= 16'b0000_0000_0000_0000;
array[43907] <= 16'b0000_0000_0000_0000;
array[43908] <= 16'b0000_0000_0000_0000;
array[43909] <= 16'b0000_0000_0000_0000;
array[43910] <= 16'b0000_0000_0000_0000;
array[43911] <= 16'b0000_0000_0000_0000;
array[43912] <= 16'b0000_0000_0000_0000;
array[43913] <= 16'b0000_0000_0000_0000;
array[43914] <= 16'b0000_0000_0000_0000;
array[43915] <= 16'b0000_0000_0000_0000;
array[43916] <= 16'b0000_0000_0000_0000;
array[43917] <= 16'b0000_0000_0000_0000;
array[43918] <= 16'b0000_0000_0000_0000;
array[43919] <= 16'b0000_0000_0000_0000;
array[43920] <= 16'b0000_0000_0000_0000;
array[43921] <= 16'b0000_0000_0000_0000;
array[43922] <= 16'b0000_0000_0000_0000;
array[43923] <= 16'b0000_0000_0000_0000;
array[43924] <= 16'b0000_0000_0000_0000;
array[43925] <= 16'b0000_0000_0000_0000;
array[43926] <= 16'b0000_0000_0000_0000;
array[43927] <= 16'b0000_0000_0000_0000;
array[43928] <= 16'b0000_0000_0000_0000;
array[43929] <= 16'b0000_0000_0000_0000;
array[43930] <= 16'b0000_0000_0000_0000;
array[43931] <= 16'b0000_0000_0000_0000;
array[43932] <= 16'b0000_0000_0000_0000;
array[43933] <= 16'b0000_0000_0000_0000;
array[43934] <= 16'b0000_0000_0000_0000;
array[43935] <= 16'b0000_0000_0000_0000;
array[43936] <= 16'b0000_0000_0000_0000;
array[43937] <= 16'b0000_0000_0000_0000;
array[43938] <= 16'b0000_0000_0000_0000;
array[43939] <= 16'b0000_0000_0000_0000;
array[43940] <= 16'b0000_0000_0000_0000;
array[43941] <= 16'b0000_0000_0000_0000;
array[43942] <= 16'b0000_0000_0000_0000;
array[43943] <= 16'b0000_0000_0000_0000;
array[43944] <= 16'b0000_0000_0000_0000;
array[43945] <= 16'b0000_0000_0000_0000;
array[43946] <= 16'b0000_0000_0000_0000;
array[43947] <= 16'b0000_0000_0000_0000;
array[43948] <= 16'b0000_0000_0000_0000;
array[43949] <= 16'b0000_0000_0000_0000;
array[43950] <= 16'b0000_0000_0000_0000;
array[43951] <= 16'b0000_0000_0000_0000;
array[43952] <= 16'b0000_0000_0000_0000;
array[43953] <= 16'b0000_0000_0000_0000;
array[43954] <= 16'b0000_0000_0000_0000;
array[43955] <= 16'b0000_0000_0000_0000;
array[43956] <= 16'b0000_0000_0000_0000;
array[43957] <= 16'b0000_0000_0000_0000;
array[43958] <= 16'b0000_0000_0000_0000;
array[43959] <= 16'b0000_0000_0000_0000;
array[43960] <= 16'b0000_0000_0000_0000;
array[43961] <= 16'b0000_0000_0000_0000;
array[43962] <= 16'b0000_0000_0000_0000;
array[43963] <= 16'b0000_0000_0000_0000;
array[43964] <= 16'b0000_0000_0000_0000;
array[43965] <= 16'b0000_0000_0000_0000;
array[43966] <= 16'b0000_0000_0000_0000;
array[43967] <= 16'b0000_0000_0000_0000;
array[43968] <= 16'b0000_0000_0000_0000;
array[43969] <= 16'b0000_0000_0000_0000;
array[43970] <= 16'b0000_0000_0000_0000;
array[43971] <= 16'b0000_0000_0000_0000;
array[43972] <= 16'b0000_0000_0000_0000;
array[43973] <= 16'b0000_0000_0000_0000;
array[43974] <= 16'b0000_0000_0000_0000;
array[43975] <= 16'b0000_0000_0000_0000;
array[43976] <= 16'b0000_0000_0000_0000;
array[43977] <= 16'b0000_0000_0000_0000;
array[43978] <= 16'b0000_0000_0000_0000;
array[43979] <= 16'b0000_0000_0000_0000;
array[43980] <= 16'b0000_0000_0000_0000;
array[43981] <= 16'b0000_0000_0000_0000;
array[43982] <= 16'b0000_0000_0000_0000;
array[43983] <= 16'b0000_0000_0000_0000;
array[43984] <= 16'b0000_0000_0000_0000;
array[43985] <= 16'b0000_0000_0000_0000;
array[43986] <= 16'b0000_0000_0000_0000;
array[43987] <= 16'b0000_0000_0000_0000;
array[43988] <= 16'b0000_0000_0000_0000;
array[43989] <= 16'b0000_0000_0000_0000;
array[43990] <= 16'b0000_0000_0000_0000;
array[43991] <= 16'b0000_0000_0000_0000;
array[43992] <= 16'b0000_0000_0000_0000;
array[43993] <= 16'b0000_0000_0000_0000;
array[43994] <= 16'b0000_0000_0000_0000;
array[43995] <= 16'b0000_0000_0000_0000;
array[43996] <= 16'b0000_0000_0000_0000;
array[43997] <= 16'b0000_0000_0000_0000;
array[43998] <= 16'b0000_0000_0000_0000;
array[43999] <= 16'b0000_0000_0000_0000;
array[44000] <= 16'b0000_0000_0000_0000;
array[44001] <= 16'b0000_0000_0000_0000;
array[44002] <= 16'b0000_0000_0000_0000;
array[44003] <= 16'b0000_0000_0000_0000;
array[44004] <= 16'b0000_0000_0000_0000;
array[44005] <= 16'b0000_0000_0000_0000;
array[44006] <= 16'b0000_0000_0000_0000;
array[44007] <= 16'b0000_0000_0000_0000;
array[44008] <= 16'b0000_0000_0000_0000;
array[44009] <= 16'b0000_0000_0000_0000;
array[44010] <= 16'b0000_0000_0000_0000;
array[44011] <= 16'b0000_0000_0000_0000;
array[44012] <= 16'b0000_0000_0000_0000;
array[44013] <= 16'b0000_0000_0000_0000;
array[44014] <= 16'b0000_0000_0000_0000;
array[44015] <= 16'b0000_0000_0000_0000;
array[44016] <= 16'b0000_0000_0000_0000;
array[44017] <= 16'b0000_0000_0000_0000;
array[44018] <= 16'b0000_0000_0000_0000;
array[44019] <= 16'b0000_0000_0000_0000;
array[44020] <= 16'b0000_0000_0000_0000;
array[44021] <= 16'b0000_0000_0000_0000;
array[44022] <= 16'b0000_0000_0000_0000;
array[44023] <= 16'b0000_0000_0000_0000;
array[44024] <= 16'b0000_0000_0000_0000;
array[44025] <= 16'b0000_0000_0000_0000;
array[44026] <= 16'b0000_0000_0000_0000;
array[44027] <= 16'b0000_0000_0000_0000;
array[44028] <= 16'b0000_0000_0000_0000;
array[44029] <= 16'b0000_0000_0000_0000;
array[44030] <= 16'b0000_0000_0000_0000;
array[44031] <= 16'b0000_0000_0000_0000;
array[44032] <= 16'b0000_0000_0000_0000;
array[44033] <= 16'b0000_0000_0000_0000;
array[44034] <= 16'b0000_0000_0000_0000;
array[44035] <= 16'b0000_0000_0000_0000;
array[44036] <= 16'b0000_0000_0000_0000;
array[44037] <= 16'b0000_0000_0000_0000;
array[44038] <= 16'b0000_0000_0000_0000;
array[44039] <= 16'b0000_0000_0000_0000;
array[44040] <= 16'b0000_0000_0000_0000;
array[44041] <= 16'b0000_0000_0000_0000;
array[44042] <= 16'b0000_0000_0000_0000;
array[44043] <= 16'b0000_0000_0000_0000;
array[44044] <= 16'b0000_0000_0000_0000;
array[44045] <= 16'b0000_0000_0000_0000;
array[44046] <= 16'b0000_0000_0000_0000;
array[44047] <= 16'b0000_0000_0000_0000;
array[44048] <= 16'b0000_0000_0000_0000;
array[44049] <= 16'b0000_0000_0000_0000;
array[44050] <= 16'b0000_0000_0000_0000;
array[44051] <= 16'b0000_0000_0000_0000;
array[44052] <= 16'b0000_0000_0000_0000;
array[44053] <= 16'b0000_0000_0000_0000;
array[44054] <= 16'b0000_0000_0000_0000;
array[44055] <= 16'b0000_0000_0000_0000;
array[44056] <= 16'b0000_0000_0000_0000;
array[44057] <= 16'b0000_0000_0000_0000;
array[44058] <= 16'b0000_0000_0000_0000;
array[44059] <= 16'b0000_0000_0000_0000;
array[44060] <= 16'b0000_0000_0000_0000;
array[44061] <= 16'b0000_0000_0000_0000;
array[44062] <= 16'b0000_0000_0000_0000;
array[44063] <= 16'b0000_0000_0000_0000;
array[44064] <= 16'b0000_0000_0000_0000;
array[44065] <= 16'b0000_0000_0000_0000;
array[44066] <= 16'b0000_0000_0000_0000;
array[44067] <= 16'b0000_0000_0000_0000;
array[44068] <= 16'b0000_0000_0000_0000;
array[44069] <= 16'b0000_0000_0000_0000;
array[44070] <= 16'b0000_0000_0000_0000;
array[44071] <= 16'b0000_0000_0000_0000;
array[44072] <= 16'b0000_0000_0000_0000;
array[44073] <= 16'b0000_0000_0000_0000;
array[44074] <= 16'b0000_0000_0000_0000;
array[44075] <= 16'b0000_0000_0000_0000;
array[44076] <= 16'b0000_0000_0000_0000;
array[44077] <= 16'b0000_0000_0000_0000;
array[44078] <= 16'b0000_0000_0000_0000;
array[44079] <= 16'b0000_0000_0000_0000;
array[44080] <= 16'b0000_0000_0000_0000;
array[44081] <= 16'b0000_0000_0000_0000;
array[44082] <= 16'b0000_0000_0000_0000;
array[44083] <= 16'b0000_0000_0000_0000;
array[44084] <= 16'b0000_0000_0000_0000;
array[44085] <= 16'b0000_0000_0000_0000;
array[44086] <= 16'b0000_0000_0000_0000;
array[44087] <= 16'b0000_0000_0000_0000;
array[44088] <= 16'b0000_0000_0000_0000;
array[44089] <= 16'b0000_0000_0000_0000;
array[44090] <= 16'b0000_0000_0000_0000;
array[44091] <= 16'b0000_0000_0000_0000;
array[44092] <= 16'b0000_0000_0000_0000;
array[44093] <= 16'b0000_0000_0000_0000;
array[44094] <= 16'b0000_0000_0000_0000;
array[44095] <= 16'b0000_0000_0000_0000;
array[44096] <= 16'b0000_0000_0000_0000;
array[44097] <= 16'b0000_0000_0000_0000;
array[44098] <= 16'b0000_0000_0000_0000;
array[44099] <= 16'b0000_0000_0000_0000;
array[44100] <= 16'b0000_0000_0000_0000;
array[44101] <= 16'b0000_0000_0000_0000;
array[44102] <= 16'b0000_0000_0000_0000;
array[44103] <= 16'b0000_0000_0000_0000;
array[44104] <= 16'b0000_0000_0000_0000;
array[44105] <= 16'b0000_0000_0000_0000;
array[44106] <= 16'b0000_0000_0000_0000;
array[44107] <= 16'b0000_0000_0000_0000;
array[44108] <= 16'b0000_0000_0000_0000;
array[44109] <= 16'b0000_0000_0000_0000;
array[44110] <= 16'b0000_0000_0000_0000;
array[44111] <= 16'b0000_0000_0000_0000;
array[44112] <= 16'b0000_0000_0000_0000;
array[44113] <= 16'b0000_0000_0000_0000;
array[44114] <= 16'b0000_0000_0000_0000;
array[44115] <= 16'b0000_0000_0000_0000;
array[44116] <= 16'b0000_0000_0000_0000;
array[44117] <= 16'b0000_0000_0000_0000;
array[44118] <= 16'b0000_0000_0000_0000;
array[44119] <= 16'b0000_0000_0000_0000;
array[44120] <= 16'b0000_0000_0000_0000;
array[44121] <= 16'b0000_0000_0000_0000;
array[44122] <= 16'b0000_0000_0000_0000;
array[44123] <= 16'b0000_0000_0000_0000;
array[44124] <= 16'b0000_0000_0000_0000;
array[44125] <= 16'b0000_0000_0000_0000;
array[44126] <= 16'b0000_0000_0000_0000;
array[44127] <= 16'b0000_0000_0000_0000;
array[44128] <= 16'b0000_0000_0000_0000;
array[44129] <= 16'b0000_0000_0000_0000;
array[44130] <= 16'b0000_0000_0000_0000;
array[44131] <= 16'b0000_0000_0000_0000;
array[44132] <= 16'b0000_0000_0000_0000;
array[44133] <= 16'b0000_0000_0000_0000;
array[44134] <= 16'b0000_0000_0000_0000;
array[44135] <= 16'b0000_0000_0000_0000;
array[44136] <= 16'b0000_0000_0000_0000;
array[44137] <= 16'b0000_0000_0000_0000;
array[44138] <= 16'b0000_0000_0000_0000;
array[44139] <= 16'b0000_0000_0000_0000;
array[44140] <= 16'b0000_0000_0000_0000;
array[44141] <= 16'b0000_0000_0000_0000;
array[44142] <= 16'b0000_0000_0000_0000;
array[44143] <= 16'b0000_0000_0000_0000;
array[44144] <= 16'b0000_0000_0000_0000;
array[44145] <= 16'b0000_0000_0000_0000;
array[44146] <= 16'b0000_0000_0000_0000;
array[44147] <= 16'b0000_0000_0000_0000;
array[44148] <= 16'b0000_0000_0000_0000;
array[44149] <= 16'b0000_0000_0000_0000;
array[44150] <= 16'b0000_0000_0000_0000;
array[44151] <= 16'b0000_0000_0000_0000;
array[44152] <= 16'b0000_0000_0000_0000;
array[44153] <= 16'b0000_0000_0000_0000;
array[44154] <= 16'b0000_0000_0000_0000;
array[44155] <= 16'b0000_0000_0000_0000;
array[44156] <= 16'b0000_0000_0000_0000;
array[44157] <= 16'b0000_0000_0000_0000;
array[44158] <= 16'b0000_0000_0000_0000;
array[44159] <= 16'b0000_0000_0000_0000;
array[44160] <= 16'b0000_0000_0000_0000;
array[44161] <= 16'b0000_0000_0000_0000;
array[44162] <= 16'b0000_0000_0000_0000;
array[44163] <= 16'b0000_0000_0000_0000;
array[44164] <= 16'b0000_0000_0000_0000;
array[44165] <= 16'b0000_0000_0000_0000;
array[44166] <= 16'b0000_0000_0000_0000;
array[44167] <= 16'b0000_0000_0000_0000;
array[44168] <= 16'b0000_0000_0000_0000;
array[44169] <= 16'b0000_0000_0000_0000;
array[44170] <= 16'b0000_0000_0000_0000;
array[44171] <= 16'b0000_0000_0000_0000;
array[44172] <= 16'b0000_0000_0000_0000;
array[44173] <= 16'b0000_0000_0000_0000;
array[44174] <= 16'b0000_0000_0000_0000;
array[44175] <= 16'b0000_0000_0000_0000;
array[44176] <= 16'b0000_0000_0000_0000;
array[44177] <= 16'b0000_0000_0000_0000;
array[44178] <= 16'b0000_0000_0000_0000;
array[44179] <= 16'b0000_0000_0000_0000;
array[44180] <= 16'b0000_0000_0000_0000;
array[44181] <= 16'b0000_0000_0000_0000;
array[44182] <= 16'b0000_0000_0000_0000;
array[44183] <= 16'b0000_0000_0000_0000;
array[44184] <= 16'b0000_0000_0000_0000;
array[44185] <= 16'b0000_0000_0000_0000;
array[44186] <= 16'b0000_0000_0000_0000;
array[44187] <= 16'b0000_0000_0000_0000;
array[44188] <= 16'b0000_0000_0000_0000;
array[44189] <= 16'b0000_0000_0000_0000;
array[44190] <= 16'b0000_0000_0000_0000;
array[44191] <= 16'b0000_0000_0000_0000;
array[44192] <= 16'b0000_0000_0000_0000;
array[44193] <= 16'b0000_0000_0000_0000;
array[44194] <= 16'b0000_0000_0000_0000;
array[44195] <= 16'b0000_0000_0000_0000;
array[44196] <= 16'b0000_0000_0000_0000;
array[44197] <= 16'b0000_0000_0000_0000;
array[44198] <= 16'b0000_0000_0000_0000;
array[44199] <= 16'b0000_0000_0000_0000;
array[44200] <= 16'b0000_0000_0000_0000;
array[44201] <= 16'b0000_0000_0000_0000;
array[44202] <= 16'b0000_0000_0000_0000;
array[44203] <= 16'b0000_0000_0000_0000;
array[44204] <= 16'b0000_0000_0000_0000;
array[44205] <= 16'b0000_0000_0000_0000;
array[44206] <= 16'b0000_0000_0000_0000;
array[44207] <= 16'b0000_0000_0000_0000;
array[44208] <= 16'b0000_0000_0000_0000;
array[44209] <= 16'b0000_0000_0000_0000;
array[44210] <= 16'b0000_0000_0000_0000;
array[44211] <= 16'b0000_0000_0000_0000;
array[44212] <= 16'b0000_0000_0000_0000;
array[44213] <= 16'b0000_0000_0000_0000;
array[44214] <= 16'b0000_0000_0000_0000;
array[44215] <= 16'b0000_0000_0000_0000;
array[44216] <= 16'b0000_0000_0000_0000;
array[44217] <= 16'b0000_0000_0000_0000;
array[44218] <= 16'b0000_0000_0000_0000;
array[44219] <= 16'b0000_0000_0000_0000;
array[44220] <= 16'b0000_0000_0000_0000;
array[44221] <= 16'b0000_0000_0000_0000;
array[44222] <= 16'b0000_0000_0000_0000;
array[44223] <= 16'b0000_0000_0000_0000;
array[44224] <= 16'b0000_0000_0000_0000;
array[44225] <= 16'b0000_0000_0000_0000;
array[44226] <= 16'b0000_0000_0000_0000;
array[44227] <= 16'b0000_0000_0000_0000;
array[44228] <= 16'b0000_0000_0000_0000;
array[44229] <= 16'b0000_0000_0000_0000;
array[44230] <= 16'b0000_0000_0000_0000;
array[44231] <= 16'b0000_0000_0000_0000;
array[44232] <= 16'b0000_0000_0000_0000;
array[44233] <= 16'b0000_0000_0000_0000;
array[44234] <= 16'b0000_0000_0000_0000;
array[44235] <= 16'b0000_0000_0000_0000;
array[44236] <= 16'b0000_0000_0000_0000;
array[44237] <= 16'b0000_0000_0000_0000;
array[44238] <= 16'b0000_0000_0000_0000;
array[44239] <= 16'b0000_0000_0000_0000;
array[44240] <= 16'b0000_0000_0000_0000;
array[44241] <= 16'b0000_0000_0000_0000;
array[44242] <= 16'b0000_0000_0000_0000;
array[44243] <= 16'b0000_0000_0000_0000;
array[44244] <= 16'b0000_0000_0000_0000;
array[44245] <= 16'b0000_0000_0000_0000;
array[44246] <= 16'b0000_0000_0000_0000;
array[44247] <= 16'b0000_0000_0000_0000;
array[44248] <= 16'b0000_0000_0000_0000;
array[44249] <= 16'b0000_0000_0000_0000;
array[44250] <= 16'b0000_0000_0000_0000;
array[44251] <= 16'b0000_0000_0000_0000;
array[44252] <= 16'b0000_0000_0000_0000;
array[44253] <= 16'b0000_0000_0000_0000;
array[44254] <= 16'b0000_0000_0000_0000;
array[44255] <= 16'b0000_0000_0000_0000;
array[44256] <= 16'b0000_0000_0000_0000;
array[44257] <= 16'b0000_0000_0000_0000;
array[44258] <= 16'b0000_0000_0000_0000;
array[44259] <= 16'b0000_0000_0000_0000;
array[44260] <= 16'b0000_0000_0000_0000;
array[44261] <= 16'b0000_0000_0000_0000;
array[44262] <= 16'b0000_0000_0000_0000;
array[44263] <= 16'b0000_0000_0000_0000;
array[44264] <= 16'b0000_0000_0000_0000;
array[44265] <= 16'b0000_0000_0000_0000;
array[44266] <= 16'b0000_0000_0000_0000;
array[44267] <= 16'b0000_0000_0000_0000;
array[44268] <= 16'b0000_0000_0000_0000;
array[44269] <= 16'b0000_0000_0000_0000;
array[44270] <= 16'b0000_0000_0000_0000;
array[44271] <= 16'b0000_0000_0000_0000;
array[44272] <= 16'b0000_0000_0000_0000;
array[44273] <= 16'b0000_0000_0000_0000;
array[44274] <= 16'b0000_0000_0000_0000;
array[44275] <= 16'b0000_0000_0000_0000;
array[44276] <= 16'b0000_0000_0000_0000;
array[44277] <= 16'b0000_0000_0000_0000;
array[44278] <= 16'b0000_0000_0000_0000;
array[44279] <= 16'b0000_0000_0000_0000;
array[44280] <= 16'b0000_0000_0000_0000;
array[44281] <= 16'b0000_0000_0000_0000;
array[44282] <= 16'b0000_0000_0000_0000;
array[44283] <= 16'b0000_0000_0000_0000;
array[44284] <= 16'b0000_0000_0000_0000;
array[44285] <= 16'b0000_0000_0000_0000;
array[44286] <= 16'b0000_0000_0000_0000;
array[44287] <= 16'b0000_0000_0000_0000;
array[44288] <= 16'b0000_0000_0000_0000;
array[44289] <= 16'b0000_0000_0000_0000;
array[44290] <= 16'b0000_0000_0000_0000;
array[44291] <= 16'b0000_0000_0000_0000;
array[44292] <= 16'b0000_0000_0000_0000;
array[44293] <= 16'b0000_0000_0000_0000;
array[44294] <= 16'b0000_0000_0000_0000;
array[44295] <= 16'b0000_0000_0000_0000;
array[44296] <= 16'b0000_0000_0000_0000;
array[44297] <= 16'b0000_0000_0000_0000;
array[44298] <= 16'b0000_0000_0000_0000;
array[44299] <= 16'b0000_0000_0000_0000;
array[44300] <= 16'b0000_0000_0000_0000;
array[44301] <= 16'b0000_0000_0000_0000;
array[44302] <= 16'b0000_0000_0000_0000;
array[44303] <= 16'b0000_0000_0000_0000;
array[44304] <= 16'b0000_0000_0000_0000;
array[44305] <= 16'b0000_0000_0000_0000;
array[44306] <= 16'b0000_0000_0000_0000;
array[44307] <= 16'b0000_0000_0000_0000;
array[44308] <= 16'b0000_0000_0000_0000;
array[44309] <= 16'b0000_0000_0000_0000;
array[44310] <= 16'b0000_0000_0000_0000;
array[44311] <= 16'b0000_0000_0000_0000;
array[44312] <= 16'b0000_0000_0000_0000;
array[44313] <= 16'b0000_0000_0000_0000;
array[44314] <= 16'b0000_0000_0000_0000;
array[44315] <= 16'b0000_0000_0000_0000;
array[44316] <= 16'b0000_0000_0000_0000;
array[44317] <= 16'b0000_0000_0000_0000;
array[44318] <= 16'b0000_0000_0000_0000;
array[44319] <= 16'b0000_0000_0000_0000;
array[44320] <= 16'b0000_0000_0000_0000;
array[44321] <= 16'b0000_0000_0000_0000;
array[44322] <= 16'b0000_0000_0000_0000;
array[44323] <= 16'b0000_0000_0000_0000;
array[44324] <= 16'b0000_0000_0000_0000;
array[44325] <= 16'b0000_0000_0000_0000;
array[44326] <= 16'b0000_0000_0000_0000;
array[44327] <= 16'b0000_0000_0000_0000;
array[44328] <= 16'b0000_0000_0000_0000;
array[44329] <= 16'b0000_0000_0000_0000;
array[44330] <= 16'b0000_0000_0000_0000;
array[44331] <= 16'b0000_0000_0000_0000;
array[44332] <= 16'b0000_0000_0000_0000;
array[44333] <= 16'b0000_0000_0000_0000;
array[44334] <= 16'b0000_0000_0000_0000;
array[44335] <= 16'b0000_0000_0000_0000;
array[44336] <= 16'b0000_0000_0000_0000;
array[44337] <= 16'b0000_0000_0000_0000;
array[44338] <= 16'b0000_0000_0000_0000;
array[44339] <= 16'b0000_0000_0000_0000;
array[44340] <= 16'b0000_0000_0000_0000;
array[44341] <= 16'b0000_0000_0000_0000;
array[44342] <= 16'b0000_0000_0000_0000;
array[44343] <= 16'b0000_0000_0000_0000;
array[44344] <= 16'b0000_0000_0000_0000;
array[44345] <= 16'b0000_0000_0000_0000;
array[44346] <= 16'b0000_0000_0000_0000;
array[44347] <= 16'b0000_0000_0000_0000;
array[44348] <= 16'b0000_0000_0000_0000;
array[44349] <= 16'b0000_0000_0000_0000;
array[44350] <= 16'b0000_0000_0000_0000;
array[44351] <= 16'b0000_0000_0000_0000;
array[44352] <= 16'b0000_0000_0000_0000;
array[44353] <= 16'b0000_0000_0000_0000;
array[44354] <= 16'b0000_0000_0000_0000;
array[44355] <= 16'b0000_0000_0000_0000;
array[44356] <= 16'b0000_0000_0000_0000;
array[44357] <= 16'b0000_0000_0000_0000;
array[44358] <= 16'b0000_0000_0000_0000;
array[44359] <= 16'b0000_0000_0000_0000;
array[44360] <= 16'b0000_0000_0000_0000;
array[44361] <= 16'b0000_0000_0000_0000;
array[44362] <= 16'b0000_0000_0000_0000;
array[44363] <= 16'b0000_0000_0000_0000;
array[44364] <= 16'b0000_0000_0000_0000;
array[44365] <= 16'b0000_0000_0000_0000;
array[44366] <= 16'b0000_0000_0000_0000;
array[44367] <= 16'b0000_0000_0000_0000;
array[44368] <= 16'b0000_0000_0000_0000;
array[44369] <= 16'b0000_0000_0000_0000;
array[44370] <= 16'b0000_0000_0000_0000;
array[44371] <= 16'b0000_0000_0000_0000;
array[44372] <= 16'b0000_0000_0000_0000;
array[44373] <= 16'b0000_0000_0000_0000;
array[44374] <= 16'b0000_0000_0000_0000;
array[44375] <= 16'b0000_0000_0000_0000;
array[44376] <= 16'b0000_0000_0000_0000;
array[44377] <= 16'b0000_0000_0000_0000;
array[44378] <= 16'b0000_0000_0000_0000;
array[44379] <= 16'b0000_0000_0000_0000;
array[44380] <= 16'b0000_0000_0000_0000;
array[44381] <= 16'b0000_0000_0000_0000;
array[44382] <= 16'b0000_0000_0000_0000;
array[44383] <= 16'b0000_0000_0000_0000;
array[44384] <= 16'b0000_0000_0000_0000;
array[44385] <= 16'b0000_0000_0000_0000;
array[44386] <= 16'b0000_0000_0000_0000;
array[44387] <= 16'b0000_0000_0000_0000;
array[44388] <= 16'b0000_0000_0000_0000;
array[44389] <= 16'b0000_0000_0000_0000;
array[44390] <= 16'b0000_0000_0000_0000;
array[44391] <= 16'b0000_0000_0000_0000;
array[44392] <= 16'b0000_0000_0000_0000;
array[44393] <= 16'b0000_0000_0000_0000;
array[44394] <= 16'b0000_0000_0000_0000;
array[44395] <= 16'b0000_0000_0000_0000;
array[44396] <= 16'b0000_0000_0000_0000;
array[44397] <= 16'b0000_0000_0000_0000;
array[44398] <= 16'b0000_0000_0000_0000;
array[44399] <= 16'b0000_0000_0000_0000;
array[44400] <= 16'b0000_0000_0000_0000;
array[44401] <= 16'b0000_0000_0000_0000;
array[44402] <= 16'b0000_0000_0000_0000;
array[44403] <= 16'b0000_0000_0000_0000;
array[44404] <= 16'b0000_0000_0000_0000;
array[44405] <= 16'b0000_0000_0000_0000;
array[44406] <= 16'b0000_0000_0000_0000;
array[44407] <= 16'b0000_0000_0000_0000;
array[44408] <= 16'b0000_0000_0000_0000;
array[44409] <= 16'b0000_0000_0000_0000;
array[44410] <= 16'b0000_0000_0000_0000;
array[44411] <= 16'b0000_0000_0000_0000;
array[44412] <= 16'b0000_0000_0000_0000;
array[44413] <= 16'b0000_0000_0000_0000;
array[44414] <= 16'b0000_0000_0000_0000;
array[44415] <= 16'b0000_0000_0000_0000;
array[44416] <= 16'b0000_0000_0000_0000;
array[44417] <= 16'b0000_0000_0000_0000;
array[44418] <= 16'b0000_0000_0000_0000;
array[44419] <= 16'b0000_0000_0000_0000;
array[44420] <= 16'b0000_0000_0000_0000;
array[44421] <= 16'b0000_0000_0000_0000;
array[44422] <= 16'b0000_0000_0000_0000;
array[44423] <= 16'b0000_0000_0000_0000;
array[44424] <= 16'b0000_0000_0000_0000;
array[44425] <= 16'b0000_0000_0000_0000;
array[44426] <= 16'b0000_0000_0000_0000;
array[44427] <= 16'b0000_0000_0000_0000;
array[44428] <= 16'b0000_0000_0000_0000;
array[44429] <= 16'b0000_0000_0000_0000;
array[44430] <= 16'b0000_0000_0000_0000;
array[44431] <= 16'b0000_0000_0000_0000;
array[44432] <= 16'b0000_0000_0000_0000;
array[44433] <= 16'b0000_0000_0000_0000;
array[44434] <= 16'b0000_0000_0000_0000;
array[44435] <= 16'b0000_0000_0000_0000;
array[44436] <= 16'b0000_0000_0000_0000;
array[44437] <= 16'b0000_0000_0000_0000;
array[44438] <= 16'b0000_0000_0000_0000;
array[44439] <= 16'b0000_0000_0000_0000;
array[44440] <= 16'b0000_0000_0000_0000;
array[44441] <= 16'b0000_0000_0000_0000;
array[44442] <= 16'b0000_0000_0000_0000;
array[44443] <= 16'b0000_0000_0000_0000;
array[44444] <= 16'b0000_0000_0000_0000;
array[44445] <= 16'b0000_0000_0000_0000;
array[44446] <= 16'b0000_0000_0000_0000;
array[44447] <= 16'b0000_0000_0000_0000;
array[44448] <= 16'b0000_0000_0000_0000;
array[44449] <= 16'b0000_0000_0000_0000;
array[44450] <= 16'b0000_0000_0000_0000;
array[44451] <= 16'b0000_0000_0000_0000;
array[44452] <= 16'b0000_0000_0000_0000;
array[44453] <= 16'b0000_0000_0000_0000;
array[44454] <= 16'b0000_0000_0000_0000;
array[44455] <= 16'b0000_0000_0000_0000;
array[44456] <= 16'b0000_0000_0000_0000;
array[44457] <= 16'b0000_0000_0000_0000;
array[44458] <= 16'b0000_0000_0000_0000;
array[44459] <= 16'b0000_0000_0000_0000;
array[44460] <= 16'b0000_0000_0000_0000;
array[44461] <= 16'b0000_0000_0000_0000;
array[44462] <= 16'b0000_0000_0000_0000;
array[44463] <= 16'b0000_0000_0000_0000;
array[44464] <= 16'b0000_0000_0000_0000;
array[44465] <= 16'b0000_0000_0000_0000;
array[44466] <= 16'b0000_0000_0000_0000;
array[44467] <= 16'b0000_0000_0000_0000;
array[44468] <= 16'b0000_0000_0000_0000;
array[44469] <= 16'b0000_0000_0000_0000;
array[44470] <= 16'b0000_0000_0000_0000;
array[44471] <= 16'b0000_0000_0000_0000;
array[44472] <= 16'b0000_0000_0000_0000;
array[44473] <= 16'b0000_0000_0000_0000;
array[44474] <= 16'b0000_0000_0000_0000;
array[44475] <= 16'b0000_0000_0000_0000;
array[44476] <= 16'b0000_0000_0000_0000;
array[44477] <= 16'b0000_0000_0000_0000;
array[44478] <= 16'b0000_0000_0000_0000;
array[44479] <= 16'b0000_0000_0000_0000;
array[44480] <= 16'b0000_0000_0000_0000;
array[44481] <= 16'b0000_0000_0000_0000;
array[44482] <= 16'b0000_0000_0000_0000;
array[44483] <= 16'b0000_0000_0000_0000;
array[44484] <= 16'b0000_0000_0000_0000;
array[44485] <= 16'b0000_0000_0000_0000;
array[44486] <= 16'b0000_0000_0000_0000;
array[44487] <= 16'b0000_0000_0000_0000;
array[44488] <= 16'b0000_0000_0000_0000;
array[44489] <= 16'b0000_0000_0000_0000;
array[44490] <= 16'b0000_0000_0000_0000;
array[44491] <= 16'b0000_0000_0000_0000;
array[44492] <= 16'b0000_0000_0000_0000;
array[44493] <= 16'b0000_0000_0000_0000;
array[44494] <= 16'b0000_0000_0000_0000;
array[44495] <= 16'b0000_0000_0000_0000;
array[44496] <= 16'b0000_0000_0000_0000;
array[44497] <= 16'b0000_0000_0000_0000;
array[44498] <= 16'b0000_0000_0000_0000;
array[44499] <= 16'b0000_0000_0000_0000;
array[44500] <= 16'b0000_0000_0000_0000;
array[44501] <= 16'b0000_0000_0000_0000;
array[44502] <= 16'b0000_0000_0000_0000;
array[44503] <= 16'b0000_0000_0000_0000;
array[44504] <= 16'b0000_0000_0000_0000;
array[44505] <= 16'b0000_0000_0000_0000;
array[44506] <= 16'b0000_0000_0000_0000;
array[44507] <= 16'b0000_0000_0000_0000;
array[44508] <= 16'b0000_0000_0000_0000;
array[44509] <= 16'b0000_0000_0000_0000;
array[44510] <= 16'b0000_0000_0000_0000;
array[44511] <= 16'b0000_0000_0000_0000;
array[44512] <= 16'b0000_0000_0000_0000;
array[44513] <= 16'b0000_0000_0000_0000;
array[44514] <= 16'b0000_0000_0000_0000;
array[44515] <= 16'b0000_0000_0000_0000;
array[44516] <= 16'b0000_0000_0000_0000;
array[44517] <= 16'b0000_0000_0000_0000;
array[44518] <= 16'b0000_0000_0000_0000;
array[44519] <= 16'b0000_0000_0000_0000;
array[44520] <= 16'b0000_0000_0000_0000;
array[44521] <= 16'b0000_0000_0000_0000;
array[44522] <= 16'b0000_0000_0000_0000;
array[44523] <= 16'b0000_0000_0000_0000;
array[44524] <= 16'b0000_0000_0000_0000;
array[44525] <= 16'b0000_0000_0000_0000;
array[44526] <= 16'b0000_0000_0000_0000;
array[44527] <= 16'b0000_0000_0000_0000;
array[44528] <= 16'b0000_0000_0000_0000;
array[44529] <= 16'b0000_0000_0000_0000;
array[44530] <= 16'b0000_0000_0000_0000;
array[44531] <= 16'b0000_0000_0000_0000;
array[44532] <= 16'b0000_0000_0000_0000;
array[44533] <= 16'b0000_0000_0000_0000;
array[44534] <= 16'b0000_0000_0000_0000;
array[44535] <= 16'b0000_0000_0000_0000;
array[44536] <= 16'b0000_0000_0000_0000;
array[44537] <= 16'b0000_0000_0000_0000;
array[44538] <= 16'b0000_0000_0000_0000;
array[44539] <= 16'b0000_0000_0000_0000;
array[44540] <= 16'b0000_0000_0000_0000;
array[44541] <= 16'b0000_0000_0000_0000;
array[44542] <= 16'b0000_0000_0000_0000;
array[44543] <= 16'b0000_0000_0000_0000;
array[44544] <= 16'b0000_0000_0000_0000;
array[44545] <= 16'b0000_0000_0000_0000;
array[44546] <= 16'b0000_0000_0000_0000;
array[44547] <= 16'b0000_0000_0000_0000;
array[44548] <= 16'b0000_0000_0000_0000;
array[44549] <= 16'b0000_0000_0000_0000;
array[44550] <= 16'b0000_0000_0000_0000;
array[44551] <= 16'b0000_0000_0000_0000;
array[44552] <= 16'b0000_0000_0000_0000;
array[44553] <= 16'b0000_0000_0000_0000;
array[44554] <= 16'b0000_0000_0000_0000;
array[44555] <= 16'b0000_0000_0000_0000;
array[44556] <= 16'b0000_0000_0000_0000;
array[44557] <= 16'b0000_0000_0000_0000;
array[44558] <= 16'b0000_0000_0000_0000;
array[44559] <= 16'b0000_0000_0000_0000;
array[44560] <= 16'b0000_0000_0000_0000;
array[44561] <= 16'b0000_0000_0000_0000;
array[44562] <= 16'b0000_0000_0000_0000;
array[44563] <= 16'b0000_0000_0000_0000;
array[44564] <= 16'b0000_0000_0000_0000;
array[44565] <= 16'b0000_0000_0000_0000;
array[44566] <= 16'b0000_0000_0000_0000;
array[44567] <= 16'b0000_0000_0000_0000;
array[44568] <= 16'b0000_0000_0000_0000;
array[44569] <= 16'b0000_0000_0000_0000;
array[44570] <= 16'b0000_0000_0000_0000;
array[44571] <= 16'b0000_0000_0000_0000;
array[44572] <= 16'b0000_0000_0000_0000;
array[44573] <= 16'b0000_0000_0000_0000;
array[44574] <= 16'b0000_0000_0000_0000;
array[44575] <= 16'b0000_0000_0000_0000;
array[44576] <= 16'b0000_0000_0000_0000;
array[44577] <= 16'b0000_0000_0000_0000;
array[44578] <= 16'b0000_0000_0000_0000;
array[44579] <= 16'b0000_0000_0000_0000;
array[44580] <= 16'b0000_0000_0000_0000;
array[44581] <= 16'b0000_0000_0000_0000;
array[44582] <= 16'b0000_0000_0000_0000;
array[44583] <= 16'b0000_0000_0000_0000;
array[44584] <= 16'b0000_0000_0000_0000;
array[44585] <= 16'b0000_0000_0000_0000;
array[44586] <= 16'b0000_0000_0000_0000;
array[44587] <= 16'b0000_0000_0000_0000;
array[44588] <= 16'b0000_0000_0000_0000;
array[44589] <= 16'b0000_0000_0000_0000;
array[44590] <= 16'b0000_0000_0000_0000;
array[44591] <= 16'b0000_0000_0000_0000;
array[44592] <= 16'b0000_0000_0000_0000;
array[44593] <= 16'b0000_0000_0000_0000;
array[44594] <= 16'b0000_0000_0000_0000;
array[44595] <= 16'b0000_0000_0000_0000;
array[44596] <= 16'b0000_0000_0000_0000;
array[44597] <= 16'b0000_0000_0000_0000;
array[44598] <= 16'b0000_0000_0000_0000;
array[44599] <= 16'b0000_0000_0000_0000;
array[44600] <= 16'b0000_0000_0000_0000;
array[44601] <= 16'b0000_0000_0000_0000;
array[44602] <= 16'b0000_0000_0000_0000;
array[44603] <= 16'b0000_0000_0000_0000;
array[44604] <= 16'b0000_0000_0000_0000;
array[44605] <= 16'b0000_0000_0000_0000;
array[44606] <= 16'b0000_0000_0000_0000;
array[44607] <= 16'b0000_0000_0000_0000;
array[44608] <= 16'b0000_0000_0000_0000;
array[44609] <= 16'b0000_0000_0000_0000;
array[44610] <= 16'b0000_0000_0000_0000;
array[44611] <= 16'b0000_0000_0000_0000;
array[44612] <= 16'b0000_0000_0000_0000;
array[44613] <= 16'b0000_0000_0000_0000;
array[44614] <= 16'b0000_0000_0000_0000;
array[44615] <= 16'b0000_0000_0000_0000;
array[44616] <= 16'b0000_0000_0000_0000;
array[44617] <= 16'b0000_0000_0000_0000;
array[44618] <= 16'b0000_0000_0000_0000;
array[44619] <= 16'b0000_0000_0000_0000;
array[44620] <= 16'b0000_0000_0000_0000;
array[44621] <= 16'b0000_0000_0000_0000;
array[44622] <= 16'b0000_0000_0000_0000;
array[44623] <= 16'b0000_0000_0000_0000;
array[44624] <= 16'b0000_0000_0000_0000;
array[44625] <= 16'b0000_0000_0000_0000;
array[44626] <= 16'b0000_0000_0000_0000;
array[44627] <= 16'b0000_0000_0000_0000;
array[44628] <= 16'b0000_0000_0000_0000;
array[44629] <= 16'b0000_0000_0000_0000;
array[44630] <= 16'b0000_0000_0000_0000;
array[44631] <= 16'b0000_0000_0000_0000;
array[44632] <= 16'b0000_0000_0000_0000;
array[44633] <= 16'b0000_0000_0000_0000;
array[44634] <= 16'b0000_0000_0000_0000;
array[44635] <= 16'b0000_0000_0000_0000;
array[44636] <= 16'b0000_0000_0000_0000;
array[44637] <= 16'b0000_0000_0000_0000;
array[44638] <= 16'b0000_0000_0000_0000;
array[44639] <= 16'b0000_0000_0000_0000;
array[44640] <= 16'b0000_0000_0000_0000;
array[44641] <= 16'b0000_0000_0000_0000;
array[44642] <= 16'b0000_0000_0000_0000;
array[44643] <= 16'b0000_0000_0000_0000;
array[44644] <= 16'b0000_0000_0000_0000;
array[44645] <= 16'b0000_0000_0000_0000;
array[44646] <= 16'b0000_0000_0000_0000;
array[44647] <= 16'b0000_0000_0000_0000;
array[44648] <= 16'b0000_0000_0000_0000;
array[44649] <= 16'b0000_0000_0000_0000;
array[44650] <= 16'b0000_0000_0000_0000;
array[44651] <= 16'b0000_0000_0000_0000;
array[44652] <= 16'b0000_0000_0000_0000;
array[44653] <= 16'b0000_0000_0000_0000;
array[44654] <= 16'b0000_0000_0000_0000;
array[44655] <= 16'b0000_0000_0000_0000;
array[44656] <= 16'b0000_0000_0000_0000;
array[44657] <= 16'b0000_0000_0000_0000;
array[44658] <= 16'b0000_0000_0000_0000;
array[44659] <= 16'b0000_0000_0000_0000;
array[44660] <= 16'b0000_0000_0000_0000;
array[44661] <= 16'b0000_0000_0000_0000;
array[44662] <= 16'b0000_0000_0000_0000;
array[44663] <= 16'b0000_0000_0000_0000;
array[44664] <= 16'b0000_0000_0000_0000;
array[44665] <= 16'b0000_0000_0000_0000;
array[44666] <= 16'b0000_0000_0000_0000;
array[44667] <= 16'b0000_0000_0000_0000;
array[44668] <= 16'b0000_0000_0000_0000;
array[44669] <= 16'b0000_0000_0000_0000;
array[44670] <= 16'b0000_0000_0000_0000;
array[44671] <= 16'b0000_0000_0000_0000;
array[44672] <= 16'b0000_0000_0000_0000;
array[44673] <= 16'b0000_0000_0000_0000;
array[44674] <= 16'b0000_0000_0000_0000;
array[44675] <= 16'b0000_0000_0000_0000;
array[44676] <= 16'b0000_0000_0000_0000;
array[44677] <= 16'b0000_0000_0000_0000;
array[44678] <= 16'b0000_0000_0000_0000;
array[44679] <= 16'b0000_0000_0000_0000;
array[44680] <= 16'b0000_0000_0000_0000;
array[44681] <= 16'b0000_0000_0000_0000;
array[44682] <= 16'b0000_0000_0000_0000;
array[44683] <= 16'b0000_0000_0000_0000;
array[44684] <= 16'b0000_0000_0000_0000;
array[44685] <= 16'b0000_0000_0000_0000;
array[44686] <= 16'b0000_0000_0000_0000;
array[44687] <= 16'b0000_0000_0000_0000;
array[44688] <= 16'b0000_0000_0000_0000;
array[44689] <= 16'b0000_0000_0000_0000;
array[44690] <= 16'b0000_0000_0000_0000;
array[44691] <= 16'b0000_0000_0000_0000;
array[44692] <= 16'b0000_0000_0000_0000;
array[44693] <= 16'b0000_0000_0000_0000;
array[44694] <= 16'b0000_0000_0000_0000;
array[44695] <= 16'b0000_0000_0000_0000;
array[44696] <= 16'b0000_0000_0000_0000;
array[44697] <= 16'b0000_0000_0000_0000;
array[44698] <= 16'b0000_0000_0000_0000;
array[44699] <= 16'b0000_0000_0000_0000;
array[44700] <= 16'b0000_0000_0000_0000;
array[44701] <= 16'b0000_0000_0000_0000;
array[44702] <= 16'b0000_0000_0000_0000;
array[44703] <= 16'b0000_0000_0000_0000;
array[44704] <= 16'b0000_0000_0000_0000;
array[44705] <= 16'b0000_0000_0000_0000;
array[44706] <= 16'b0000_0000_0000_0000;
array[44707] <= 16'b0000_0000_0000_0000;
array[44708] <= 16'b0000_0000_0000_0000;
array[44709] <= 16'b0000_0000_0000_0000;
array[44710] <= 16'b0000_0000_0000_0000;
array[44711] <= 16'b0000_0000_0000_0000;
array[44712] <= 16'b0000_0000_0000_0000;
array[44713] <= 16'b0000_0000_0000_0000;
array[44714] <= 16'b0000_0000_0000_0000;
array[44715] <= 16'b0000_0000_0000_0000;
array[44716] <= 16'b0000_0000_0000_0000;
array[44717] <= 16'b0000_0000_0000_0000;
array[44718] <= 16'b0000_0000_0000_0000;
array[44719] <= 16'b0000_0000_0000_0000;
array[44720] <= 16'b0000_0000_0000_0000;
array[44721] <= 16'b0000_0000_0000_0000;
array[44722] <= 16'b0000_0000_0000_0000;
array[44723] <= 16'b0000_0000_0000_0000;
array[44724] <= 16'b0000_0000_0000_0000;
array[44725] <= 16'b0000_0000_0000_0000;
array[44726] <= 16'b0000_0000_0000_0000;
array[44727] <= 16'b0000_0000_0000_0000;
array[44728] <= 16'b0000_0000_0000_0000;
array[44729] <= 16'b0000_0000_0000_0000;
array[44730] <= 16'b0000_0000_0000_0000;
array[44731] <= 16'b0000_0000_0000_0000;
array[44732] <= 16'b0000_0000_0000_0000;
array[44733] <= 16'b0000_0000_0000_0000;
array[44734] <= 16'b0000_0000_0000_0000;
array[44735] <= 16'b0000_0000_0000_0000;
array[44736] <= 16'b0000_0000_0000_0000;
array[44737] <= 16'b0000_0000_0000_0000;
array[44738] <= 16'b0000_0000_0000_0000;
array[44739] <= 16'b0000_0000_0000_0000;
array[44740] <= 16'b0000_0000_0000_0000;
array[44741] <= 16'b0000_0000_0000_0000;
array[44742] <= 16'b0000_0000_0000_0000;
array[44743] <= 16'b0000_0000_0000_0000;
array[44744] <= 16'b0000_0000_0000_0000;
array[44745] <= 16'b0000_0000_0000_0000;
array[44746] <= 16'b0000_0000_0000_0000;
array[44747] <= 16'b0000_0000_0000_0000;
array[44748] <= 16'b0000_0000_0000_0000;
array[44749] <= 16'b0000_0000_0000_0000;
array[44750] <= 16'b0000_0000_0000_0000;
array[44751] <= 16'b0000_0000_0000_0000;
array[44752] <= 16'b0000_0000_0000_0000;
array[44753] <= 16'b0000_0000_0000_0000;
array[44754] <= 16'b0000_0000_0000_0000;
array[44755] <= 16'b0000_0000_0000_0000;
array[44756] <= 16'b0000_0000_0000_0000;
array[44757] <= 16'b0000_0000_0000_0000;
array[44758] <= 16'b0000_0000_0000_0000;
array[44759] <= 16'b0000_0000_0000_0000;
array[44760] <= 16'b0000_0000_0000_0000;
array[44761] <= 16'b0000_0000_0000_0000;
array[44762] <= 16'b0000_0000_0000_0000;
array[44763] <= 16'b0000_0000_0000_0000;
array[44764] <= 16'b0000_0000_0000_0000;
array[44765] <= 16'b0000_0000_0000_0000;
array[44766] <= 16'b0000_0000_0000_0000;
array[44767] <= 16'b0000_0000_0000_0000;
array[44768] <= 16'b0000_0000_0000_0000;
array[44769] <= 16'b0000_0000_0000_0000;
array[44770] <= 16'b0000_0000_0000_0000;
array[44771] <= 16'b0000_0000_0000_0000;
array[44772] <= 16'b0000_0000_0000_0000;
array[44773] <= 16'b0000_0000_0000_0000;
array[44774] <= 16'b0000_0000_0000_0000;
array[44775] <= 16'b0000_0000_0000_0000;
array[44776] <= 16'b0000_0000_0000_0000;
array[44777] <= 16'b0000_0000_0000_0000;
array[44778] <= 16'b0000_0000_0000_0000;
array[44779] <= 16'b0000_0000_0000_0000;
array[44780] <= 16'b0000_0000_0000_0000;
array[44781] <= 16'b0000_0000_0000_0000;
array[44782] <= 16'b0000_0000_0000_0000;
array[44783] <= 16'b0000_0000_0000_0000;
array[44784] <= 16'b0000_0000_0000_0000;
array[44785] <= 16'b0000_0000_0000_0000;
array[44786] <= 16'b0000_0000_0000_0000;
array[44787] <= 16'b0000_0000_0000_0000;
array[44788] <= 16'b0000_0000_0000_0000;
array[44789] <= 16'b0000_0000_0000_0000;
array[44790] <= 16'b0000_0000_0000_0000;
array[44791] <= 16'b0000_0000_0000_0000;
array[44792] <= 16'b0000_0000_0000_0000;
array[44793] <= 16'b0000_0000_0000_0000;
array[44794] <= 16'b0000_0000_0000_0000;
array[44795] <= 16'b0000_0000_0000_0000;
array[44796] <= 16'b0000_0000_0000_0000;
array[44797] <= 16'b0000_0000_0000_0000;
array[44798] <= 16'b0000_0000_0000_0000;
array[44799] <= 16'b0000_0000_0000_0000;
array[44800] <= 16'b0000_0000_0000_0000;
array[44801] <= 16'b0000_0000_0000_0000;
array[44802] <= 16'b0000_0000_0000_0000;
array[44803] <= 16'b0000_0000_0000_0000;
array[44804] <= 16'b0000_0000_0000_0000;
array[44805] <= 16'b0000_0000_0000_0000;
array[44806] <= 16'b0000_0000_0000_0000;
array[44807] <= 16'b0000_0000_0000_0000;
array[44808] <= 16'b0000_0000_0000_0000;
array[44809] <= 16'b0000_0000_0000_0000;
array[44810] <= 16'b0000_0000_0000_0000;
array[44811] <= 16'b0000_0000_0000_0000;
array[44812] <= 16'b0000_0000_0000_0000;
array[44813] <= 16'b0000_0000_0000_0000;
array[44814] <= 16'b0000_0000_0000_0000;
array[44815] <= 16'b0000_0000_0000_0000;
array[44816] <= 16'b0000_0000_0000_0000;
array[44817] <= 16'b0000_0000_0000_0000;
array[44818] <= 16'b0000_0000_0000_0000;
array[44819] <= 16'b0000_0000_0000_0000;
array[44820] <= 16'b0000_0000_0000_0000;
array[44821] <= 16'b0000_0000_0000_0000;
array[44822] <= 16'b0000_0000_0000_0000;
array[44823] <= 16'b0000_0000_0000_0000;
array[44824] <= 16'b0000_0000_0000_0000;
array[44825] <= 16'b0000_0000_0000_0000;
array[44826] <= 16'b0000_0000_0000_0000;
array[44827] <= 16'b0000_0000_0000_0000;
array[44828] <= 16'b0000_0000_0000_0000;
array[44829] <= 16'b0000_0000_0000_0000;
array[44830] <= 16'b0000_0000_0000_0000;
array[44831] <= 16'b0000_0000_0000_0000;
array[44832] <= 16'b0000_0000_0000_0000;
array[44833] <= 16'b0000_0000_0000_0000;
array[44834] <= 16'b0000_0000_0000_0000;
array[44835] <= 16'b0000_0000_0000_0000;
array[44836] <= 16'b0000_0000_0000_0000;
array[44837] <= 16'b0000_0000_0000_0000;
array[44838] <= 16'b0000_0000_0000_0000;
array[44839] <= 16'b0000_0000_0000_0000;
array[44840] <= 16'b0000_0000_0000_0000;
array[44841] <= 16'b0000_0000_0000_0000;
array[44842] <= 16'b0000_0000_0000_0000;
array[44843] <= 16'b0000_0000_0000_0000;
array[44844] <= 16'b0000_0000_0000_0000;
array[44845] <= 16'b0000_0000_0000_0000;
array[44846] <= 16'b0000_0000_0000_0000;
array[44847] <= 16'b0000_0000_0000_0000;
array[44848] <= 16'b0000_0000_0000_0000;
array[44849] <= 16'b0000_0000_0000_0000;
array[44850] <= 16'b0000_0000_0000_0000;
array[44851] <= 16'b0000_0000_0000_0000;
array[44852] <= 16'b0000_0000_0000_0000;
array[44853] <= 16'b0000_0000_0000_0000;
array[44854] <= 16'b0000_0000_0000_0000;
array[44855] <= 16'b0000_0000_0000_0000;
array[44856] <= 16'b0000_0000_0000_0000;
array[44857] <= 16'b0000_0000_0000_0000;
array[44858] <= 16'b0000_0000_0000_0000;
array[44859] <= 16'b0000_0000_0000_0000;
array[44860] <= 16'b0000_0000_0000_0000;
array[44861] <= 16'b0000_0000_0000_0000;
array[44862] <= 16'b0000_0000_0000_0000;
array[44863] <= 16'b0000_0000_0000_0000;
array[44864] <= 16'b0000_0000_0000_0000;
array[44865] <= 16'b0000_0000_0000_0000;
array[44866] <= 16'b0000_0000_0000_0000;
array[44867] <= 16'b0000_0000_0000_0000;
array[44868] <= 16'b0000_0000_0000_0000;
array[44869] <= 16'b0000_0000_0000_0000;
array[44870] <= 16'b0000_0000_0000_0000;
array[44871] <= 16'b0000_0000_0000_0000;
array[44872] <= 16'b0000_0000_0000_0000;
array[44873] <= 16'b0000_0000_0000_0000;
array[44874] <= 16'b0000_0000_0000_0000;
array[44875] <= 16'b0000_0000_0000_0000;
array[44876] <= 16'b0000_0000_0000_0000;
array[44877] <= 16'b0000_0000_0000_0000;
array[44878] <= 16'b0000_0000_0000_0000;
array[44879] <= 16'b0000_0000_0000_0000;
array[44880] <= 16'b0000_0000_0000_0000;
array[44881] <= 16'b0000_0000_0000_0000;
array[44882] <= 16'b0000_0000_0000_0000;
array[44883] <= 16'b0000_0000_0000_0000;
array[44884] <= 16'b0000_0000_0000_0000;
array[44885] <= 16'b0000_0000_0000_0000;
array[44886] <= 16'b0000_0000_0000_0000;
array[44887] <= 16'b0000_0000_0000_0000;
array[44888] <= 16'b0000_0000_0000_0000;
array[44889] <= 16'b0000_0000_0000_0000;
array[44890] <= 16'b0000_0000_0000_0000;
array[44891] <= 16'b0000_0000_0000_0000;
array[44892] <= 16'b0000_0000_0000_0000;
array[44893] <= 16'b0000_0000_0000_0000;
array[44894] <= 16'b0000_0000_0000_0000;
array[44895] <= 16'b0000_0000_0000_0000;
array[44896] <= 16'b0000_0000_0000_0000;
array[44897] <= 16'b0000_0000_0000_0000;
array[44898] <= 16'b0000_0000_0000_0000;
array[44899] <= 16'b0000_0000_0000_0000;
array[44900] <= 16'b0000_0000_0000_0000;
array[44901] <= 16'b0000_0000_0000_0000;
array[44902] <= 16'b0000_0000_0000_0000;
array[44903] <= 16'b0000_0000_0000_0000;
array[44904] <= 16'b0000_0000_0000_0000;
array[44905] <= 16'b0000_0000_0000_0000;
array[44906] <= 16'b0000_0000_0000_0000;
array[44907] <= 16'b0000_0000_0000_0000;
array[44908] <= 16'b0000_0000_0000_0000;
array[44909] <= 16'b0000_0000_0000_0000;
array[44910] <= 16'b0000_0000_0000_0000;
array[44911] <= 16'b0000_0000_0000_0000;
array[44912] <= 16'b0000_0000_0000_0000;
array[44913] <= 16'b0000_0000_0000_0000;
array[44914] <= 16'b0000_0000_0000_0000;
array[44915] <= 16'b0000_0000_0000_0000;
array[44916] <= 16'b0000_0000_0000_0000;
array[44917] <= 16'b0000_0000_0000_0000;
array[44918] <= 16'b0000_0000_0000_0000;
array[44919] <= 16'b0000_0000_0000_0000;
array[44920] <= 16'b0000_0000_0000_0000;
array[44921] <= 16'b0000_0000_0000_0000;
array[44922] <= 16'b0000_0000_0000_0000;
array[44923] <= 16'b0000_0000_0000_0000;
array[44924] <= 16'b0000_0000_0000_0000;
array[44925] <= 16'b0000_0000_0000_0000;
array[44926] <= 16'b0000_0000_0000_0000;
array[44927] <= 16'b0000_0000_0000_0000;
array[44928] <= 16'b0000_0000_0000_0000;
array[44929] <= 16'b0000_0000_0000_0000;
array[44930] <= 16'b0000_0000_0000_0000;
array[44931] <= 16'b0000_0000_0000_0000;
array[44932] <= 16'b0000_0000_0000_0000;
array[44933] <= 16'b0000_0000_0000_0000;
array[44934] <= 16'b0000_0000_0000_0000;
array[44935] <= 16'b0000_0000_0000_0000;
array[44936] <= 16'b0000_0000_0000_0000;
array[44937] <= 16'b0000_0000_0000_0000;
array[44938] <= 16'b0000_0000_0000_0000;
array[44939] <= 16'b0000_0000_0000_0000;
array[44940] <= 16'b0000_0000_0000_0000;
array[44941] <= 16'b0000_0000_0000_0000;
array[44942] <= 16'b0000_0000_0000_0000;
array[44943] <= 16'b0000_0000_0000_0000;
array[44944] <= 16'b0000_0000_0000_0000;
array[44945] <= 16'b0000_0000_0000_0000;
array[44946] <= 16'b0000_0000_0000_0000;
array[44947] <= 16'b0000_0000_0000_0000;
array[44948] <= 16'b0000_0000_0000_0000;
array[44949] <= 16'b0000_0000_0000_0000;
array[44950] <= 16'b0000_0000_0000_0000;
array[44951] <= 16'b0000_0000_0000_0000;
array[44952] <= 16'b0000_0000_0000_0000;
array[44953] <= 16'b0000_0000_0000_0000;
array[44954] <= 16'b0000_0000_0000_0000;
array[44955] <= 16'b0000_0000_0000_0000;
array[44956] <= 16'b0000_0000_0000_0000;
array[44957] <= 16'b0000_0000_0000_0000;
array[44958] <= 16'b0000_0000_0000_0000;
array[44959] <= 16'b0000_0000_0000_0000;
array[44960] <= 16'b0000_0000_0000_0000;
array[44961] <= 16'b0000_0000_0000_0000;
array[44962] <= 16'b0000_0000_0000_0000;
array[44963] <= 16'b0000_0000_0000_0000;
array[44964] <= 16'b0000_0000_0000_0000;
array[44965] <= 16'b0000_0000_0000_0000;
array[44966] <= 16'b0000_0000_0000_0000;
array[44967] <= 16'b0000_0000_0000_0000;
array[44968] <= 16'b0000_0000_0000_0000;
array[44969] <= 16'b0000_0000_0000_0000;
array[44970] <= 16'b0000_0000_0000_0000;
array[44971] <= 16'b0000_0000_0000_0000;
array[44972] <= 16'b0000_0000_0000_0000;
array[44973] <= 16'b0000_0000_0000_0000;
array[44974] <= 16'b0000_0000_0000_0000;
array[44975] <= 16'b0000_0000_0000_0000;
array[44976] <= 16'b0000_0000_0000_0000;
array[44977] <= 16'b0000_0000_0000_0000;
array[44978] <= 16'b0000_0000_0000_0000;
array[44979] <= 16'b0000_0000_0000_0000;
array[44980] <= 16'b0000_0000_0000_0000;
array[44981] <= 16'b0000_0000_0000_0000;
array[44982] <= 16'b0000_0000_0000_0000;
array[44983] <= 16'b0000_0000_0000_0000;
array[44984] <= 16'b0000_0000_0000_0000;
array[44985] <= 16'b0000_0000_0000_0000;
array[44986] <= 16'b0000_0000_0000_0000;
array[44987] <= 16'b0000_0000_0000_0000;
array[44988] <= 16'b0000_0000_0000_0000;
array[44989] <= 16'b0000_0000_0000_0000;
array[44990] <= 16'b0000_0000_0000_0000;
array[44991] <= 16'b0000_0000_0000_0000;
array[44992] <= 16'b0000_0000_0000_0000;
array[44993] <= 16'b0000_0000_0000_0000;
array[44994] <= 16'b0000_0000_0000_0000;
array[44995] <= 16'b0000_0000_0000_0000;
array[44996] <= 16'b0000_0000_0000_0000;
array[44997] <= 16'b0000_0000_0000_0000;
array[44998] <= 16'b0000_0000_0000_0000;
array[44999] <= 16'b0000_0000_0000_0000;
array[45000] <= 16'b0000_0000_0000_0000;
array[45001] <= 16'b0000_0000_0000_0000;
array[45002] <= 16'b0000_0000_0000_0000;
array[45003] <= 16'b0000_0000_0000_0000;
array[45004] <= 16'b0000_0000_0000_0000;
array[45005] <= 16'b0000_0000_0000_0000;
array[45006] <= 16'b0000_0000_0000_0000;
array[45007] <= 16'b0000_0000_0000_0000;
array[45008] <= 16'b0000_0000_0000_0000;
array[45009] <= 16'b0000_0000_0000_0000;
array[45010] <= 16'b0000_0000_0000_0000;
array[45011] <= 16'b0000_0000_0000_0000;
array[45012] <= 16'b0000_0000_0000_0000;
array[45013] <= 16'b0000_0000_0000_0000;
array[45014] <= 16'b0000_0000_0000_0000;
array[45015] <= 16'b0000_0000_0000_0000;
array[45016] <= 16'b0000_0000_0000_0000;
array[45017] <= 16'b0000_0000_0000_0000;
array[45018] <= 16'b0000_0000_0000_0000;
array[45019] <= 16'b0000_0000_0000_0000;
array[45020] <= 16'b0000_0000_0000_0000;
array[45021] <= 16'b0000_0000_0000_0000;
array[45022] <= 16'b0000_0000_0000_0000;
array[45023] <= 16'b0000_0000_0000_0000;
array[45024] <= 16'b0000_0000_0000_0000;
array[45025] <= 16'b0000_0000_0000_0000;
array[45026] <= 16'b0000_0000_0000_0000;
array[45027] <= 16'b0000_0000_0000_0000;
array[45028] <= 16'b0000_0000_0000_0000;
array[45029] <= 16'b0000_0000_0000_0000;
array[45030] <= 16'b0000_0000_0000_0000;
array[45031] <= 16'b0000_0000_0000_0000;
array[45032] <= 16'b0000_0000_0000_0000;
array[45033] <= 16'b0000_0000_0000_0000;
array[45034] <= 16'b0000_0000_0000_0000;
array[45035] <= 16'b0000_0000_0000_0000;
array[45036] <= 16'b0000_0000_0000_0000;
array[45037] <= 16'b0000_0000_0000_0000;
array[45038] <= 16'b0000_0000_0000_0000;
array[45039] <= 16'b0000_0000_0000_0000;
array[45040] <= 16'b0000_0000_0000_0000;
array[45041] <= 16'b0000_0000_0000_0000;
array[45042] <= 16'b0000_0000_0000_0000;
array[45043] <= 16'b0000_0000_0000_0000;
array[45044] <= 16'b0000_0000_0000_0000;
array[45045] <= 16'b0000_0000_0000_0000;
array[45046] <= 16'b0000_0000_0000_0000;
array[45047] <= 16'b0000_0000_0000_0000;
array[45048] <= 16'b0000_0000_0000_0000;
array[45049] <= 16'b0000_0000_0000_0000;
array[45050] <= 16'b0000_0000_0000_0000;
array[45051] <= 16'b0000_0000_0000_0000;
array[45052] <= 16'b0000_0000_0000_0000;
array[45053] <= 16'b0000_0000_0000_0000;
array[45054] <= 16'b0000_0000_0000_0000;
array[45055] <= 16'b0000_0000_0000_0000;
array[45056] <= 16'b0000_0000_0000_0000;
array[45057] <= 16'b0000_0000_0000_0000;
array[45058] <= 16'b0000_0000_0000_0000;
array[45059] <= 16'b0000_0000_0000_0000;
array[45060] <= 16'b0000_0000_0000_0000;
array[45061] <= 16'b0000_0000_0000_0000;
array[45062] <= 16'b0000_0000_0000_0000;
array[45063] <= 16'b0000_0000_0000_0000;
array[45064] <= 16'b0000_0000_0000_0000;
array[45065] <= 16'b0000_0000_0000_0000;
array[45066] <= 16'b0000_0000_0000_0000;
array[45067] <= 16'b0000_0000_0000_0000;
array[45068] <= 16'b0000_0000_0000_0000;
array[45069] <= 16'b0000_0000_0000_0000;
array[45070] <= 16'b0000_0000_0000_0000;
array[45071] <= 16'b0000_0000_0000_0000;
array[45072] <= 16'b0000_0000_0000_0000;
array[45073] <= 16'b0000_0000_0000_0000;
array[45074] <= 16'b0000_0000_0000_0000;
array[45075] <= 16'b0000_0000_0000_0000;
array[45076] <= 16'b0000_0000_0000_0000;
array[45077] <= 16'b0000_0000_0000_0000;
array[45078] <= 16'b0000_0000_0000_0000;
array[45079] <= 16'b0000_0000_0000_0000;
array[45080] <= 16'b0000_0000_0000_0000;
array[45081] <= 16'b0000_0000_0000_0000;
array[45082] <= 16'b0000_0000_0000_0000;
array[45083] <= 16'b0000_0000_0000_0000;
array[45084] <= 16'b0000_0000_0000_0000;
array[45085] <= 16'b0000_0000_0000_0000;
array[45086] <= 16'b0000_0000_0000_0000;
array[45087] <= 16'b0000_0000_0000_0000;
array[45088] <= 16'b0000_0000_0000_0000;
array[45089] <= 16'b0000_0000_0000_0000;
array[45090] <= 16'b0000_0000_0000_0000;
array[45091] <= 16'b0000_0000_0000_0000;
array[45092] <= 16'b0000_0000_0000_0000;
array[45093] <= 16'b0000_0000_0000_0000;
array[45094] <= 16'b0000_0000_0000_0000;
array[45095] <= 16'b0000_0000_0000_0000;
array[45096] <= 16'b0000_0000_0000_0000;
array[45097] <= 16'b0000_0000_0000_0000;
array[45098] <= 16'b0000_0000_0000_0000;
array[45099] <= 16'b0000_0000_0000_0000;
array[45100] <= 16'b0000_0000_0000_0000;
array[45101] <= 16'b0000_0000_0000_0000;
array[45102] <= 16'b0000_0000_0000_0000;
array[45103] <= 16'b0000_0000_0000_0000;
array[45104] <= 16'b0000_0000_0000_0000;
array[45105] <= 16'b0000_0000_0000_0000;
array[45106] <= 16'b0000_0000_0000_0000;
array[45107] <= 16'b0000_0000_0000_0000;
array[45108] <= 16'b0000_0000_0000_0000;
array[45109] <= 16'b0000_0000_0000_0000;
array[45110] <= 16'b0000_0000_0000_0000;
array[45111] <= 16'b0000_0000_0000_0000;
array[45112] <= 16'b0000_0000_0000_0000;
array[45113] <= 16'b0000_0000_0000_0000;
array[45114] <= 16'b0000_0000_0000_0000;
array[45115] <= 16'b0000_0000_0000_0000;
array[45116] <= 16'b0000_0000_0000_0000;
array[45117] <= 16'b0000_0000_0000_0000;
array[45118] <= 16'b0000_0000_0000_0000;
array[45119] <= 16'b0000_0000_0000_0000;
array[45120] <= 16'b0000_0000_0000_0000;
array[45121] <= 16'b0000_0000_0000_0000;
array[45122] <= 16'b0000_0000_0000_0000;
array[45123] <= 16'b0000_0000_0000_0000;
array[45124] <= 16'b0000_0000_0000_0000;
array[45125] <= 16'b0000_0000_0000_0000;
array[45126] <= 16'b0000_0000_0000_0000;
array[45127] <= 16'b0000_0000_0000_0000;
array[45128] <= 16'b0000_0000_0000_0000;
array[45129] <= 16'b0000_0000_0000_0000;
array[45130] <= 16'b0000_0000_0000_0000;
array[45131] <= 16'b0000_0000_0000_0000;
array[45132] <= 16'b0000_0000_0000_0000;
array[45133] <= 16'b0000_0000_0000_0000;
array[45134] <= 16'b0000_0000_0000_0000;
array[45135] <= 16'b0000_0000_0000_0000;
array[45136] <= 16'b0000_0000_0000_0000;
array[45137] <= 16'b0000_0000_0000_0000;
array[45138] <= 16'b0000_0000_0000_0000;
array[45139] <= 16'b0000_0000_0000_0000;
array[45140] <= 16'b0000_0000_0000_0000;
array[45141] <= 16'b0000_0000_0000_0000;
array[45142] <= 16'b0000_0000_0000_0000;
array[45143] <= 16'b0000_0000_0000_0000;
array[45144] <= 16'b0000_0000_0000_0000;
array[45145] <= 16'b0000_0000_0000_0000;
array[45146] <= 16'b0000_0000_0000_0000;
array[45147] <= 16'b0000_0000_0000_0000;
array[45148] <= 16'b0000_0000_0000_0000;
array[45149] <= 16'b0000_0000_0000_0000;
array[45150] <= 16'b0000_0000_0000_0000;
array[45151] <= 16'b0000_0000_0000_0000;
array[45152] <= 16'b0000_0000_0000_0000;
array[45153] <= 16'b0000_0000_0000_0000;
array[45154] <= 16'b0000_0000_0000_0000;
array[45155] <= 16'b0000_0000_0000_0000;
array[45156] <= 16'b0000_0000_0000_0000;
array[45157] <= 16'b0000_0000_0000_0000;
array[45158] <= 16'b0000_0000_0000_0000;
array[45159] <= 16'b0000_0000_0000_0000;
array[45160] <= 16'b0000_0000_0000_0000;
array[45161] <= 16'b0000_0000_0000_0000;
array[45162] <= 16'b0000_0000_0000_0000;
array[45163] <= 16'b0000_0000_0000_0000;
array[45164] <= 16'b0000_0000_0000_0000;
array[45165] <= 16'b0000_0000_0000_0000;
array[45166] <= 16'b0000_0000_0000_0000;
array[45167] <= 16'b0000_0000_0000_0000;
array[45168] <= 16'b0000_0000_0000_0000;
array[45169] <= 16'b0000_0000_0000_0000;
array[45170] <= 16'b0000_0000_0000_0000;
array[45171] <= 16'b0000_0000_0000_0000;
array[45172] <= 16'b0000_0000_0000_0000;
array[45173] <= 16'b0000_0000_0000_0000;
array[45174] <= 16'b0000_0000_0000_0000;
array[45175] <= 16'b0000_0000_0000_0000;
array[45176] <= 16'b0000_0000_0000_0000;
array[45177] <= 16'b0000_0000_0000_0000;
array[45178] <= 16'b0000_0000_0000_0000;
array[45179] <= 16'b0000_0000_0000_0000;
array[45180] <= 16'b0000_0000_0000_0000;
array[45181] <= 16'b0000_0000_0000_0000;
array[45182] <= 16'b0000_0000_0000_0000;
array[45183] <= 16'b0000_0000_0000_0000;
array[45184] <= 16'b0000_0000_0000_0000;
array[45185] <= 16'b0000_0000_0000_0000;
array[45186] <= 16'b0000_0000_0000_0000;
array[45187] <= 16'b0000_0000_0000_0000;
array[45188] <= 16'b0000_0000_0000_0000;
array[45189] <= 16'b0000_0000_0000_0000;
array[45190] <= 16'b0000_0000_0000_0000;
array[45191] <= 16'b0000_0000_0000_0000;
array[45192] <= 16'b0000_0000_0000_0000;
array[45193] <= 16'b0000_0000_0000_0000;
array[45194] <= 16'b0000_0000_0000_0000;
array[45195] <= 16'b0000_0000_0000_0000;
array[45196] <= 16'b0000_0000_0000_0000;
array[45197] <= 16'b0000_0000_0000_0000;
array[45198] <= 16'b0000_0000_0000_0000;
array[45199] <= 16'b0000_0000_0000_0000;
array[45200] <= 16'b0000_0000_0000_0000;
array[45201] <= 16'b0000_0000_0000_0000;
array[45202] <= 16'b0000_0000_0000_0000;
array[45203] <= 16'b0000_0000_0000_0000;
array[45204] <= 16'b0000_0000_0000_0000;
array[45205] <= 16'b0000_0000_0000_0000;
array[45206] <= 16'b0000_0000_0000_0000;
array[45207] <= 16'b0000_0000_0000_0000;
array[45208] <= 16'b0000_0000_0000_0000;
array[45209] <= 16'b0000_0000_0000_0000;
array[45210] <= 16'b0000_0000_0000_0000;
array[45211] <= 16'b0000_0000_0000_0000;
array[45212] <= 16'b0000_0000_0000_0000;
array[45213] <= 16'b0000_0000_0000_0000;
array[45214] <= 16'b0000_0000_0000_0000;
array[45215] <= 16'b0000_0000_0000_0000;
array[45216] <= 16'b0000_0000_0000_0000;
array[45217] <= 16'b0000_0000_0000_0000;
array[45218] <= 16'b0000_0000_0000_0000;
array[45219] <= 16'b0000_0000_0000_0000;
array[45220] <= 16'b0000_0000_0000_0000;
array[45221] <= 16'b0000_0000_0000_0000;
array[45222] <= 16'b0000_0000_0000_0000;
array[45223] <= 16'b0000_0000_0000_0000;
array[45224] <= 16'b0000_0000_0000_0000;
array[45225] <= 16'b0000_0000_0000_0000;
array[45226] <= 16'b0000_0000_0000_0000;
array[45227] <= 16'b0000_0000_0000_0000;
array[45228] <= 16'b0000_0000_0000_0000;
array[45229] <= 16'b0000_0000_0000_0000;
array[45230] <= 16'b0000_0000_0000_0000;
array[45231] <= 16'b0000_0000_0000_0000;
array[45232] <= 16'b0000_0000_0000_0000;
array[45233] <= 16'b0000_0000_0000_0000;
array[45234] <= 16'b0000_0000_0000_0000;
array[45235] <= 16'b0000_0000_0000_0000;
array[45236] <= 16'b0000_0000_0000_0000;
array[45237] <= 16'b0000_0000_0000_0000;
array[45238] <= 16'b0000_0000_0000_0000;
array[45239] <= 16'b0000_0000_0000_0000;
array[45240] <= 16'b0000_0000_0000_0000;
array[45241] <= 16'b0000_0000_0000_0000;
array[45242] <= 16'b0000_0000_0000_0000;
array[45243] <= 16'b0000_0000_0000_0000;
array[45244] <= 16'b0000_0000_0000_0000;
array[45245] <= 16'b0000_0000_0000_0000;
array[45246] <= 16'b0000_0000_0000_0000;
array[45247] <= 16'b0000_0000_0000_0000;
array[45248] <= 16'b0000_0000_0000_0000;
array[45249] <= 16'b0000_0000_0000_0000;
array[45250] <= 16'b0000_0000_0000_0000;
array[45251] <= 16'b0000_0000_0000_0000;
array[45252] <= 16'b0000_0000_0000_0000;
array[45253] <= 16'b0000_0000_0000_0000;
array[45254] <= 16'b0000_0000_0000_0000;
array[45255] <= 16'b0000_0000_0000_0000;
array[45256] <= 16'b0000_0000_0000_0000;
array[45257] <= 16'b0000_0000_0000_0000;
array[45258] <= 16'b0000_0000_0000_0000;
array[45259] <= 16'b0000_0000_0000_0000;
array[45260] <= 16'b0000_0000_0000_0000;
array[45261] <= 16'b0000_0000_0000_0000;
array[45262] <= 16'b0000_0000_0000_0000;
array[45263] <= 16'b0000_0000_0000_0000;
array[45264] <= 16'b0000_0000_0000_0000;
array[45265] <= 16'b0000_0000_0000_0000;
array[45266] <= 16'b0000_0000_0000_0000;
array[45267] <= 16'b0000_0000_0000_0000;
array[45268] <= 16'b0000_0000_0000_0000;
array[45269] <= 16'b0000_0000_0000_0000;
array[45270] <= 16'b0000_0000_0000_0000;
array[45271] <= 16'b0000_0000_0000_0000;
array[45272] <= 16'b0000_0000_0000_0000;
array[45273] <= 16'b0000_0000_0000_0000;
array[45274] <= 16'b0000_0000_0000_0000;
array[45275] <= 16'b0000_0000_0000_0000;
array[45276] <= 16'b0000_0000_0000_0000;
array[45277] <= 16'b0000_0000_0000_0000;
array[45278] <= 16'b0000_0000_0000_0000;
array[45279] <= 16'b0000_0000_0000_0000;
array[45280] <= 16'b0000_0000_0000_0000;
array[45281] <= 16'b0000_0000_0000_0000;
array[45282] <= 16'b0000_0000_0000_0000;
array[45283] <= 16'b0000_0000_0000_0000;
array[45284] <= 16'b0000_0000_0000_0000;
array[45285] <= 16'b0000_0000_0000_0000;
array[45286] <= 16'b0000_0000_0000_0000;
array[45287] <= 16'b0000_0000_0000_0000;
array[45288] <= 16'b0000_0000_0000_0000;
array[45289] <= 16'b0000_0000_0000_0000;
array[45290] <= 16'b0000_0000_0000_0000;
array[45291] <= 16'b0000_0000_0000_0000;
array[45292] <= 16'b0000_0000_0000_0000;
array[45293] <= 16'b0000_0000_0000_0000;
array[45294] <= 16'b0000_0000_0000_0000;
array[45295] <= 16'b0000_0000_0000_0000;
array[45296] <= 16'b0000_0000_0000_0000;
array[45297] <= 16'b0000_0000_0000_0000;
array[45298] <= 16'b0000_0000_0000_0000;
array[45299] <= 16'b0000_0000_0000_0000;
array[45300] <= 16'b0000_0000_0000_0000;
array[45301] <= 16'b0000_0000_0000_0000;
array[45302] <= 16'b0000_0000_0000_0000;
array[45303] <= 16'b0000_0000_0000_0000;
array[45304] <= 16'b0000_0000_0000_0000;
array[45305] <= 16'b0000_0000_0000_0000;
array[45306] <= 16'b0000_0000_0000_0000;
array[45307] <= 16'b0000_0000_0000_0000;
array[45308] <= 16'b0000_0000_0000_0000;
array[45309] <= 16'b0000_0000_0000_0000;
array[45310] <= 16'b0000_0000_0000_0000;
array[45311] <= 16'b0000_0000_0000_0000;
array[45312] <= 16'b0000_0000_0000_0000;
array[45313] <= 16'b0000_0000_0000_0000;
array[45314] <= 16'b0000_0000_0000_0000;
array[45315] <= 16'b0000_0000_0000_0000;
array[45316] <= 16'b0000_0000_0000_0000;
array[45317] <= 16'b0000_0000_0000_0000;
array[45318] <= 16'b0000_0000_0000_0000;
array[45319] <= 16'b0000_0000_0000_0000;
array[45320] <= 16'b0000_0000_0000_0000;
array[45321] <= 16'b0000_0000_0000_0000;
array[45322] <= 16'b0000_0000_0000_0000;
array[45323] <= 16'b0000_0000_0000_0000;
array[45324] <= 16'b0000_0000_0000_0000;
array[45325] <= 16'b0000_0000_0000_0000;
array[45326] <= 16'b0000_0000_0000_0000;
array[45327] <= 16'b0000_0000_0000_0000;
array[45328] <= 16'b0000_0000_0000_0000;
array[45329] <= 16'b0000_0000_0000_0000;
array[45330] <= 16'b0000_0000_0000_0000;
array[45331] <= 16'b0000_0000_0000_0000;
array[45332] <= 16'b0000_0000_0000_0000;
array[45333] <= 16'b0000_0000_0000_0000;
array[45334] <= 16'b0000_0000_0000_0000;
array[45335] <= 16'b0000_0000_0000_0000;
array[45336] <= 16'b0000_0000_0000_0000;
array[45337] <= 16'b0000_0000_0000_0000;
array[45338] <= 16'b0000_0000_0000_0000;
array[45339] <= 16'b0000_0000_0000_0000;
array[45340] <= 16'b0000_0000_0000_0000;
array[45341] <= 16'b0000_0000_0000_0000;
array[45342] <= 16'b0000_0000_0000_0000;
array[45343] <= 16'b0000_0000_0000_0000;
array[45344] <= 16'b0000_0000_0000_0000;
array[45345] <= 16'b0000_0000_0000_0000;
array[45346] <= 16'b0000_0000_0000_0000;
array[45347] <= 16'b0000_0000_0000_0000;
array[45348] <= 16'b0000_0000_0000_0000;
array[45349] <= 16'b0000_0000_0000_0000;
array[45350] <= 16'b0000_0000_0000_0000;
array[45351] <= 16'b0000_0000_0000_0000;
array[45352] <= 16'b0000_0000_0000_0000;
array[45353] <= 16'b0000_0000_0000_0000;
array[45354] <= 16'b0000_0000_0000_0000;
array[45355] <= 16'b0000_0000_0000_0000;
array[45356] <= 16'b0000_0000_0000_0000;
array[45357] <= 16'b0000_0000_0000_0000;
array[45358] <= 16'b0000_0000_0000_0000;
array[45359] <= 16'b0000_0000_0000_0000;
array[45360] <= 16'b0000_0000_0000_0000;
array[45361] <= 16'b0000_0000_0000_0000;
array[45362] <= 16'b0000_0000_0000_0000;
array[45363] <= 16'b0000_0000_0000_0000;
array[45364] <= 16'b0000_0000_0000_0000;
array[45365] <= 16'b0000_0000_0000_0000;
array[45366] <= 16'b0000_0000_0000_0000;
array[45367] <= 16'b0000_0000_0000_0000;
array[45368] <= 16'b0000_0000_0000_0000;
array[45369] <= 16'b0000_0000_0000_0000;
array[45370] <= 16'b0000_0000_0000_0000;
array[45371] <= 16'b0000_0000_0000_0000;
array[45372] <= 16'b0000_0000_0000_0000;
array[45373] <= 16'b0000_0000_0000_0000;
array[45374] <= 16'b0000_0000_0000_0000;
array[45375] <= 16'b0000_0000_0000_0000;
array[45376] <= 16'b0000_0000_0000_0000;
array[45377] <= 16'b0000_0000_0000_0000;
array[45378] <= 16'b0000_0000_0000_0000;
array[45379] <= 16'b0000_0000_0000_0000;
array[45380] <= 16'b0000_0000_0000_0000;
array[45381] <= 16'b0000_0000_0000_0000;
array[45382] <= 16'b0000_0000_0000_0000;
array[45383] <= 16'b0000_0000_0000_0000;
array[45384] <= 16'b0000_0000_0000_0000;
array[45385] <= 16'b0000_0000_0000_0000;
array[45386] <= 16'b0000_0000_0000_0000;
array[45387] <= 16'b0000_0000_0000_0000;
array[45388] <= 16'b0000_0000_0000_0000;
array[45389] <= 16'b0000_0000_0000_0000;
array[45390] <= 16'b0000_0000_0000_0000;
array[45391] <= 16'b0000_0000_0000_0000;
array[45392] <= 16'b0000_0000_0000_0000;
array[45393] <= 16'b0000_0000_0000_0000;
array[45394] <= 16'b0000_0000_0000_0000;
array[45395] <= 16'b0000_0000_0000_0000;
array[45396] <= 16'b0000_0000_0000_0000;
array[45397] <= 16'b0000_0000_0000_0000;
array[45398] <= 16'b0000_0000_0000_0000;
array[45399] <= 16'b0000_0000_0000_0000;
array[45400] <= 16'b0000_0000_0000_0000;
array[45401] <= 16'b0000_0000_0000_0000;
array[45402] <= 16'b0000_0000_0000_0000;
array[45403] <= 16'b0000_0000_0000_0000;
array[45404] <= 16'b0000_0000_0000_0000;
array[45405] <= 16'b0000_0000_0000_0000;
array[45406] <= 16'b0000_0000_0000_0000;
array[45407] <= 16'b0000_0000_0000_0000;
array[45408] <= 16'b0000_0000_0000_0000;
array[45409] <= 16'b0000_0000_0000_0000;
array[45410] <= 16'b0000_0000_0000_0000;
array[45411] <= 16'b0000_0000_0000_0000;
array[45412] <= 16'b0000_0000_0000_0000;
array[45413] <= 16'b0000_0000_0000_0000;
array[45414] <= 16'b0000_0000_0000_0000;
array[45415] <= 16'b0000_0000_0000_0000;
array[45416] <= 16'b0000_0000_0000_0000;
array[45417] <= 16'b0000_0000_0000_0000;
array[45418] <= 16'b0000_0000_0000_0000;
array[45419] <= 16'b0000_0000_0000_0000;
array[45420] <= 16'b0000_0000_0000_0000;
array[45421] <= 16'b0000_0000_0000_0000;
array[45422] <= 16'b0000_0000_0000_0000;
array[45423] <= 16'b0000_0000_0000_0000;
array[45424] <= 16'b0000_0000_0000_0000;
array[45425] <= 16'b0000_0000_0000_0000;
array[45426] <= 16'b0000_0000_0000_0000;
array[45427] <= 16'b0000_0000_0000_0000;
array[45428] <= 16'b0000_0000_0000_0000;
array[45429] <= 16'b0000_0000_0000_0000;
array[45430] <= 16'b0000_0000_0000_0000;
array[45431] <= 16'b0000_0000_0000_0000;
array[45432] <= 16'b0000_0000_0000_0000;
array[45433] <= 16'b0000_0000_0000_0000;
array[45434] <= 16'b0000_0000_0000_0000;
array[45435] <= 16'b0000_0000_0000_0000;
array[45436] <= 16'b0000_0000_0000_0000;
array[45437] <= 16'b0000_0000_0000_0000;
array[45438] <= 16'b0000_0000_0000_0000;
array[45439] <= 16'b0000_0000_0000_0000;
array[45440] <= 16'b0000_0000_0000_0000;
array[45441] <= 16'b0000_0000_0000_0000;
array[45442] <= 16'b0000_0000_0000_0000;
array[45443] <= 16'b0000_0000_0000_0000;
array[45444] <= 16'b0000_0000_0000_0000;
array[45445] <= 16'b0000_0000_0000_0000;
array[45446] <= 16'b0000_0000_0000_0000;
array[45447] <= 16'b0000_0000_0000_0000;
array[45448] <= 16'b0000_0000_0000_0000;
array[45449] <= 16'b0000_0000_0000_0000;
array[45450] <= 16'b0000_0000_0000_0000;
array[45451] <= 16'b0000_0000_0000_0000;
array[45452] <= 16'b0000_0000_0000_0000;
array[45453] <= 16'b0000_0000_0000_0000;
array[45454] <= 16'b0000_0000_0000_0000;
array[45455] <= 16'b0000_0000_0000_0000;
array[45456] <= 16'b0000_0000_0000_0000;
array[45457] <= 16'b0000_0000_0000_0000;
array[45458] <= 16'b0000_0000_0000_0000;
array[45459] <= 16'b0000_0000_0000_0000;
array[45460] <= 16'b0000_0000_0000_0000;
array[45461] <= 16'b0000_0000_0000_0000;
array[45462] <= 16'b0000_0000_0000_0000;
array[45463] <= 16'b0000_0000_0000_0000;
array[45464] <= 16'b0000_0000_0000_0000;
array[45465] <= 16'b0000_0000_0000_0000;
array[45466] <= 16'b0000_0000_0000_0000;
array[45467] <= 16'b0000_0000_0000_0000;
array[45468] <= 16'b0000_0000_0000_0000;
array[45469] <= 16'b0000_0000_0000_0000;
array[45470] <= 16'b0000_0000_0000_0000;
array[45471] <= 16'b0000_0000_0000_0000;
array[45472] <= 16'b0000_0000_0000_0000;
array[45473] <= 16'b0000_0000_0000_0000;
array[45474] <= 16'b0000_0000_0000_0000;
array[45475] <= 16'b0000_0000_0000_0000;
array[45476] <= 16'b0000_0000_0000_0000;
array[45477] <= 16'b0000_0000_0000_0000;
array[45478] <= 16'b0000_0000_0000_0000;
array[45479] <= 16'b0000_0000_0000_0000;
array[45480] <= 16'b0000_0000_0000_0000;
array[45481] <= 16'b0000_0000_0000_0000;
array[45482] <= 16'b0000_0000_0000_0000;
array[45483] <= 16'b0000_0000_0000_0000;
array[45484] <= 16'b0000_0000_0000_0000;
array[45485] <= 16'b0000_0000_0000_0000;
array[45486] <= 16'b0000_0000_0000_0000;
array[45487] <= 16'b0000_0000_0000_0000;
array[45488] <= 16'b0000_0000_0000_0000;
array[45489] <= 16'b0000_0000_0000_0000;
array[45490] <= 16'b0000_0000_0000_0000;
array[45491] <= 16'b0000_0000_0000_0000;
array[45492] <= 16'b0000_0000_0000_0000;
array[45493] <= 16'b0000_0000_0000_0000;
array[45494] <= 16'b0000_0000_0000_0000;
array[45495] <= 16'b0000_0000_0000_0000;
array[45496] <= 16'b0000_0000_0000_0000;
array[45497] <= 16'b0000_0000_0000_0000;
array[45498] <= 16'b0000_0000_0000_0000;
array[45499] <= 16'b0000_0000_0000_0000;
array[45500] <= 16'b0000_0000_0000_0000;
array[45501] <= 16'b0000_0000_0000_0000;
array[45502] <= 16'b0000_0000_0000_0000;
array[45503] <= 16'b0000_0000_0000_0000;
array[45504] <= 16'b0000_0000_0000_0000;
array[45505] <= 16'b0000_0000_0000_0000;
array[45506] <= 16'b0000_0000_0000_0000;
array[45507] <= 16'b0000_0000_0000_0000;
array[45508] <= 16'b0000_0000_0000_0000;
array[45509] <= 16'b0000_0000_0000_0000;
array[45510] <= 16'b0000_0000_0000_0000;
array[45511] <= 16'b0000_0000_0000_0000;
array[45512] <= 16'b0000_0000_0000_0000;
array[45513] <= 16'b0000_0000_0000_0000;
array[45514] <= 16'b0000_0000_0000_0000;
array[45515] <= 16'b0000_0000_0000_0000;
array[45516] <= 16'b0000_0000_0000_0000;
array[45517] <= 16'b0000_0000_0000_0000;
array[45518] <= 16'b0000_0000_0000_0000;
array[45519] <= 16'b0000_0000_0000_0000;
array[45520] <= 16'b0000_0000_0000_0000;
array[45521] <= 16'b0000_0000_0000_0000;
array[45522] <= 16'b0000_0000_0000_0000;
array[45523] <= 16'b0000_0000_0000_0000;
array[45524] <= 16'b0000_0000_0000_0000;
array[45525] <= 16'b0000_0000_0000_0000;
array[45526] <= 16'b0000_0000_0000_0000;
array[45527] <= 16'b0000_0000_0000_0000;
array[45528] <= 16'b0000_0000_0000_0000;
array[45529] <= 16'b0000_0000_0000_0000;
array[45530] <= 16'b0000_0000_0000_0000;
array[45531] <= 16'b0000_0000_0000_0000;
array[45532] <= 16'b0000_0000_0000_0000;
array[45533] <= 16'b0000_0000_0000_0000;
array[45534] <= 16'b0000_0000_0000_0000;
array[45535] <= 16'b0000_0000_0000_0000;
array[45536] <= 16'b0000_0000_0000_0000;
array[45537] <= 16'b0000_0000_0000_0000;
array[45538] <= 16'b0000_0000_0000_0000;
array[45539] <= 16'b0000_0000_0000_0000;
array[45540] <= 16'b0000_0000_0000_0000;
array[45541] <= 16'b0000_0000_0000_0000;
array[45542] <= 16'b0000_0000_0000_0000;
array[45543] <= 16'b0000_0000_0000_0000;
array[45544] <= 16'b0000_0000_0000_0000;
array[45545] <= 16'b0000_0000_0000_0000;
array[45546] <= 16'b0000_0000_0000_0000;
array[45547] <= 16'b0000_0000_0000_0000;
array[45548] <= 16'b0000_0000_0000_0000;
array[45549] <= 16'b0000_0000_0000_0000;
array[45550] <= 16'b0000_0000_0000_0000;
array[45551] <= 16'b0000_0000_0000_0000;
array[45552] <= 16'b0000_0000_0000_0000;
array[45553] <= 16'b0000_0000_0000_0000;
array[45554] <= 16'b0000_0000_0000_0000;
array[45555] <= 16'b0000_0000_0000_0000;
array[45556] <= 16'b0000_0000_0000_0000;
array[45557] <= 16'b0000_0000_0000_0000;
array[45558] <= 16'b0000_0000_0000_0000;
array[45559] <= 16'b0000_0000_0000_0000;
array[45560] <= 16'b0000_0000_0000_0000;
array[45561] <= 16'b0000_0000_0000_0000;
array[45562] <= 16'b0000_0000_0000_0000;
array[45563] <= 16'b0000_0000_0000_0000;
array[45564] <= 16'b0000_0000_0000_0000;
array[45565] <= 16'b0000_0000_0000_0000;
array[45566] <= 16'b0000_0000_0000_0000;
array[45567] <= 16'b0000_0000_0000_0000;
array[45568] <= 16'b0000_0000_0000_0000;
array[45569] <= 16'b0000_0000_0000_0000;
array[45570] <= 16'b0000_0000_0000_0000;
array[45571] <= 16'b0000_0000_0000_0000;
array[45572] <= 16'b0000_0000_0000_0000;
array[45573] <= 16'b0000_0000_0000_0000;
array[45574] <= 16'b0000_0000_0000_0000;
array[45575] <= 16'b0000_0000_0000_0000;
array[45576] <= 16'b0000_0000_0000_0000;
array[45577] <= 16'b0000_0000_0000_0000;
array[45578] <= 16'b0000_0000_0000_0000;
array[45579] <= 16'b0000_0000_0000_0000;
array[45580] <= 16'b0000_0000_0000_0000;
array[45581] <= 16'b0000_0000_0000_0000;
array[45582] <= 16'b0000_0000_0000_0000;
array[45583] <= 16'b0000_0000_0000_0000;
array[45584] <= 16'b0000_0000_0000_0000;
array[45585] <= 16'b0000_0000_0000_0000;
array[45586] <= 16'b0000_0000_0000_0000;
array[45587] <= 16'b0000_0000_0000_0000;
array[45588] <= 16'b0000_0000_0000_0000;
array[45589] <= 16'b0000_0000_0000_0000;
array[45590] <= 16'b0000_0000_0000_0000;
array[45591] <= 16'b0000_0000_0000_0000;
array[45592] <= 16'b0000_0000_0000_0000;
array[45593] <= 16'b0000_0000_0000_0000;
array[45594] <= 16'b0000_0000_0000_0000;
array[45595] <= 16'b0000_0000_0000_0000;
array[45596] <= 16'b0000_0000_0000_0000;
array[45597] <= 16'b0000_0000_0000_0000;
array[45598] <= 16'b0000_0000_0000_0000;
array[45599] <= 16'b0000_0000_0000_0000;
array[45600] <= 16'b0000_0000_0000_0000;
array[45601] <= 16'b0000_0000_0000_0000;
array[45602] <= 16'b0000_0000_0000_0000;
array[45603] <= 16'b0000_0000_0000_0000;
array[45604] <= 16'b0000_0000_0000_0000;
array[45605] <= 16'b0000_0000_0000_0000;
array[45606] <= 16'b0000_0000_0000_0000;
array[45607] <= 16'b0000_0000_0000_0000;
array[45608] <= 16'b0000_0000_0000_0000;
array[45609] <= 16'b0000_0000_0000_0000;
array[45610] <= 16'b0000_0000_0000_0000;
array[45611] <= 16'b0000_0000_0000_0000;
array[45612] <= 16'b0000_0000_0000_0000;
array[45613] <= 16'b0000_0000_0000_0000;
array[45614] <= 16'b0000_0000_0000_0000;
array[45615] <= 16'b0000_0000_0000_0000;
array[45616] <= 16'b0000_0000_0000_0000;
array[45617] <= 16'b0000_0000_0000_0000;
array[45618] <= 16'b0000_0000_0000_0000;
array[45619] <= 16'b0000_0000_0000_0000;
array[45620] <= 16'b0000_0000_0000_0000;
array[45621] <= 16'b0000_0000_0000_0000;
array[45622] <= 16'b0000_0000_0000_0000;
array[45623] <= 16'b0000_0000_0000_0000;
array[45624] <= 16'b0000_0000_0000_0000;
array[45625] <= 16'b0000_0000_0000_0000;
array[45626] <= 16'b0000_0000_0000_0000;
array[45627] <= 16'b0000_0000_0000_0000;
array[45628] <= 16'b0000_0000_0000_0000;
array[45629] <= 16'b0000_0000_0000_0000;
array[45630] <= 16'b0000_0000_0000_0000;
array[45631] <= 16'b0000_0000_0000_0000;
array[45632] <= 16'b0000_0000_0000_0000;
array[45633] <= 16'b0000_0000_0000_0000;
array[45634] <= 16'b0000_0000_0000_0000;
array[45635] <= 16'b0000_0000_0000_0000;
array[45636] <= 16'b0000_0000_0000_0000;
array[45637] <= 16'b0000_0000_0000_0000;
array[45638] <= 16'b0000_0000_0000_0000;
array[45639] <= 16'b0000_0000_0000_0000;
array[45640] <= 16'b0000_0000_0000_0000;
array[45641] <= 16'b0000_0000_0000_0000;
array[45642] <= 16'b0000_0000_0000_0000;
array[45643] <= 16'b0000_0000_0000_0000;
array[45644] <= 16'b0000_0000_0000_0000;
array[45645] <= 16'b0000_0000_0000_0000;
array[45646] <= 16'b0000_0000_0000_0000;
array[45647] <= 16'b0000_0000_0000_0000;
array[45648] <= 16'b0000_0000_0000_0000;
array[45649] <= 16'b0000_0000_0000_0000;
array[45650] <= 16'b0000_0000_0000_0000;
array[45651] <= 16'b0000_0000_0000_0000;
array[45652] <= 16'b0000_0000_0000_0000;
array[45653] <= 16'b0000_0000_0000_0000;
array[45654] <= 16'b0000_0000_0000_0000;
array[45655] <= 16'b0000_0000_0000_0000;
array[45656] <= 16'b0000_0000_0000_0000;
array[45657] <= 16'b0000_0000_0000_0000;
array[45658] <= 16'b0000_0000_0000_0000;
array[45659] <= 16'b0000_0000_0000_0000;
array[45660] <= 16'b0000_0000_0000_0000;
array[45661] <= 16'b0000_0000_0000_0000;
array[45662] <= 16'b0000_0000_0000_0000;
array[45663] <= 16'b0000_0000_0000_0000;
array[45664] <= 16'b0000_0000_0000_0000;
array[45665] <= 16'b0000_0000_0000_0000;
array[45666] <= 16'b0000_0000_0000_0000;
array[45667] <= 16'b0000_0000_0000_0000;
array[45668] <= 16'b0000_0000_0000_0000;
array[45669] <= 16'b0000_0000_0000_0000;
array[45670] <= 16'b0000_0000_0000_0000;
array[45671] <= 16'b0000_0000_0000_0000;
array[45672] <= 16'b0000_0000_0000_0000;
array[45673] <= 16'b0000_0000_0000_0000;
array[45674] <= 16'b0000_0000_0000_0000;
array[45675] <= 16'b0000_0000_0000_0000;
array[45676] <= 16'b0000_0000_0000_0000;
array[45677] <= 16'b0000_0000_0000_0000;
array[45678] <= 16'b0000_0000_0000_0000;
array[45679] <= 16'b0000_0000_0000_0000;
array[45680] <= 16'b0000_0000_0000_0000;
array[45681] <= 16'b0000_0000_0000_0000;
array[45682] <= 16'b0000_0000_0000_0000;
array[45683] <= 16'b0000_0000_0000_0000;
array[45684] <= 16'b0000_0000_0000_0000;
array[45685] <= 16'b0000_0000_0000_0000;
array[45686] <= 16'b0000_0000_0000_0000;
array[45687] <= 16'b0000_0000_0000_0000;
array[45688] <= 16'b0000_0000_0000_0000;
array[45689] <= 16'b0000_0000_0000_0000;
array[45690] <= 16'b0000_0000_0000_0000;
array[45691] <= 16'b0000_0000_0000_0000;
array[45692] <= 16'b0000_0000_0000_0000;
array[45693] <= 16'b0000_0000_0000_0000;
array[45694] <= 16'b0000_0000_0000_0000;
array[45695] <= 16'b0000_0000_0000_0000;
array[45696] <= 16'b0000_0000_0000_0000;
array[45697] <= 16'b0000_0000_0000_0000;
array[45698] <= 16'b0000_0000_0000_0000;
array[45699] <= 16'b0000_0000_0000_0000;
array[45700] <= 16'b0000_0000_0000_0000;
array[45701] <= 16'b0000_0000_0000_0000;
array[45702] <= 16'b0000_0000_0000_0000;
array[45703] <= 16'b0000_0000_0000_0000;
array[45704] <= 16'b0000_0000_0000_0000;
array[45705] <= 16'b0000_0000_0000_0000;
array[45706] <= 16'b0000_0000_0000_0000;
array[45707] <= 16'b0000_0000_0000_0000;
array[45708] <= 16'b0000_0000_0000_0000;
array[45709] <= 16'b0000_0000_0000_0000;
array[45710] <= 16'b0000_0000_0000_0000;
array[45711] <= 16'b0000_0000_0000_0000;
array[45712] <= 16'b0000_0000_0000_0000;
array[45713] <= 16'b0000_0000_0000_0000;
array[45714] <= 16'b0000_0000_0000_0000;
array[45715] <= 16'b0000_0000_0000_0000;
array[45716] <= 16'b0000_0000_0000_0000;
array[45717] <= 16'b0000_0000_0000_0000;
array[45718] <= 16'b0000_0000_0000_0000;
array[45719] <= 16'b0000_0000_0000_0000;
array[45720] <= 16'b0000_0000_0000_0000;
array[45721] <= 16'b0000_0000_0000_0000;
array[45722] <= 16'b0000_0000_0000_0000;
array[45723] <= 16'b0000_0000_0000_0000;
array[45724] <= 16'b0000_0000_0000_0000;
array[45725] <= 16'b0000_0000_0000_0000;
array[45726] <= 16'b0000_0000_0000_0000;
array[45727] <= 16'b0000_0000_0000_0000;
array[45728] <= 16'b0000_0000_0000_0000;
array[45729] <= 16'b0000_0000_0000_0000;
array[45730] <= 16'b0000_0000_0000_0000;
array[45731] <= 16'b0000_0000_0000_0000;
array[45732] <= 16'b0000_0000_0000_0000;
array[45733] <= 16'b0000_0000_0000_0000;
array[45734] <= 16'b0000_0000_0000_0000;
array[45735] <= 16'b0000_0000_0000_0000;
array[45736] <= 16'b0000_0000_0000_0000;
array[45737] <= 16'b0000_0000_0000_0000;
array[45738] <= 16'b0000_0000_0000_0000;
array[45739] <= 16'b0000_0000_0000_0000;
array[45740] <= 16'b0000_0000_0000_0000;
array[45741] <= 16'b0000_0000_0000_0000;
array[45742] <= 16'b0000_0000_0000_0000;
array[45743] <= 16'b0000_0000_0000_0000;
array[45744] <= 16'b0000_0000_0000_0000;
array[45745] <= 16'b0000_0000_0000_0000;
array[45746] <= 16'b0000_0000_0000_0000;
array[45747] <= 16'b0000_0000_0000_0000;
array[45748] <= 16'b0000_0000_0000_0000;
array[45749] <= 16'b0000_0000_0000_0000;
array[45750] <= 16'b0000_0000_0000_0000;
array[45751] <= 16'b0000_0000_0000_0000;
array[45752] <= 16'b0000_0000_0000_0000;
array[45753] <= 16'b0000_0000_0000_0000;
array[45754] <= 16'b0000_0000_0000_0000;
array[45755] <= 16'b0000_0000_0000_0000;
array[45756] <= 16'b0000_0000_0000_0000;
array[45757] <= 16'b0000_0000_0000_0000;
array[45758] <= 16'b0000_0000_0000_0000;
array[45759] <= 16'b0000_0000_0000_0000;
array[45760] <= 16'b0000_0000_0000_0000;
array[45761] <= 16'b0000_0000_0000_0000;
array[45762] <= 16'b0000_0000_0000_0000;
array[45763] <= 16'b0000_0000_0000_0000;
array[45764] <= 16'b0000_0000_0000_0000;
array[45765] <= 16'b0000_0000_0000_0000;
array[45766] <= 16'b0000_0000_0000_0000;
array[45767] <= 16'b0000_0000_0000_0000;
array[45768] <= 16'b0000_0000_0000_0000;
array[45769] <= 16'b0000_0000_0000_0000;
array[45770] <= 16'b0000_0000_0000_0000;
array[45771] <= 16'b0000_0000_0000_0000;
array[45772] <= 16'b0000_0000_0000_0000;
array[45773] <= 16'b0000_0000_0000_0000;
array[45774] <= 16'b0000_0000_0000_0000;
array[45775] <= 16'b0000_0000_0000_0000;
array[45776] <= 16'b0000_0000_0000_0000;
array[45777] <= 16'b0000_0000_0000_0000;
array[45778] <= 16'b0000_0000_0000_0000;
array[45779] <= 16'b0000_0000_0000_0000;
array[45780] <= 16'b0000_0000_0000_0000;
array[45781] <= 16'b0000_0000_0000_0000;
array[45782] <= 16'b0000_0000_0000_0000;
array[45783] <= 16'b0000_0000_0000_0000;
array[45784] <= 16'b0000_0000_0000_0000;
array[45785] <= 16'b0000_0000_0000_0000;
array[45786] <= 16'b0000_0000_0000_0000;
array[45787] <= 16'b0000_0000_0000_0000;
array[45788] <= 16'b0000_0000_0000_0000;
array[45789] <= 16'b0000_0000_0000_0000;
array[45790] <= 16'b0000_0000_0000_0000;
array[45791] <= 16'b0000_0000_0000_0000;
array[45792] <= 16'b0000_0000_0000_0000;
array[45793] <= 16'b0000_0000_0000_0000;
array[45794] <= 16'b0000_0000_0000_0000;
array[45795] <= 16'b0000_0000_0000_0000;
array[45796] <= 16'b0000_0000_0000_0000;
array[45797] <= 16'b0000_0000_0000_0000;
array[45798] <= 16'b0000_0000_0000_0000;
array[45799] <= 16'b0000_0000_0000_0000;
array[45800] <= 16'b0000_0000_0000_0000;
array[45801] <= 16'b0000_0000_0000_0000;
array[45802] <= 16'b0000_0000_0000_0000;
array[45803] <= 16'b0000_0000_0000_0000;
array[45804] <= 16'b0000_0000_0000_0000;
array[45805] <= 16'b0000_0000_0000_0000;
array[45806] <= 16'b0000_0000_0000_0000;
array[45807] <= 16'b0000_0000_0000_0000;
array[45808] <= 16'b0000_0000_0000_0000;
array[45809] <= 16'b0000_0000_0000_0000;
array[45810] <= 16'b0000_0000_0000_0000;
array[45811] <= 16'b0000_0000_0000_0000;
array[45812] <= 16'b0000_0000_0000_0000;
array[45813] <= 16'b0000_0000_0000_0000;
array[45814] <= 16'b0000_0000_0000_0000;
array[45815] <= 16'b0000_0000_0000_0000;
array[45816] <= 16'b0000_0000_0000_0000;
array[45817] <= 16'b0000_0000_0000_0000;
array[45818] <= 16'b0000_0000_0000_0000;
array[45819] <= 16'b0000_0000_0000_0000;
array[45820] <= 16'b0000_0000_0000_0000;
array[45821] <= 16'b0000_0000_0000_0000;
array[45822] <= 16'b0000_0000_0000_0000;
array[45823] <= 16'b0000_0000_0000_0000;
array[45824] <= 16'b0000_0000_0000_0000;
array[45825] <= 16'b0000_0000_0000_0000;
array[45826] <= 16'b0000_0000_0000_0000;
array[45827] <= 16'b0000_0000_0000_0000;
array[45828] <= 16'b0000_0000_0000_0000;
array[45829] <= 16'b0000_0000_0000_0000;
array[45830] <= 16'b0000_0000_0000_0000;
array[45831] <= 16'b0000_0000_0000_0000;
array[45832] <= 16'b0000_0000_0000_0000;
array[45833] <= 16'b0000_0000_0000_0000;
array[45834] <= 16'b0000_0000_0000_0000;
array[45835] <= 16'b0000_0000_0000_0000;
array[45836] <= 16'b0000_0000_0000_0000;
array[45837] <= 16'b0000_0000_0000_0000;
array[45838] <= 16'b0000_0000_0000_0000;
array[45839] <= 16'b0000_0000_0000_0000;
array[45840] <= 16'b0000_0000_0000_0000;
array[45841] <= 16'b0000_0000_0000_0000;
array[45842] <= 16'b0000_0000_0000_0000;
array[45843] <= 16'b0000_0000_0000_0000;
array[45844] <= 16'b0000_0000_0000_0000;
array[45845] <= 16'b0000_0000_0000_0000;
array[45846] <= 16'b0000_0000_0000_0000;
array[45847] <= 16'b0000_0000_0000_0000;
array[45848] <= 16'b0000_0000_0000_0000;
array[45849] <= 16'b0000_0000_0000_0000;
array[45850] <= 16'b0000_0000_0000_0000;
array[45851] <= 16'b0000_0000_0000_0000;
array[45852] <= 16'b0000_0000_0000_0000;
array[45853] <= 16'b0000_0000_0000_0000;
array[45854] <= 16'b0000_0000_0000_0000;
array[45855] <= 16'b0000_0000_0000_0000;
array[45856] <= 16'b0000_0000_0000_0000;
array[45857] <= 16'b0000_0000_0000_0000;
array[45858] <= 16'b0000_0000_0000_0000;
array[45859] <= 16'b0000_0000_0000_0000;
array[45860] <= 16'b0000_0000_0000_0000;
array[45861] <= 16'b0000_0000_0000_0000;
array[45862] <= 16'b0000_0000_0000_0000;
array[45863] <= 16'b0000_0000_0000_0000;
array[45864] <= 16'b0000_0000_0000_0000;
array[45865] <= 16'b0000_0000_0000_0000;
array[45866] <= 16'b0000_0000_0000_0000;
array[45867] <= 16'b0000_0000_0000_0000;
array[45868] <= 16'b0000_0000_0000_0000;
array[45869] <= 16'b0000_0000_0000_0000;
array[45870] <= 16'b0000_0000_0000_0000;
array[45871] <= 16'b0000_0000_0000_0000;
array[45872] <= 16'b0000_0000_0000_0000;
array[45873] <= 16'b0000_0000_0000_0000;
array[45874] <= 16'b0000_0000_0000_0000;
array[45875] <= 16'b0000_0000_0000_0000;
array[45876] <= 16'b0000_0000_0000_0000;
array[45877] <= 16'b0000_0000_0000_0000;
array[45878] <= 16'b0000_0000_0000_0000;
array[45879] <= 16'b0000_0000_0000_0000;
array[45880] <= 16'b0000_0000_0000_0000;
array[45881] <= 16'b0000_0000_0000_0000;
array[45882] <= 16'b0000_0000_0000_0000;
array[45883] <= 16'b0000_0000_0000_0000;
array[45884] <= 16'b0000_0000_0000_0000;
array[45885] <= 16'b0000_0000_0000_0000;
array[45886] <= 16'b0000_0000_0000_0000;
array[45887] <= 16'b0000_0000_0000_0000;
array[45888] <= 16'b0000_0000_0000_0000;
array[45889] <= 16'b0000_0000_0000_0000;
array[45890] <= 16'b0000_0000_0000_0000;
array[45891] <= 16'b0000_0000_0000_0000;
array[45892] <= 16'b0000_0000_0000_0000;
array[45893] <= 16'b0000_0000_0000_0000;
array[45894] <= 16'b0000_0000_0000_0000;
array[45895] <= 16'b0000_0000_0000_0000;
array[45896] <= 16'b0000_0000_0000_0000;
array[45897] <= 16'b0000_0000_0000_0000;
array[45898] <= 16'b0000_0000_0000_0000;
array[45899] <= 16'b0000_0000_0000_0000;
array[45900] <= 16'b0000_0000_0000_0000;
array[45901] <= 16'b0000_0000_0000_0000;
array[45902] <= 16'b0000_0000_0000_0000;
array[45903] <= 16'b0000_0000_0000_0000;
array[45904] <= 16'b0000_0000_0000_0000;
array[45905] <= 16'b0000_0000_0000_0000;
array[45906] <= 16'b0000_0000_0000_0000;
array[45907] <= 16'b0000_0000_0000_0000;
array[45908] <= 16'b0000_0000_0000_0000;
array[45909] <= 16'b0000_0000_0000_0000;
array[45910] <= 16'b0000_0000_0000_0000;
array[45911] <= 16'b0000_0000_0000_0000;
array[45912] <= 16'b0000_0000_0000_0000;
array[45913] <= 16'b0000_0000_0000_0000;
array[45914] <= 16'b0000_0000_0000_0000;
array[45915] <= 16'b0000_0000_0000_0000;
array[45916] <= 16'b0000_0000_0000_0000;
array[45917] <= 16'b0000_0000_0000_0000;
array[45918] <= 16'b0000_0000_0000_0000;
array[45919] <= 16'b0000_0000_0000_0000;
array[45920] <= 16'b0000_0000_0000_0000;
array[45921] <= 16'b0000_0000_0000_0000;
array[45922] <= 16'b0000_0000_0000_0000;
array[45923] <= 16'b0000_0000_0000_0000;
array[45924] <= 16'b0000_0000_0000_0000;
array[45925] <= 16'b0000_0000_0000_0000;
array[45926] <= 16'b0000_0000_0000_0000;
array[45927] <= 16'b0000_0000_0000_0000;
array[45928] <= 16'b0000_0000_0000_0000;
array[45929] <= 16'b0000_0000_0000_0000;
array[45930] <= 16'b0000_0000_0000_0000;
array[45931] <= 16'b0000_0000_0000_0000;
array[45932] <= 16'b0000_0000_0000_0000;
array[45933] <= 16'b0000_0000_0000_0000;
array[45934] <= 16'b0000_0000_0000_0000;
array[45935] <= 16'b0000_0000_0000_0000;
array[45936] <= 16'b0000_0000_0000_0000;
array[45937] <= 16'b0000_0000_0000_0000;
array[45938] <= 16'b0000_0000_0000_0000;
array[45939] <= 16'b0000_0000_0000_0000;
array[45940] <= 16'b0000_0000_0000_0000;
array[45941] <= 16'b0000_0000_0000_0000;
array[45942] <= 16'b0000_0000_0000_0000;
array[45943] <= 16'b0000_0000_0000_0000;
array[45944] <= 16'b0000_0000_0000_0000;
array[45945] <= 16'b0000_0000_0000_0000;
array[45946] <= 16'b0000_0000_0000_0000;
array[45947] <= 16'b0000_0000_0000_0000;
array[45948] <= 16'b0000_0000_0000_0000;
array[45949] <= 16'b0000_0000_0000_0000;
array[45950] <= 16'b0000_0000_0000_0000;
array[45951] <= 16'b0000_0000_0000_0000;
array[45952] <= 16'b0000_0000_0000_0000;
array[45953] <= 16'b0000_0000_0000_0000;
array[45954] <= 16'b0000_0000_0000_0000;
array[45955] <= 16'b0000_0000_0000_0000;
array[45956] <= 16'b0000_0000_0000_0000;
array[45957] <= 16'b0000_0000_0000_0000;
array[45958] <= 16'b0000_0000_0000_0000;
array[45959] <= 16'b0000_0000_0000_0000;
array[45960] <= 16'b0000_0000_0000_0000;
array[45961] <= 16'b0000_0000_0000_0000;
array[45962] <= 16'b0000_0000_0000_0000;
array[45963] <= 16'b0000_0000_0000_0000;
array[45964] <= 16'b0000_0000_0000_0000;
array[45965] <= 16'b0000_0000_0000_0000;
array[45966] <= 16'b0000_0000_0000_0000;
array[45967] <= 16'b0000_0000_0000_0000;
array[45968] <= 16'b0000_0000_0000_0000;
array[45969] <= 16'b0000_0000_0000_0000;
array[45970] <= 16'b0000_0000_0000_0000;
array[45971] <= 16'b0000_0000_0000_0000;
array[45972] <= 16'b0000_0000_0000_0000;
array[45973] <= 16'b0000_0000_0000_0000;
array[45974] <= 16'b0000_0000_0000_0000;
array[45975] <= 16'b0000_0000_0000_0000;
array[45976] <= 16'b0000_0000_0000_0000;
array[45977] <= 16'b0000_0000_0000_0000;
array[45978] <= 16'b0000_0000_0000_0000;
array[45979] <= 16'b0000_0000_0000_0000;
array[45980] <= 16'b0000_0000_0000_0000;
array[45981] <= 16'b0000_0000_0000_0000;
array[45982] <= 16'b0000_0000_0000_0000;
array[45983] <= 16'b0000_0000_0000_0000;
array[45984] <= 16'b0000_0000_0000_0000;
array[45985] <= 16'b0000_0000_0000_0000;
array[45986] <= 16'b0000_0000_0000_0000;
array[45987] <= 16'b0000_0000_0000_0000;
array[45988] <= 16'b0000_0000_0000_0000;
array[45989] <= 16'b0000_0000_0000_0000;
array[45990] <= 16'b0000_0000_0000_0000;
array[45991] <= 16'b0000_0000_0000_0000;
array[45992] <= 16'b0000_0000_0000_0000;
array[45993] <= 16'b0000_0000_0000_0000;
array[45994] <= 16'b0000_0000_0000_0000;
array[45995] <= 16'b0000_0000_0000_0000;
array[45996] <= 16'b0000_0000_0000_0000;
array[45997] <= 16'b0000_0000_0000_0000;
array[45998] <= 16'b0000_0000_0000_0000;
array[45999] <= 16'b0000_0000_0000_0000;
array[46000] <= 16'b0000_0000_0000_0000;
array[46001] <= 16'b0000_0000_0000_0000;
array[46002] <= 16'b0000_0000_0000_0000;
array[46003] <= 16'b0000_0000_0000_0000;
array[46004] <= 16'b0000_0000_0000_0000;
array[46005] <= 16'b0000_0000_0000_0000;
array[46006] <= 16'b0000_0000_0000_0000;
array[46007] <= 16'b0000_0000_0000_0000;
array[46008] <= 16'b0000_0000_0000_0000;
array[46009] <= 16'b0000_0000_0000_0000;
array[46010] <= 16'b0000_0000_0000_0000;
array[46011] <= 16'b0000_0000_0000_0000;
array[46012] <= 16'b0000_0000_0000_0000;
array[46013] <= 16'b0000_0000_0000_0000;
array[46014] <= 16'b0000_0000_0000_0000;
array[46015] <= 16'b0000_0000_0000_0000;
array[46016] <= 16'b0000_0000_0000_0000;
array[46017] <= 16'b0000_0000_0000_0000;
array[46018] <= 16'b0000_0000_0000_0000;
array[46019] <= 16'b0000_0000_0000_0000;
array[46020] <= 16'b0000_0000_0000_0000;
array[46021] <= 16'b0000_0000_0000_0000;
array[46022] <= 16'b0000_0000_0000_0000;
array[46023] <= 16'b0000_0000_0000_0000;
array[46024] <= 16'b0000_0000_0000_0000;
array[46025] <= 16'b0000_0000_0000_0000;
array[46026] <= 16'b0000_0000_0000_0000;
array[46027] <= 16'b0000_0000_0000_0000;
array[46028] <= 16'b0000_0000_0000_0000;
array[46029] <= 16'b0000_0000_0000_0000;
array[46030] <= 16'b0000_0000_0000_0000;
array[46031] <= 16'b0000_0000_0000_0000;
array[46032] <= 16'b0000_0000_0000_0000;
array[46033] <= 16'b0000_0000_0000_0000;
array[46034] <= 16'b0000_0000_0000_0000;
array[46035] <= 16'b0000_0000_0000_0000;
array[46036] <= 16'b0000_0000_0000_0000;
array[46037] <= 16'b0000_0000_0000_0000;
array[46038] <= 16'b0000_0000_0000_0000;
array[46039] <= 16'b0000_0000_0000_0000;
array[46040] <= 16'b0000_0000_0000_0000;
array[46041] <= 16'b0000_0000_0000_0000;
array[46042] <= 16'b0000_0000_0000_0000;
array[46043] <= 16'b0000_0000_0000_0000;
array[46044] <= 16'b0000_0000_0000_0000;
array[46045] <= 16'b0000_0000_0000_0000;
array[46046] <= 16'b0000_0000_0000_0000;
array[46047] <= 16'b0000_0000_0000_0000;
array[46048] <= 16'b0000_0000_0000_0000;
array[46049] <= 16'b0000_0000_0000_0000;
array[46050] <= 16'b0000_0000_0000_0000;
array[46051] <= 16'b0000_0000_0000_0000;
array[46052] <= 16'b0000_0000_0000_0000;
array[46053] <= 16'b0000_0000_0000_0000;
array[46054] <= 16'b0000_0000_0000_0000;
array[46055] <= 16'b0000_0000_0000_0000;
array[46056] <= 16'b0000_0000_0000_0000;
array[46057] <= 16'b0000_0000_0000_0000;
array[46058] <= 16'b0000_0000_0000_0000;
array[46059] <= 16'b0000_0000_0000_0000;
array[46060] <= 16'b0000_0000_0000_0000;
array[46061] <= 16'b0000_0000_0000_0000;
array[46062] <= 16'b0000_0000_0000_0000;
array[46063] <= 16'b0000_0000_0000_0000;
array[46064] <= 16'b0000_0000_0000_0000;
array[46065] <= 16'b0000_0000_0000_0000;
array[46066] <= 16'b0000_0000_0000_0000;
array[46067] <= 16'b0000_0000_0000_0000;
array[46068] <= 16'b0000_0000_0000_0000;
array[46069] <= 16'b0000_0000_0000_0000;
array[46070] <= 16'b0000_0000_0000_0000;
array[46071] <= 16'b0000_0000_0000_0000;
array[46072] <= 16'b0000_0000_0000_0000;
array[46073] <= 16'b0000_0000_0000_0000;
array[46074] <= 16'b0000_0000_0000_0000;
array[46075] <= 16'b0000_0000_0000_0000;
array[46076] <= 16'b0000_0000_0000_0000;
array[46077] <= 16'b0000_0000_0000_0000;
array[46078] <= 16'b0000_0000_0000_0000;
array[46079] <= 16'b0000_0000_0000_0000;
array[46080] <= 16'b0000_0000_0000_0000;
array[46081] <= 16'b0000_0000_0000_0000;
array[46082] <= 16'b0000_0000_0000_0000;
array[46083] <= 16'b0000_0000_0000_0000;
array[46084] <= 16'b0000_0000_0000_0000;
array[46085] <= 16'b0000_0000_0000_0000;
array[46086] <= 16'b0000_0000_0000_0000;
array[46087] <= 16'b0000_0000_0000_0000;
array[46088] <= 16'b0000_0000_0000_0000;
array[46089] <= 16'b0000_0000_0000_0000;
array[46090] <= 16'b0000_0000_0000_0000;
array[46091] <= 16'b0000_0000_0000_0000;
array[46092] <= 16'b0000_0000_0000_0000;
array[46093] <= 16'b0000_0000_0000_0000;
array[46094] <= 16'b0000_0000_0000_0000;
array[46095] <= 16'b0000_0000_0000_0000;
array[46096] <= 16'b0000_0000_0000_0000;
array[46097] <= 16'b0000_0000_0000_0000;
array[46098] <= 16'b0000_0000_0000_0000;
array[46099] <= 16'b0000_0000_0000_0000;
array[46100] <= 16'b0000_0000_0000_0000;
array[46101] <= 16'b0000_0000_0000_0000;
array[46102] <= 16'b0000_0000_0000_0000;
array[46103] <= 16'b0000_0000_0000_0000;
array[46104] <= 16'b0000_0000_0000_0000;
array[46105] <= 16'b0000_0000_0000_0000;
array[46106] <= 16'b0000_0000_0000_0000;
array[46107] <= 16'b0000_0000_0000_0000;
array[46108] <= 16'b0000_0000_0000_0000;
array[46109] <= 16'b0000_0000_0000_0000;
array[46110] <= 16'b0000_0000_0000_0000;
array[46111] <= 16'b0000_0000_0000_0000;
array[46112] <= 16'b0000_0000_0000_0000;
array[46113] <= 16'b0000_0000_0000_0000;
array[46114] <= 16'b0000_0000_0000_0000;
array[46115] <= 16'b0000_0000_0000_0000;
array[46116] <= 16'b0000_0000_0000_0000;
array[46117] <= 16'b0000_0000_0000_0000;
array[46118] <= 16'b0000_0000_0000_0000;
array[46119] <= 16'b0000_0000_0000_0000;
array[46120] <= 16'b0000_0000_0000_0000;
array[46121] <= 16'b0000_0000_0000_0000;
array[46122] <= 16'b0000_0000_0000_0000;
array[46123] <= 16'b0000_0000_0000_0000;
array[46124] <= 16'b0000_0000_0000_0000;
array[46125] <= 16'b0000_0000_0000_0000;
array[46126] <= 16'b0000_0000_0000_0000;
array[46127] <= 16'b0000_0000_0000_0000;
array[46128] <= 16'b0000_0000_0000_0000;
array[46129] <= 16'b0000_0000_0000_0000;
array[46130] <= 16'b0000_0000_0000_0000;
array[46131] <= 16'b0000_0000_0000_0000;
array[46132] <= 16'b0000_0000_0000_0000;
array[46133] <= 16'b0000_0000_0000_0000;
array[46134] <= 16'b0000_0000_0000_0000;
array[46135] <= 16'b0000_0000_0000_0000;
array[46136] <= 16'b0000_0000_0000_0000;
array[46137] <= 16'b0000_0000_0000_0000;
array[46138] <= 16'b0000_0000_0000_0000;
array[46139] <= 16'b0000_0000_0000_0000;
array[46140] <= 16'b0000_0000_0000_0000;
array[46141] <= 16'b0000_0000_0000_0000;
array[46142] <= 16'b0000_0000_0000_0000;
array[46143] <= 16'b0000_0000_0000_0000;
array[46144] <= 16'b0000_0000_0000_0000;
array[46145] <= 16'b0000_0000_0000_0000;
array[46146] <= 16'b0000_0000_0000_0000;
array[46147] <= 16'b0000_0000_0000_0000;
array[46148] <= 16'b0000_0000_0000_0000;
array[46149] <= 16'b0000_0000_0000_0000;
array[46150] <= 16'b0000_0000_0000_0000;
array[46151] <= 16'b0000_0000_0000_0000;
array[46152] <= 16'b0000_0000_0000_0000;
array[46153] <= 16'b0000_0000_0000_0000;
array[46154] <= 16'b0000_0000_0000_0000;
array[46155] <= 16'b0000_0000_0000_0000;
array[46156] <= 16'b0000_0000_0000_0000;
array[46157] <= 16'b0000_0000_0000_0000;
array[46158] <= 16'b0000_0000_0000_0000;
array[46159] <= 16'b0000_0000_0000_0000;
array[46160] <= 16'b0000_0000_0000_0000;
array[46161] <= 16'b0000_0000_0000_0000;
array[46162] <= 16'b0000_0000_0000_0000;
array[46163] <= 16'b0000_0000_0000_0000;
array[46164] <= 16'b0000_0000_0000_0000;
array[46165] <= 16'b0000_0000_0000_0000;
array[46166] <= 16'b0000_0000_0000_0000;
array[46167] <= 16'b0000_0000_0000_0000;
array[46168] <= 16'b0000_0000_0000_0000;
array[46169] <= 16'b0000_0000_0000_0000;
array[46170] <= 16'b0000_0000_0000_0000;
array[46171] <= 16'b0000_0000_0000_0000;
array[46172] <= 16'b0000_0000_0000_0000;
array[46173] <= 16'b0000_0000_0000_0000;
array[46174] <= 16'b0000_0000_0000_0000;
array[46175] <= 16'b0000_0000_0000_0000;
array[46176] <= 16'b0000_0000_0000_0000;
array[46177] <= 16'b0000_0000_0000_0000;
array[46178] <= 16'b0000_0000_0000_0000;
array[46179] <= 16'b0000_0000_0000_0000;
array[46180] <= 16'b0000_0000_0000_0000;
array[46181] <= 16'b0000_0000_0000_0000;
array[46182] <= 16'b0000_0000_0000_0000;
array[46183] <= 16'b0000_0000_0000_0000;
array[46184] <= 16'b0000_0000_0000_0000;
array[46185] <= 16'b0000_0000_0000_0000;
array[46186] <= 16'b0000_0000_0000_0000;
array[46187] <= 16'b0000_0000_0000_0000;
array[46188] <= 16'b0000_0000_0000_0000;
array[46189] <= 16'b0000_0000_0000_0000;
array[46190] <= 16'b0000_0000_0000_0000;
array[46191] <= 16'b0000_0000_0000_0000;
array[46192] <= 16'b0000_0000_0000_0000;
array[46193] <= 16'b0000_0000_0000_0000;
array[46194] <= 16'b0000_0000_0000_0000;
array[46195] <= 16'b0000_0000_0000_0000;
array[46196] <= 16'b0000_0000_0000_0000;
array[46197] <= 16'b0000_0000_0000_0000;
array[46198] <= 16'b0000_0000_0000_0000;
array[46199] <= 16'b0000_0000_0000_0000;
array[46200] <= 16'b0000_0000_0000_0000;
array[46201] <= 16'b0000_0000_0000_0000;
array[46202] <= 16'b0000_0000_0000_0000;
array[46203] <= 16'b0000_0000_0000_0000;
array[46204] <= 16'b0000_0000_0000_0000;
array[46205] <= 16'b0000_0000_0000_0000;
array[46206] <= 16'b0000_0000_0000_0000;
array[46207] <= 16'b0000_0000_0000_0000;
array[46208] <= 16'b0000_0000_0000_0000;
array[46209] <= 16'b0000_0000_0000_0000;
array[46210] <= 16'b0000_0000_0000_0000;
array[46211] <= 16'b0000_0000_0000_0000;
array[46212] <= 16'b0000_0000_0000_0000;
array[46213] <= 16'b0000_0000_0000_0000;
array[46214] <= 16'b0000_0000_0000_0000;
array[46215] <= 16'b0000_0000_0000_0000;
array[46216] <= 16'b0000_0000_0000_0000;
array[46217] <= 16'b0000_0000_0000_0000;
array[46218] <= 16'b0000_0000_0000_0000;
array[46219] <= 16'b0000_0000_0000_0000;
array[46220] <= 16'b0000_0000_0000_0000;
array[46221] <= 16'b0000_0000_0000_0000;
array[46222] <= 16'b0000_0000_0000_0000;
array[46223] <= 16'b0000_0000_0000_0000;
array[46224] <= 16'b0000_0000_0000_0000;
array[46225] <= 16'b0000_0000_0000_0000;
array[46226] <= 16'b0000_0000_0000_0000;
array[46227] <= 16'b0000_0000_0000_0000;
array[46228] <= 16'b0000_0000_0000_0000;
array[46229] <= 16'b0000_0000_0000_0000;
array[46230] <= 16'b0000_0000_0000_0000;
array[46231] <= 16'b0000_0000_0000_0000;
array[46232] <= 16'b0000_0000_0000_0000;
array[46233] <= 16'b0000_0000_0000_0000;
array[46234] <= 16'b0000_0000_0000_0000;
array[46235] <= 16'b0000_0000_0000_0000;
array[46236] <= 16'b0000_0000_0000_0000;
array[46237] <= 16'b0000_0000_0000_0000;
array[46238] <= 16'b0000_0000_0000_0000;
array[46239] <= 16'b0000_0000_0000_0000;
array[46240] <= 16'b0000_0000_0000_0000;
array[46241] <= 16'b0000_0000_0000_0000;
array[46242] <= 16'b0000_0000_0000_0000;
array[46243] <= 16'b0000_0000_0000_0000;
array[46244] <= 16'b0000_0000_0000_0000;
array[46245] <= 16'b0000_0000_0000_0000;
array[46246] <= 16'b0000_0000_0000_0000;
array[46247] <= 16'b0000_0000_0000_0000;
array[46248] <= 16'b0000_0000_0000_0000;
array[46249] <= 16'b0000_0000_0000_0000;
array[46250] <= 16'b0000_0000_0000_0000;
array[46251] <= 16'b0000_0000_0000_0000;
array[46252] <= 16'b0000_0000_0000_0000;
array[46253] <= 16'b0000_0000_0000_0000;
array[46254] <= 16'b0000_0000_0000_0000;
array[46255] <= 16'b0000_0000_0000_0000;
array[46256] <= 16'b0000_0000_0000_0000;
array[46257] <= 16'b0000_0000_0000_0000;
array[46258] <= 16'b0000_0000_0000_0000;
array[46259] <= 16'b0000_0000_0000_0000;
array[46260] <= 16'b0000_0000_0000_0000;
array[46261] <= 16'b0000_0000_0000_0000;
array[46262] <= 16'b0000_0000_0000_0000;
array[46263] <= 16'b0000_0000_0000_0000;
array[46264] <= 16'b0000_0000_0000_0000;
array[46265] <= 16'b0000_0000_0000_0000;
array[46266] <= 16'b0000_0000_0000_0000;
array[46267] <= 16'b0000_0000_0000_0000;
array[46268] <= 16'b0000_0000_0000_0000;
array[46269] <= 16'b0000_0000_0000_0000;
array[46270] <= 16'b0000_0000_0000_0000;
array[46271] <= 16'b0000_0000_0000_0000;
array[46272] <= 16'b0000_0000_0000_0000;
array[46273] <= 16'b0000_0000_0000_0000;
array[46274] <= 16'b0000_0000_0000_0000;
array[46275] <= 16'b0000_0000_0000_0000;
array[46276] <= 16'b0000_0000_0000_0000;
array[46277] <= 16'b0000_0000_0000_0000;
array[46278] <= 16'b0000_0000_0000_0000;
array[46279] <= 16'b0000_0000_0000_0000;
array[46280] <= 16'b0000_0000_0000_0000;
array[46281] <= 16'b0000_0000_0000_0000;
array[46282] <= 16'b0000_0000_0000_0000;
array[46283] <= 16'b0000_0000_0000_0000;
array[46284] <= 16'b0000_0000_0000_0000;
array[46285] <= 16'b0000_0000_0000_0000;
array[46286] <= 16'b0000_0000_0000_0000;
array[46287] <= 16'b0000_0000_0000_0000;
array[46288] <= 16'b0000_0000_0000_0000;
array[46289] <= 16'b0000_0000_0000_0000;
array[46290] <= 16'b0000_0000_0000_0000;
array[46291] <= 16'b0000_0000_0000_0000;
array[46292] <= 16'b0000_0000_0000_0000;
array[46293] <= 16'b0000_0000_0000_0000;
array[46294] <= 16'b0000_0000_0000_0000;
array[46295] <= 16'b0000_0000_0000_0000;
array[46296] <= 16'b0000_0000_0000_0000;
array[46297] <= 16'b0000_0000_0000_0000;
array[46298] <= 16'b0000_0000_0000_0000;
array[46299] <= 16'b0000_0000_0000_0000;
array[46300] <= 16'b0000_0000_0000_0000;
array[46301] <= 16'b0000_0000_0000_0000;
array[46302] <= 16'b0000_0000_0000_0000;
array[46303] <= 16'b0000_0000_0000_0000;
array[46304] <= 16'b0000_0000_0000_0000;
array[46305] <= 16'b0000_0000_0000_0000;
array[46306] <= 16'b0000_0000_0000_0000;
array[46307] <= 16'b0000_0000_0000_0000;
array[46308] <= 16'b0000_0000_0000_0000;
array[46309] <= 16'b0000_0000_0000_0000;
array[46310] <= 16'b0000_0000_0000_0000;
array[46311] <= 16'b0000_0000_0000_0000;
array[46312] <= 16'b0000_0000_0000_0000;
array[46313] <= 16'b0000_0000_0000_0000;
array[46314] <= 16'b0000_0000_0000_0000;
array[46315] <= 16'b0000_0000_0000_0000;
array[46316] <= 16'b0000_0000_0000_0000;
array[46317] <= 16'b0000_0000_0000_0000;
array[46318] <= 16'b0000_0000_0000_0000;
array[46319] <= 16'b0000_0000_0000_0000;
array[46320] <= 16'b0000_0000_0000_0000;
array[46321] <= 16'b0000_0000_0000_0000;
array[46322] <= 16'b0000_0000_0000_0000;
array[46323] <= 16'b0000_0000_0000_0000;
array[46324] <= 16'b0000_0000_0000_0000;
array[46325] <= 16'b0000_0000_0000_0000;
array[46326] <= 16'b0000_0000_0000_0000;
array[46327] <= 16'b0000_0000_0000_0000;
array[46328] <= 16'b0000_0000_0000_0000;
array[46329] <= 16'b0000_0000_0000_0000;
array[46330] <= 16'b0000_0000_0000_0000;
array[46331] <= 16'b0000_0000_0000_0000;
array[46332] <= 16'b0000_0000_0000_0000;
array[46333] <= 16'b0000_0000_0000_0000;
array[46334] <= 16'b0000_0000_0000_0000;
array[46335] <= 16'b0000_0000_0000_0000;
array[46336] <= 16'b0000_0000_0000_0000;
array[46337] <= 16'b0000_0000_0000_0000;
array[46338] <= 16'b0000_0000_0000_0000;
array[46339] <= 16'b0000_0000_0000_0000;
array[46340] <= 16'b0000_0000_0000_0000;
array[46341] <= 16'b0000_0000_0000_0000;
array[46342] <= 16'b0000_0000_0000_0000;
array[46343] <= 16'b0000_0000_0000_0000;
array[46344] <= 16'b0000_0000_0000_0000;
array[46345] <= 16'b0000_0000_0000_0000;
array[46346] <= 16'b0000_0000_0000_0000;
array[46347] <= 16'b0000_0000_0000_0000;
array[46348] <= 16'b0000_0000_0000_0000;
array[46349] <= 16'b0000_0000_0000_0000;
array[46350] <= 16'b0000_0000_0000_0000;
array[46351] <= 16'b0000_0000_0000_0000;
array[46352] <= 16'b0000_0000_0000_0000;
array[46353] <= 16'b0000_0000_0000_0000;
array[46354] <= 16'b0000_0000_0000_0000;
array[46355] <= 16'b0000_0000_0000_0000;
array[46356] <= 16'b0000_0000_0000_0000;
array[46357] <= 16'b0000_0000_0000_0000;
array[46358] <= 16'b0000_0000_0000_0000;
array[46359] <= 16'b0000_0000_0000_0000;
array[46360] <= 16'b0000_0000_0000_0000;
array[46361] <= 16'b0000_0000_0000_0000;
array[46362] <= 16'b0000_0000_0000_0000;
array[46363] <= 16'b0000_0000_0000_0000;
array[46364] <= 16'b0000_0000_0000_0000;
array[46365] <= 16'b0000_0000_0000_0000;
array[46366] <= 16'b0000_0000_0000_0000;
array[46367] <= 16'b0000_0000_0000_0000;
array[46368] <= 16'b0000_0000_0000_0000;
array[46369] <= 16'b0000_0000_0000_0000;
array[46370] <= 16'b0000_0000_0000_0000;
array[46371] <= 16'b0000_0000_0000_0000;
array[46372] <= 16'b0000_0000_0000_0000;
array[46373] <= 16'b0000_0000_0000_0000;
array[46374] <= 16'b0000_0000_0000_0000;
array[46375] <= 16'b0000_0000_0000_0000;
array[46376] <= 16'b0000_0000_0000_0000;
array[46377] <= 16'b0000_0000_0000_0000;
array[46378] <= 16'b0000_0000_0000_0000;
array[46379] <= 16'b0000_0000_0000_0000;
array[46380] <= 16'b0000_0000_0000_0000;
array[46381] <= 16'b0000_0000_0000_0000;
array[46382] <= 16'b0000_0000_0000_0000;
array[46383] <= 16'b0000_0000_0000_0000;
array[46384] <= 16'b0000_0000_0000_0000;
array[46385] <= 16'b0000_0000_0000_0000;
array[46386] <= 16'b0000_0000_0000_0000;
array[46387] <= 16'b0000_0000_0000_0000;
array[46388] <= 16'b0000_0000_0000_0000;
array[46389] <= 16'b0000_0000_0000_0000;
array[46390] <= 16'b0000_0000_0000_0000;
array[46391] <= 16'b0000_0000_0000_0000;
array[46392] <= 16'b0000_0000_0000_0000;
array[46393] <= 16'b0000_0000_0000_0000;
array[46394] <= 16'b0000_0000_0000_0000;
array[46395] <= 16'b0000_0000_0000_0000;
array[46396] <= 16'b0000_0000_0000_0000;
array[46397] <= 16'b0000_0000_0000_0000;
array[46398] <= 16'b0000_0000_0000_0000;
array[46399] <= 16'b0000_0000_0000_0000;
array[46400] <= 16'b0000_0000_0000_0000;
array[46401] <= 16'b0000_0000_0000_0000;
array[46402] <= 16'b0000_0000_0000_0000;
array[46403] <= 16'b0000_0000_0000_0000;
array[46404] <= 16'b0000_0000_0000_0000;
array[46405] <= 16'b0000_0000_0000_0000;
array[46406] <= 16'b0000_0000_0000_0000;
array[46407] <= 16'b0000_0000_0000_0000;
array[46408] <= 16'b0000_0000_0000_0000;
array[46409] <= 16'b0000_0000_0000_0000;
array[46410] <= 16'b0000_0000_0000_0000;
array[46411] <= 16'b0000_0000_0000_0000;
array[46412] <= 16'b0000_0000_0000_0000;
array[46413] <= 16'b0000_0000_0000_0000;
array[46414] <= 16'b0000_0000_0000_0000;
array[46415] <= 16'b0000_0000_0000_0000;
array[46416] <= 16'b0000_0000_0000_0000;
array[46417] <= 16'b0000_0000_0000_0000;
array[46418] <= 16'b0000_0000_0000_0000;
array[46419] <= 16'b0000_0000_0000_0000;
array[46420] <= 16'b0000_0000_0000_0000;
array[46421] <= 16'b0000_0000_0000_0000;
array[46422] <= 16'b0000_0000_0000_0000;
array[46423] <= 16'b0000_0000_0000_0000;
array[46424] <= 16'b0000_0000_0000_0000;
array[46425] <= 16'b0000_0000_0000_0000;
array[46426] <= 16'b0000_0000_0000_0000;
array[46427] <= 16'b0000_0000_0000_0000;
array[46428] <= 16'b0000_0000_0000_0000;
array[46429] <= 16'b0000_0000_0000_0000;
array[46430] <= 16'b0000_0000_0000_0000;
array[46431] <= 16'b0000_0000_0000_0000;
array[46432] <= 16'b0000_0000_0000_0000;
array[46433] <= 16'b0000_0000_0000_0000;
array[46434] <= 16'b0000_0000_0000_0000;
array[46435] <= 16'b0000_0000_0000_0000;
array[46436] <= 16'b0000_0000_0000_0000;
array[46437] <= 16'b0000_0000_0000_0000;
array[46438] <= 16'b0000_0000_0000_0000;
array[46439] <= 16'b0000_0000_0000_0000;
array[46440] <= 16'b0000_0000_0000_0000;
array[46441] <= 16'b0000_0000_0000_0000;
array[46442] <= 16'b0000_0000_0000_0000;
array[46443] <= 16'b0000_0000_0000_0000;
array[46444] <= 16'b0000_0000_0000_0000;
array[46445] <= 16'b0000_0000_0000_0000;
array[46446] <= 16'b0000_0000_0000_0000;
array[46447] <= 16'b0000_0000_0000_0000;
array[46448] <= 16'b0000_0000_0000_0000;
array[46449] <= 16'b0000_0000_0000_0000;
array[46450] <= 16'b0000_0000_0000_0000;
array[46451] <= 16'b0000_0000_0000_0000;
array[46452] <= 16'b0000_0000_0000_0000;
array[46453] <= 16'b0000_0000_0000_0000;
array[46454] <= 16'b0000_0000_0000_0000;
array[46455] <= 16'b0000_0000_0000_0000;
array[46456] <= 16'b0000_0000_0000_0000;
array[46457] <= 16'b0000_0000_0000_0000;
array[46458] <= 16'b0000_0000_0000_0000;
array[46459] <= 16'b0000_0000_0000_0000;
array[46460] <= 16'b0000_0000_0000_0000;
array[46461] <= 16'b0000_0000_0000_0000;
array[46462] <= 16'b0000_0000_0000_0000;
array[46463] <= 16'b0000_0000_0000_0000;
array[46464] <= 16'b0000_0000_0000_0000;
array[46465] <= 16'b0000_0000_0000_0000;
array[46466] <= 16'b0000_0000_0000_0000;
array[46467] <= 16'b0000_0000_0000_0000;
array[46468] <= 16'b0000_0000_0000_0000;
array[46469] <= 16'b0000_0000_0000_0000;
array[46470] <= 16'b0000_0000_0000_0000;
array[46471] <= 16'b0000_0000_0000_0000;
array[46472] <= 16'b0000_0000_0000_0000;
array[46473] <= 16'b0000_0000_0000_0000;
array[46474] <= 16'b0000_0000_0000_0000;
array[46475] <= 16'b0000_0000_0000_0000;
array[46476] <= 16'b0000_0000_0000_0000;
array[46477] <= 16'b0000_0000_0000_0000;
array[46478] <= 16'b0000_0000_0000_0000;
array[46479] <= 16'b0000_0000_0000_0000;
array[46480] <= 16'b0000_0000_0000_0000;
array[46481] <= 16'b0000_0000_0000_0000;
array[46482] <= 16'b0000_0000_0000_0000;
array[46483] <= 16'b0000_0000_0000_0000;
array[46484] <= 16'b0000_0000_0000_0000;
array[46485] <= 16'b0000_0000_0000_0000;
array[46486] <= 16'b0000_0000_0000_0000;
array[46487] <= 16'b0000_0000_0000_0000;
array[46488] <= 16'b0000_0000_0000_0000;
array[46489] <= 16'b0000_0000_0000_0000;
array[46490] <= 16'b0000_0000_0000_0000;
array[46491] <= 16'b0000_0000_0000_0000;
array[46492] <= 16'b0000_0000_0000_0000;
array[46493] <= 16'b0000_0000_0000_0000;
array[46494] <= 16'b0000_0000_0000_0000;
array[46495] <= 16'b0000_0000_0000_0000;
array[46496] <= 16'b0000_0000_0000_0000;
array[46497] <= 16'b0000_0000_0000_0000;
array[46498] <= 16'b0000_0000_0000_0000;
array[46499] <= 16'b0000_0000_0000_0000;
array[46500] <= 16'b0000_0000_0000_0000;
array[46501] <= 16'b0000_0000_0000_0000;
array[46502] <= 16'b0000_0000_0000_0000;
array[46503] <= 16'b0000_0000_0000_0000;
array[46504] <= 16'b0000_0000_0000_0000;
array[46505] <= 16'b0000_0000_0000_0000;
array[46506] <= 16'b0000_0000_0000_0000;
array[46507] <= 16'b0000_0000_0000_0000;
array[46508] <= 16'b0000_0000_0000_0000;
array[46509] <= 16'b0000_0000_0000_0000;
array[46510] <= 16'b0000_0000_0000_0000;
array[46511] <= 16'b0000_0000_0000_0000;
array[46512] <= 16'b0000_0000_0000_0000;
array[46513] <= 16'b0000_0000_0000_0000;
array[46514] <= 16'b0000_0000_0000_0000;
array[46515] <= 16'b0000_0000_0000_0000;
array[46516] <= 16'b0000_0000_0000_0000;
array[46517] <= 16'b0000_0000_0000_0000;
array[46518] <= 16'b0000_0000_0000_0000;
array[46519] <= 16'b0000_0000_0000_0000;
array[46520] <= 16'b0000_0000_0000_0000;
array[46521] <= 16'b0000_0000_0000_0000;
array[46522] <= 16'b0000_0000_0000_0000;
array[46523] <= 16'b0000_0000_0000_0000;
array[46524] <= 16'b0000_0000_0000_0000;
array[46525] <= 16'b0000_0000_0000_0000;
array[46526] <= 16'b0000_0000_0000_0000;
array[46527] <= 16'b0000_0000_0000_0000;
array[46528] <= 16'b0000_0000_0000_0000;
array[46529] <= 16'b0000_0000_0000_0000;
array[46530] <= 16'b0000_0000_0000_0000;
array[46531] <= 16'b0000_0000_0000_0000;
array[46532] <= 16'b0000_0000_0000_0000;
array[46533] <= 16'b0000_0000_0000_0000;
array[46534] <= 16'b0000_0000_0000_0000;
array[46535] <= 16'b0000_0000_0000_0000;
array[46536] <= 16'b0000_0000_0000_0000;
array[46537] <= 16'b0000_0000_0000_0000;
array[46538] <= 16'b0000_0000_0000_0000;
array[46539] <= 16'b0000_0000_0000_0000;
array[46540] <= 16'b0000_0000_0000_0000;
array[46541] <= 16'b0000_0000_0000_0000;
array[46542] <= 16'b0000_0000_0000_0000;
array[46543] <= 16'b0000_0000_0000_0000;
array[46544] <= 16'b0000_0000_0000_0000;
array[46545] <= 16'b0000_0000_0000_0000;
array[46546] <= 16'b0000_0000_0000_0000;
array[46547] <= 16'b0000_0000_0000_0000;
array[46548] <= 16'b0000_0000_0000_0000;
array[46549] <= 16'b0000_0000_0000_0000;
array[46550] <= 16'b0000_0000_0000_0000;
array[46551] <= 16'b0000_0000_0000_0000;
array[46552] <= 16'b0000_0000_0000_0000;
array[46553] <= 16'b0000_0000_0000_0000;
array[46554] <= 16'b0000_0000_0000_0000;
array[46555] <= 16'b0000_0000_0000_0000;
array[46556] <= 16'b0000_0000_0000_0000;
array[46557] <= 16'b0000_0000_0000_0000;
array[46558] <= 16'b0000_0000_0000_0000;
array[46559] <= 16'b0000_0000_0000_0000;
array[46560] <= 16'b0000_0000_0000_0000;
array[46561] <= 16'b0000_0000_0000_0000;
array[46562] <= 16'b0000_0000_0000_0000;
array[46563] <= 16'b0000_0000_0000_0000;
array[46564] <= 16'b0000_0000_0000_0000;
array[46565] <= 16'b0000_0000_0000_0000;
array[46566] <= 16'b0000_0000_0000_0000;
array[46567] <= 16'b0000_0000_0000_0000;
array[46568] <= 16'b0000_0000_0000_0000;
array[46569] <= 16'b0000_0000_0000_0000;
array[46570] <= 16'b0000_0000_0000_0000;
array[46571] <= 16'b0000_0000_0000_0000;
array[46572] <= 16'b0000_0000_0000_0000;
array[46573] <= 16'b0000_0000_0000_0000;
array[46574] <= 16'b0000_0000_0000_0000;
array[46575] <= 16'b0000_0000_0000_0000;
array[46576] <= 16'b0000_0000_0000_0000;
array[46577] <= 16'b0000_0000_0000_0000;
array[46578] <= 16'b0000_0000_0000_0000;
array[46579] <= 16'b0000_0000_0000_0000;
array[46580] <= 16'b0000_0000_0000_0000;
array[46581] <= 16'b0000_0000_0000_0000;
array[46582] <= 16'b0000_0000_0000_0000;
array[46583] <= 16'b0000_0000_0000_0000;
array[46584] <= 16'b0000_0000_0000_0000;
array[46585] <= 16'b0000_0000_0000_0000;
array[46586] <= 16'b0000_0000_0000_0000;
array[46587] <= 16'b0000_0000_0000_0000;
array[46588] <= 16'b0000_0000_0000_0000;
array[46589] <= 16'b0000_0000_0000_0000;
array[46590] <= 16'b0000_0000_0000_0000;
array[46591] <= 16'b0000_0000_0000_0000;
array[46592] <= 16'b0000_0000_0000_0000;
array[46593] <= 16'b0000_0000_0000_0000;
array[46594] <= 16'b0000_0000_0000_0000;
array[46595] <= 16'b0000_0000_0000_0000;
array[46596] <= 16'b0000_0000_0000_0000;
array[46597] <= 16'b0000_0000_0000_0000;
array[46598] <= 16'b0000_0000_0000_0000;
array[46599] <= 16'b0000_0000_0000_0000;
array[46600] <= 16'b0000_0000_0000_0000;
array[46601] <= 16'b0000_0000_0000_0000;
array[46602] <= 16'b0000_0000_0000_0000;
array[46603] <= 16'b0000_0000_0000_0000;
array[46604] <= 16'b0000_0000_0000_0000;
array[46605] <= 16'b0000_0000_0000_0000;
array[46606] <= 16'b0000_0000_0000_0000;
array[46607] <= 16'b0000_0000_0000_0000;
array[46608] <= 16'b0000_0000_0000_0000;
array[46609] <= 16'b0000_0000_0000_0000;
array[46610] <= 16'b0000_0000_0000_0000;
array[46611] <= 16'b0000_0000_0000_0000;
array[46612] <= 16'b0000_0000_0000_0000;
array[46613] <= 16'b0000_0000_0000_0000;
array[46614] <= 16'b0000_0000_0000_0000;
array[46615] <= 16'b0000_0000_0000_0000;
array[46616] <= 16'b0000_0000_0000_0000;
array[46617] <= 16'b0000_0000_0000_0000;
array[46618] <= 16'b0000_0000_0000_0000;
array[46619] <= 16'b0000_0000_0000_0000;
array[46620] <= 16'b0000_0000_0000_0000;
array[46621] <= 16'b0000_0000_0000_0000;
array[46622] <= 16'b0000_0000_0000_0000;
array[46623] <= 16'b0000_0000_0000_0000;
array[46624] <= 16'b0000_0000_0000_0000;
array[46625] <= 16'b0000_0000_0000_0000;
array[46626] <= 16'b0000_0000_0000_0000;
array[46627] <= 16'b0000_0000_0000_0000;
array[46628] <= 16'b0000_0000_0000_0000;
array[46629] <= 16'b0000_0000_0000_0000;
array[46630] <= 16'b0000_0000_0000_0000;
array[46631] <= 16'b0000_0000_0000_0000;
array[46632] <= 16'b0000_0000_0000_0000;
array[46633] <= 16'b0000_0000_0000_0000;
array[46634] <= 16'b0000_0000_0000_0000;
array[46635] <= 16'b0000_0000_0000_0000;
array[46636] <= 16'b0000_0000_0000_0000;
array[46637] <= 16'b0000_0000_0000_0000;
array[46638] <= 16'b0000_0000_0000_0000;
array[46639] <= 16'b0000_0000_0000_0000;
array[46640] <= 16'b0000_0000_0000_0000;
array[46641] <= 16'b0000_0000_0000_0000;
array[46642] <= 16'b0000_0000_0000_0000;
array[46643] <= 16'b0000_0000_0000_0000;
array[46644] <= 16'b0000_0000_0000_0000;
array[46645] <= 16'b0000_0000_0000_0000;
array[46646] <= 16'b0000_0000_0000_0000;
array[46647] <= 16'b0000_0000_0000_0000;
array[46648] <= 16'b0000_0000_0000_0000;
array[46649] <= 16'b0000_0000_0000_0000;
array[46650] <= 16'b0000_0000_0000_0000;
array[46651] <= 16'b0000_0000_0000_0000;
array[46652] <= 16'b0000_0000_0000_0000;
array[46653] <= 16'b0000_0000_0000_0000;
array[46654] <= 16'b0000_0000_0000_0000;
array[46655] <= 16'b0000_0000_0000_0000;
array[46656] <= 16'b0000_0000_0000_0000;
array[46657] <= 16'b0000_0000_0000_0000;
array[46658] <= 16'b0000_0000_0000_0000;
array[46659] <= 16'b0000_0000_0000_0000;
array[46660] <= 16'b0000_0000_0000_0000;
array[46661] <= 16'b0000_0000_0000_0000;
array[46662] <= 16'b0000_0000_0000_0000;
array[46663] <= 16'b0000_0000_0000_0000;
array[46664] <= 16'b0000_0000_0000_0000;
array[46665] <= 16'b0000_0000_0000_0000;
array[46666] <= 16'b0000_0000_0000_0000;
array[46667] <= 16'b0000_0000_0000_0000;
array[46668] <= 16'b0000_0000_0000_0000;
array[46669] <= 16'b0000_0000_0000_0000;
array[46670] <= 16'b0000_0000_0000_0000;
array[46671] <= 16'b0000_0000_0000_0000;
array[46672] <= 16'b0000_0000_0000_0000;
array[46673] <= 16'b0000_0000_0000_0000;
array[46674] <= 16'b0000_0000_0000_0000;
array[46675] <= 16'b0000_0000_0000_0000;
array[46676] <= 16'b0000_0000_0000_0000;
array[46677] <= 16'b0000_0000_0000_0000;
array[46678] <= 16'b0000_0000_0000_0000;
array[46679] <= 16'b0000_0000_0000_0000;
array[46680] <= 16'b0000_0000_0000_0000;
array[46681] <= 16'b0000_0000_0000_0000;
array[46682] <= 16'b0000_0000_0000_0000;
array[46683] <= 16'b0000_0000_0000_0000;
array[46684] <= 16'b0000_0000_0000_0000;
array[46685] <= 16'b0000_0000_0000_0000;
array[46686] <= 16'b0000_0000_0000_0000;
array[46687] <= 16'b0000_0000_0000_0000;
array[46688] <= 16'b0000_0000_0000_0000;
array[46689] <= 16'b0000_0000_0000_0000;
array[46690] <= 16'b0000_0000_0000_0000;
array[46691] <= 16'b0000_0000_0000_0000;
array[46692] <= 16'b0000_0000_0000_0000;
array[46693] <= 16'b0000_0000_0000_0000;
array[46694] <= 16'b0000_0000_0000_0000;
array[46695] <= 16'b0000_0000_0000_0000;
array[46696] <= 16'b0000_0000_0000_0000;
array[46697] <= 16'b0000_0000_0000_0000;
array[46698] <= 16'b0000_0000_0000_0000;
array[46699] <= 16'b0000_0000_0000_0000;
array[46700] <= 16'b0000_0000_0000_0000;
array[46701] <= 16'b0000_0000_0000_0000;
array[46702] <= 16'b0000_0000_0000_0000;
array[46703] <= 16'b0000_0000_0000_0000;
array[46704] <= 16'b0000_0000_0000_0000;
array[46705] <= 16'b0000_0000_0000_0000;
array[46706] <= 16'b0000_0000_0000_0000;
array[46707] <= 16'b0000_0000_0000_0000;
array[46708] <= 16'b0000_0000_0000_0000;
array[46709] <= 16'b0000_0000_0000_0000;
array[46710] <= 16'b0000_0000_0000_0000;
array[46711] <= 16'b0000_0000_0000_0000;
array[46712] <= 16'b0000_0000_0000_0000;
array[46713] <= 16'b0000_0000_0000_0000;
array[46714] <= 16'b0000_0000_0000_0000;
array[46715] <= 16'b0000_0000_0000_0000;
array[46716] <= 16'b0000_0000_0000_0000;
array[46717] <= 16'b0000_0000_0000_0000;
array[46718] <= 16'b0000_0000_0000_0000;
array[46719] <= 16'b0000_0000_0000_0000;
array[46720] <= 16'b0000_0000_0000_0000;
array[46721] <= 16'b0000_0000_0000_0000;
array[46722] <= 16'b0000_0000_0000_0000;
array[46723] <= 16'b0000_0000_0000_0000;
array[46724] <= 16'b0000_0000_0000_0000;
array[46725] <= 16'b0000_0000_0000_0000;
array[46726] <= 16'b0000_0000_0000_0000;
array[46727] <= 16'b0000_0000_0000_0000;
array[46728] <= 16'b0000_0000_0000_0000;
array[46729] <= 16'b0000_0000_0000_0000;
array[46730] <= 16'b0000_0000_0000_0000;
array[46731] <= 16'b0000_0000_0000_0000;
array[46732] <= 16'b0000_0000_0000_0000;
array[46733] <= 16'b0000_0000_0000_0000;
array[46734] <= 16'b0000_0000_0000_0000;
array[46735] <= 16'b0000_0000_0000_0000;
array[46736] <= 16'b0000_0000_0000_0000;
array[46737] <= 16'b0000_0000_0000_0000;
array[46738] <= 16'b0000_0000_0000_0000;
array[46739] <= 16'b0000_0000_0000_0000;
array[46740] <= 16'b0000_0000_0000_0000;
array[46741] <= 16'b0000_0000_0000_0000;
array[46742] <= 16'b0000_0000_0000_0000;
array[46743] <= 16'b0000_0000_0000_0000;
array[46744] <= 16'b0000_0000_0000_0000;
array[46745] <= 16'b0000_0000_0000_0000;
array[46746] <= 16'b0000_0000_0000_0000;
array[46747] <= 16'b0000_0000_0000_0000;
array[46748] <= 16'b0000_0000_0000_0000;
array[46749] <= 16'b0000_0000_0000_0000;
array[46750] <= 16'b0000_0000_0000_0000;
array[46751] <= 16'b0000_0000_0000_0000;
array[46752] <= 16'b0000_0000_0000_0000;
array[46753] <= 16'b0000_0000_0000_0000;
array[46754] <= 16'b0000_0000_0000_0000;
array[46755] <= 16'b0000_0000_0000_0000;
array[46756] <= 16'b0000_0000_0000_0000;
array[46757] <= 16'b0000_0000_0000_0000;
array[46758] <= 16'b0000_0000_0000_0000;
array[46759] <= 16'b0000_0000_0000_0000;
array[46760] <= 16'b0000_0000_0000_0000;
array[46761] <= 16'b0000_0000_0000_0000;
array[46762] <= 16'b0000_0000_0000_0000;
array[46763] <= 16'b0000_0000_0000_0000;
array[46764] <= 16'b0000_0000_0000_0000;
array[46765] <= 16'b0000_0000_0000_0000;
array[46766] <= 16'b0000_0000_0000_0000;
array[46767] <= 16'b0000_0000_0000_0000;
array[46768] <= 16'b0000_0000_0000_0000;
array[46769] <= 16'b0000_0000_0000_0000;
array[46770] <= 16'b0000_0000_0000_0000;
array[46771] <= 16'b0000_0000_0000_0000;
array[46772] <= 16'b0000_0000_0000_0000;
array[46773] <= 16'b0000_0000_0000_0000;
array[46774] <= 16'b0000_0000_0000_0000;
array[46775] <= 16'b0000_0000_0000_0000;
array[46776] <= 16'b0000_0000_0000_0000;
array[46777] <= 16'b0000_0000_0000_0000;
array[46778] <= 16'b0000_0000_0000_0000;
array[46779] <= 16'b0000_0000_0000_0000;
array[46780] <= 16'b0000_0000_0000_0000;
array[46781] <= 16'b0000_0000_0000_0000;
array[46782] <= 16'b0000_0000_0000_0000;
array[46783] <= 16'b0000_0000_0000_0000;
array[46784] <= 16'b0000_0000_0000_0000;
array[46785] <= 16'b0000_0000_0000_0000;
array[46786] <= 16'b0000_0000_0000_0000;
array[46787] <= 16'b0000_0000_0000_0000;
array[46788] <= 16'b0000_0000_0000_0000;
array[46789] <= 16'b0000_0000_0000_0000;
array[46790] <= 16'b0000_0000_0000_0000;
array[46791] <= 16'b0000_0000_0000_0000;
array[46792] <= 16'b0000_0000_0000_0000;
array[46793] <= 16'b0000_0000_0000_0000;
array[46794] <= 16'b0000_0000_0000_0000;
array[46795] <= 16'b0000_0000_0000_0000;
array[46796] <= 16'b0000_0000_0000_0000;
array[46797] <= 16'b0000_0000_0000_0000;
array[46798] <= 16'b0000_0000_0000_0000;
array[46799] <= 16'b0000_0000_0000_0000;
array[46800] <= 16'b0000_0000_0000_0000;
array[46801] <= 16'b0000_0000_0000_0000;
array[46802] <= 16'b0000_0000_0000_0000;
array[46803] <= 16'b0000_0000_0000_0000;
array[46804] <= 16'b0000_0000_0000_0000;
array[46805] <= 16'b0000_0000_0000_0000;
array[46806] <= 16'b0000_0000_0000_0000;
array[46807] <= 16'b0000_0000_0000_0000;
array[46808] <= 16'b0000_0000_0000_0000;
array[46809] <= 16'b0000_0000_0000_0000;
array[46810] <= 16'b0000_0000_0000_0000;
array[46811] <= 16'b0000_0000_0000_0000;
array[46812] <= 16'b0000_0000_0000_0000;
array[46813] <= 16'b0000_0000_0000_0000;
array[46814] <= 16'b0000_0000_0000_0000;
array[46815] <= 16'b0000_0000_0000_0000;
array[46816] <= 16'b0000_0000_0000_0000;
array[46817] <= 16'b0000_0000_0000_0000;
array[46818] <= 16'b0000_0000_0000_0000;
array[46819] <= 16'b0000_0000_0000_0000;
array[46820] <= 16'b0000_0000_0000_0000;
array[46821] <= 16'b0000_0000_0000_0000;
array[46822] <= 16'b0000_0000_0000_0000;
array[46823] <= 16'b0000_0000_0000_0000;
array[46824] <= 16'b0000_0000_0000_0000;
array[46825] <= 16'b0000_0000_0000_0000;
array[46826] <= 16'b0000_0000_0000_0000;
array[46827] <= 16'b0000_0000_0000_0000;
array[46828] <= 16'b0000_0000_0000_0000;
array[46829] <= 16'b0000_0000_0000_0000;
array[46830] <= 16'b0000_0000_0000_0000;
array[46831] <= 16'b0000_0000_0000_0000;
array[46832] <= 16'b0000_0000_0000_0000;
array[46833] <= 16'b0000_0000_0000_0000;
array[46834] <= 16'b0000_0000_0000_0000;
array[46835] <= 16'b0000_0000_0000_0000;
array[46836] <= 16'b0000_0000_0000_0000;
array[46837] <= 16'b0000_0000_0000_0000;
array[46838] <= 16'b0000_0000_0000_0000;
array[46839] <= 16'b0000_0000_0000_0000;
array[46840] <= 16'b0000_0000_0000_0000;
array[46841] <= 16'b0000_0000_0000_0000;
array[46842] <= 16'b0000_0000_0000_0000;
array[46843] <= 16'b0000_0000_0000_0000;
array[46844] <= 16'b0000_0000_0000_0000;
array[46845] <= 16'b0000_0000_0000_0000;
array[46846] <= 16'b0000_0000_0000_0000;
array[46847] <= 16'b0000_0000_0000_0000;
array[46848] <= 16'b0000_0000_0000_0000;
array[46849] <= 16'b0000_0000_0000_0000;
array[46850] <= 16'b0000_0000_0000_0000;
array[46851] <= 16'b0000_0000_0000_0000;
array[46852] <= 16'b0000_0000_0000_0000;
array[46853] <= 16'b0000_0000_0000_0000;
array[46854] <= 16'b0000_0000_0000_0000;
array[46855] <= 16'b0000_0000_0000_0000;
array[46856] <= 16'b0000_0000_0000_0000;
array[46857] <= 16'b0000_0000_0000_0000;
array[46858] <= 16'b0000_0000_0000_0000;
array[46859] <= 16'b0000_0000_0000_0000;
array[46860] <= 16'b0000_0000_0000_0000;
array[46861] <= 16'b0000_0000_0000_0000;
array[46862] <= 16'b0000_0000_0000_0000;
array[46863] <= 16'b0000_0000_0000_0000;
array[46864] <= 16'b0000_0000_0000_0000;
array[46865] <= 16'b0000_0000_0000_0000;
array[46866] <= 16'b0000_0000_0000_0000;
array[46867] <= 16'b0000_0000_0000_0000;
array[46868] <= 16'b0000_0000_0000_0000;
array[46869] <= 16'b0000_0000_0000_0000;
array[46870] <= 16'b0000_0000_0000_0000;
array[46871] <= 16'b0000_0000_0000_0000;
array[46872] <= 16'b0000_0000_0000_0000;
array[46873] <= 16'b0000_0000_0000_0000;
array[46874] <= 16'b0000_0000_0000_0000;
array[46875] <= 16'b0000_0000_0000_0000;
array[46876] <= 16'b0000_0000_0000_0000;
array[46877] <= 16'b0000_0000_0000_0000;
array[46878] <= 16'b0000_0000_0000_0000;
array[46879] <= 16'b0000_0000_0000_0000;
array[46880] <= 16'b0000_0000_0000_0000;
array[46881] <= 16'b0000_0000_0000_0000;
array[46882] <= 16'b0000_0000_0000_0000;
array[46883] <= 16'b0000_0000_0000_0000;
array[46884] <= 16'b0000_0000_0000_0000;
array[46885] <= 16'b0000_0000_0000_0000;
array[46886] <= 16'b0000_0000_0000_0000;
array[46887] <= 16'b0000_0000_0000_0000;
array[46888] <= 16'b0000_0000_0000_0000;
array[46889] <= 16'b0000_0000_0000_0000;
array[46890] <= 16'b0000_0000_0000_0000;
array[46891] <= 16'b0000_0000_0000_0000;
array[46892] <= 16'b0000_0000_0000_0000;
array[46893] <= 16'b0000_0000_0000_0000;
array[46894] <= 16'b0000_0000_0000_0000;
array[46895] <= 16'b0000_0000_0000_0000;
array[46896] <= 16'b0000_0000_0000_0000;
array[46897] <= 16'b0000_0000_0000_0000;
array[46898] <= 16'b0000_0000_0000_0000;
array[46899] <= 16'b0000_0000_0000_0000;
array[46900] <= 16'b0000_0000_0000_0000;
array[46901] <= 16'b0000_0000_0000_0000;
array[46902] <= 16'b0000_0000_0000_0000;
array[46903] <= 16'b0000_0000_0000_0000;
array[46904] <= 16'b0000_0000_0000_0000;
array[46905] <= 16'b0000_0000_0000_0000;
array[46906] <= 16'b0000_0000_0000_0000;
array[46907] <= 16'b0000_0000_0000_0000;
array[46908] <= 16'b0000_0000_0000_0000;
array[46909] <= 16'b0000_0000_0000_0000;
array[46910] <= 16'b0000_0000_0000_0000;
array[46911] <= 16'b0000_0000_0000_0000;
array[46912] <= 16'b0000_0000_0000_0000;
array[46913] <= 16'b0000_0000_0000_0000;
array[46914] <= 16'b0000_0000_0000_0000;
array[46915] <= 16'b0000_0000_0000_0000;
array[46916] <= 16'b0000_0000_0000_0000;
array[46917] <= 16'b0000_0000_0000_0000;
array[46918] <= 16'b0000_0000_0000_0000;
array[46919] <= 16'b0000_0000_0000_0000;
array[46920] <= 16'b0000_0000_0000_0000;
array[46921] <= 16'b0000_0000_0000_0000;
array[46922] <= 16'b0000_0000_0000_0000;
array[46923] <= 16'b0000_0000_0000_0000;
array[46924] <= 16'b0000_0000_0000_0000;
array[46925] <= 16'b0000_0000_0000_0000;
array[46926] <= 16'b0000_0000_0000_0000;
array[46927] <= 16'b0000_0000_0000_0000;
array[46928] <= 16'b0000_0000_0000_0000;
array[46929] <= 16'b0000_0000_0000_0000;
array[46930] <= 16'b0000_0000_0000_0000;
array[46931] <= 16'b0000_0000_0000_0000;
array[46932] <= 16'b0000_0000_0000_0000;
array[46933] <= 16'b0000_0000_0000_0000;
array[46934] <= 16'b0000_0000_0000_0000;
array[46935] <= 16'b0000_0000_0000_0000;
array[46936] <= 16'b0000_0000_0000_0000;
array[46937] <= 16'b0000_0000_0000_0000;
array[46938] <= 16'b0000_0000_0000_0000;
array[46939] <= 16'b0000_0000_0000_0000;
array[46940] <= 16'b0000_0000_0000_0000;
array[46941] <= 16'b0000_0000_0000_0000;
array[46942] <= 16'b0000_0000_0000_0000;
array[46943] <= 16'b0000_0000_0000_0000;
array[46944] <= 16'b0000_0000_0000_0000;
array[46945] <= 16'b0000_0000_0000_0000;
array[46946] <= 16'b0000_0000_0000_0000;
array[46947] <= 16'b0000_0000_0000_0000;
array[46948] <= 16'b0000_0000_0000_0000;
array[46949] <= 16'b0000_0000_0000_0000;
array[46950] <= 16'b0000_0000_0000_0000;
array[46951] <= 16'b0000_0000_0000_0000;
array[46952] <= 16'b0000_0000_0000_0000;
array[46953] <= 16'b0000_0000_0000_0000;
array[46954] <= 16'b0000_0000_0000_0000;
array[46955] <= 16'b0000_0000_0000_0000;
array[46956] <= 16'b0000_0000_0000_0000;
array[46957] <= 16'b0000_0000_0000_0000;
array[46958] <= 16'b0000_0000_0000_0000;
array[46959] <= 16'b0000_0000_0000_0000;
array[46960] <= 16'b0000_0000_0000_0000;
array[46961] <= 16'b0000_0000_0000_0000;
array[46962] <= 16'b0000_0000_0000_0000;
array[46963] <= 16'b0000_0000_0000_0000;
array[46964] <= 16'b0000_0000_0000_0000;
array[46965] <= 16'b0000_0000_0000_0000;
array[46966] <= 16'b0000_0000_0000_0000;
array[46967] <= 16'b0000_0000_0000_0000;
array[46968] <= 16'b0000_0000_0000_0000;
array[46969] <= 16'b0000_0000_0000_0000;
array[46970] <= 16'b0000_0000_0000_0000;
array[46971] <= 16'b0000_0000_0000_0000;
array[46972] <= 16'b0000_0000_0000_0000;
array[46973] <= 16'b0000_0000_0000_0000;
array[46974] <= 16'b0000_0000_0000_0000;
array[46975] <= 16'b0000_0000_0000_0000;
array[46976] <= 16'b0000_0000_0000_0000;
array[46977] <= 16'b0000_0000_0000_0000;
array[46978] <= 16'b0000_0000_0000_0000;
array[46979] <= 16'b0000_0000_0000_0000;
array[46980] <= 16'b0000_0000_0000_0000;
array[46981] <= 16'b0000_0000_0000_0000;
array[46982] <= 16'b0000_0000_0000_0000;
array[46983] <= 16'b0000_0000_0000_0000;
array[46984] <= 16'b0000_0000_0000_0000;
array[46985] <= 16'b0000_0000_0000_0000;
array[46986] <= 16'b0000_0000_0000_0000;
array[46987] <= 16'b0000_0000_0000_0000;
array[46988] <= 16'b0000_0000_0000_0000;
array[46989] <= 16'b0000_0000_0000_0000;
array[46990] <= 16'b0000_0000_0000_0000;
array[46991] <= 16'b0000_0000_0000_0000;
array[46992] <= 16'b0000_0000_0000_0000;
array[46993] <= 16'b0000_0000_0000_0000;
array[46994] <= 16'b0000_0000_0000_0000;
array[46995] <= 16'b0000_0000_0000_0000;
array[46996] <= 16'b0000_0000_0000_0000;
array[46997] <= 16'b0000_0000_0000_0000;
array[46998] <= 16'b0000_0000_0000_0000;
array[46999] <= 16'b0000_0000_0000_0000;
array[47000] <= 16'b0000_0000_0000_0000;
array[47001] <= 16'b0000_0000_0000_0000;
array[47002] <= 16'b0000_0000_0000_0000;
array[47003] <= 16'b0000_0000_0000_0000;
array[47004] <= 16'b0000_0000_0000_0000;
array[47005] <= 16'b0000_0000_0000_0000;
array[47006] <= 16'b0000_0000_0000_0000;
array[47007] <= 16'b0000_0000_0000_0000;
array[47008] <= 16'b0000_0000_0000_0000;
array[47009] <= 16'b0000_0000_0000_0000;
array[47010] <= 16'b0000_0000_0000_0000;
array[47011] <= 16'b0000_0000_0000_0000;
array[47012] <= 16'b0000_0000_0000_0000;
array[47013] <= 16'b0000_0000_0000_0000;
array[47014] <= 16'b0000_0000_0000_0000;
array[47015] <= 16'b0000_0000_0000_0000;
array[47016] <= 16'b0000_0000_0000_0000;
array[47017] <= 16'b0000_0000_0000_0000;
array[47018] <= 16'b0000_0000_0000_0000;
array[47019] <= 16'b0000_0000_0000_0000;
array[47020] <= 16'b0000_0000_0000_0000;
array[47021] <= 16'b0000_0000_0000_0000;
array[47022] <= 16'b0000_0000_0000_0000;
array[47023] <= 16'b0000_0000_0000_0000;
array[47024] <= 16'b0000_0000_0000_0000;
array[47025] <= 16'b0000_0000_0000_0000;
array[47026] <= 16'b0000_0000_0000_0000;
array[47027] <= 16'b0000_0000_0000_0000;
array[47028] <= 16'b0000_0000_0000_0000;
array[47029] <= 16'b0000_0000_0000_0000;
array[47030] <= 16'b0000_0000_0000_0000;
array[47031] <= 16'b0000_0000_0000_0000;
array[47032] <= 16'b0000_0000_0000_0000;
array[47033] <= 16'b0000_0000_0000_0000;
array[47034] <= 16'b0000_0000_0000_0000;
array[47035] <= 16'b0000_0000_0000_0000;
array[47036] <= 16'b0000_0000_0000_0000;
array[47037] <= 16'b0000_0000_0000_0000;
array[47038] <= 16'b0000_0000_0000_0000;
array[47039] <= 16'b0000_0000_0000_0000;
array[47040] <= 16'b0000_0000_0000_0000;
array[47041] <= 16'b0000_0000_0000_0000;
array[47042] <= 16'b0000_0000_0000_0000;
array[47043] <= 16'b0000_0000_0000_0000;
array[47044] <= 16'b0000_0000_0000_0000;
array[47045] <= 16'b0000_0000_0000_0000;
array[47046] <= 16'b0000_0000_0000_0000;
array[47047] <= 16'b0000_0000_0000_0000;
array[47048] <= 16'b0000_0000_0000_0000;
array[47049] <= 16'b0000_0000_0000_0000;
array[47050] <= 16'b0000_0000_0000_0000;
array[47051] <= 16'b0000_0000_0000_0000;
array[47052] <= 16'b0000_0000_0000_0000;
array[47053] <= 16'b0000_0000_0000_0000;
array[47054] <= 16'b0000_0000_0000_0000;
array[47055] <= 16'b0000_0000_0000_0000;
array[47056] <= 16'b0000_0000_0000_0000;
array[47057] <= 16'b0000_0000_0000_0000;
array[47058] <= 16'b0000_0000_0000_0000;
array[47059] <= 16'b0000_0000_0000_0000;
array[47060] <= 16'b0000_0000_0000_0000;
array[47061] <= 16'b0000_0000_0000_0000;
array[47062] <= 16'b0000_0000_0000_0000;
array[47063] <= 16'b0000_0000_0000_0000;
array[47064] <= 16'b0000_0000_0000_0000;
array[47065] <= 16'b0000_0000_0000_0000;
array[47066] <= 16'b0000_0000_0000_0000;
array[47067] <= 16'b0000_0000_0000_0000;
array[47068] <= 16'b0000_0000_0000_0000;
array[47069] <= 16'b0000_0000_0000_0000;
array[47070] <= 16'b0000_0000_0000_0000;
array[47071] <= 16'b0000_0000_0000_0000;
array[47072] <= 16'b0000_0000_0000_0000;
array[47073] <= 16'b0000_0000_0000_0000;
array[47074] <= 16'b0000_0000_0000_0000;
array[47075] <= 16'b0000_0000_0000_0000;
array[47076] <= 16'b0000_0000_0000_0000;
array[47077] <= 16'b0000_0000_0000_0000;
array[47078] <= 16'b0000_0000_0000_0000;
array[47079] <= 16'b0000_0000_0000_0000;
array[47080] <= 16'b0000_0000_0000_0000;
array[47081] <= 16'b0000_0000_0000_0000;
array[47082] <= 16'b0000_0000_0000_0000;
array[47083] <= 16'b0000_0000_0000_0000;
array[47084] <= 16'b0000_0000_0000_0000;
array[47085] <= 16'b0000_0000_0000_0000;
array[47086] <= 16'b0000_0000_0000_0000;
array[47087] <= 16'b0000_0000_0000_0000;
array[47088] <= 16'b0000_0000_0000_0000;
array[47089] <= 16'b0000_0000_0000_0000;
array[47090] <= 16'b0000_0000_0000_0000;
array[47091] <= 16'b0000_0000_0000_0000;
array[47092] <= 16'b0000_0000_0000_0000;
array[47093] <= 16'b0000_0000_0000_0000;
array[47094] <= 16'b0000_0000_0000_0000;
array[47095] <= 16'b0000_0000_0000_0000;
array[47096] <= 16'b0000_0000_0000_0000;
array[47097] <= 16'b0000_0000_0000_0000;
array[47098] <= 16'b0000_0000_0000_0000;
array[47099] <= 16'b0000_0000_0000_0000;
array[47100] <= 16'b0000_0000_0000_0000;
array[47101] <= 16'b0000_0000_0000_0000;
array[47102] <= 16'b0000_0000_0000_0000;
array[47103] <= 16'b0000_0000_0000_0000;
array[47104] <= 16'b0000_0000_0000_0000;
array[47105] <= 16'b0000_0000_0000_0000;
array[47106] <= 16'b0000_0000_0000_0000;
array[47107] <= 16'b0000_0000_0000_0000;
array[47108] <= 16'b0000_0000_0000_0000;
array[47109] <= 16'b0000_0000_0000_0000;
array[47110] <= 16'b0000_0000_0000_0000;
array[47111] <= 16'b0000_0000_0000_0000;
array[47112] <= 16'b0000_0000_0000_0000;
array[47113] <= 16'b0000_0000_0000_0000;
array[47114] <= 16'b0000_0000_0000_0000;
array[47115] <= 16'b0000_0000_0000_0000;
array[47116] <= 16'b0000_0000_0000_0000;
array[47117] <= 16'b0000_0000_0000_0000;
array[47118] <= 16'b0000_0000_0000_0000;
array[47119] <= 16'b0000_0000_0000_0000;
array[47120] <= 16'b0000_0000_0000_0000;
array[47121] <= 16'b0000_0000_0000_0000;
array[47122] <= 16'b0000_0000_0000_0000;
array[47123] <= 16'b0000_0000_0000_0000;
array[47124] <= 16'b0000_0000_0000_0000;
array[47125] <= 16'b0000_0000_0000_0000;
array[47126] <= 16'b0000_0000_0000_0000;
array[47127] <= 16'b0000_0000_0000_0000;
array[47128] <= 16'b0000_0000_0000_0000;
array[47129] <= 16'b0000_0000_0000_0000;
array[47130] <= 16'b0000_0000_0000_0000;
array[47131] <= 16'b0000_0000_0000_0000;
array[47132] <= 16'b0000_0000_0000_0000;
array[47133] <= 16'b0000_0000_0000_0000;
array[47134] <= 16'b0000_0000_0000_0000;
array[47135] <= 16'b0000_0000_0000_0000;
array[47136] <= 16'b0000_0000_0000_0000;
array[47137] <= 16'b0000_0000_0000_0000;
array[47138] <= 16'b0000_0000_0000_0000;
array[47139] <= 16'b0000_0000_0000_0000;
array[47140] <= 16'b0000_0000_0000_0000;
array[47141] <= 16'b0000_0000_0000_0000;
array[47142] <= 16'b0000_0000_0000_0000;
array[47143] <= 16'b0000_0000_0000_0000;
array[47144] <= 16'b0000_0000_0000_0000;
array[47145] <= 16'b0000_0000_0000_0000;
array[47146] <= 16'b0000_0000_0000_0000;
array[47147] <= 16'b0000_0000_0000_0000;
array[47148] <= 16'b0000_0000_0000_0000;
array[47149] <= 16'b0000_0000_0000_0000;
array[47150] <= 16'b0000_0000_0000_0000;
array[47151] <= 16'b0000_0000_0000_0000;
array[47152] <= 16'b0000_0000_0000_0000;
array[47153] <= 16'b0000_0000_0000_0000;
array[47154] <= 16'b0000_0000_0000_0000;
array[47155] <= 16'b0000_0000_0000_0000;
array[47156] <= 16'b0000_0000_0000_0000;
array[47157] <= 16'b0000_0000_0000_0000;
array[47158] <= 16'b0000_0000_0000_0000;
array[47159] <= 16'b0000_0000_0000_0000;
array[47160] <= 16'b0000_0000_0000_0000;
array[47161] <= 16'b0000_0000_0000_0000;
array[47162] <= 16'b0000_0000_0000_0000;
array[47163] <= 16'b0000_0000_0000_0000;
array[47164] <= 16'b0000_0000_0000_0000;
array[47165] <= 16'b0000_0000_0000_0000;
array[47166] <= 16'b0000_0000_0000_0000;
array[47167] <= 16'b0000_0000_0000_0000;
array[47168] <= 16'b0000_0000_0000_0000;
array[47169] <= 16'b0000_0000_0000_0000;
array[47170] <= 16'b0000_0000_0000_0000;
array[47171] <= 16'b0000_0000_0000_0000;
array[47172] <= 16'b0000_0000_0000_0000;
array[47173] <= 16'b0000_0000_0000_0000;
array[47174] <= 16'b0000_0000_0000_0000;
array[47175] <= 16'b0000_0000_0000_0000;
array[47176] <= 16'b0000_0000_0000_0000;
array[47177] <= 16'b0000_0000_0000_0000;
array[47178] <= 16'b0000_0000_0000_0000;
array[47179] <= 16'b0000_0000_0000_0000;
array[47180] <= 16'b0000_0000_0000_0000;
array[47181] <= 16'b0000_0000_0000_0000;
array[47182] <= 16'b0000_0000_0000_0000;
array[47183] <= 16'b0000_0000_0000_0000;
array[47184] <= 16'b0000_0000_0000_0000;
array[47185] <= 16'b0000_0000_0000_0000;
array[47186] <= 16'b0000_0000_0000_0000;
array[47187] <= 16'b0000_0000_0000_0000;
array[47188] <= 16'b0000_0000_0000_0000;
array[47189] <= 16'b0000_0000_0000_0000;
array[47190] <= 16'b0000_0000_0000_0000;
array[47191] <= 16'b0000_0000_0000_0000;
array[47192] <= 16'b0000_0000_0000_0000;
array[47193] <= 16'b0000_0000_0000_0000;
array[47194] <= 16'b0000_0000_0000_0000;
array[47195] <= 16'b0000_0000_0000_0000;
array[47196] <= 16'b0000_0000_0000_0000;
array[47197] <= 16'b0000_0000_0000_0000;
array[47198] <= 16'b0000_0000_0000_0000;
array[47199] <= 16'b0000_0000_0000_0000;
array[47200] <= 16'b0000_0000_0000_0000;
array[47201] <= 16'b0000_0000_0000_0000;
array[47202] <= 16'b0000_0000_0000_0000;
array[47203] <= 16'b0000_0000_0000_0000;
array[47204] <= 16'b0000_0000_0000_0000;
array[47205] <= 16'b0000_0000_0000_0000;
array[47206] <= 16'b0000_0000_0000_0000;
array[47207] <= 16'b0000_0000_0000_0000;
array[47208] <= 16'b0000_0000_0000_0000;
array[47209] <= 16'b0000_0000_0000_0000;
array[47210] <= 16'b0000_0000_0000_0000;
array[47211] <= 16'b0000_0000_0000_0000;
array[47212] <= 16'b0000_0000_0000_0000;
array[47213] <= 16'b0000_0000_0000_0000;
array[47214] <= 16'b0000_0000_0000_0000;
array[47215] <= 16'b0000_0000_0000_0000;
array[47216] <= 16'b0000_0000_0000_0000;
array[47217] <= 16'b0000_0000_0000_0000;
array[47218] <= 16'b0000_0000_0000_0000;
array[47219] <= 16'b0000_0000_0000_0000;
array[47220] <= 16'b0000_0000_0000_0000;
array[47221] <= 16'b0000_0000_0000_0000;
array[47222] <= 16'b0000_0000_0000_0000;
array[47223] <= 16'b0000_0000_0000_0000;
array[47224] <= 16'b0000_0000_0000_0000;
array[47225] <= 16'b0000_0000_0000_0000;
array[47226] <= 16'b0000_0000_0000_0000;
array[47227] <= 16'b0000_0000_0000_0000;
array[47228] <= 16'b0000_0000_0000_0000;
array[47229] <= 16'b0000_0000_0000_0000;
array[47230] <= 16'b0000_0000_0000_0000;
array[47231] <= 16'b0000_0000_0000_0000;
array[47232] <= 16'b0000_0000_0000_0000;
array[47233] <= 16'b0000_0000_0000_0000;
array[47234] <= 16'b0000_0000_0000_0000;
array[47235] <= 16'b0000_0000_0000_0000;
array[47236] <= 16'b0000_0000_0000_0000;
array[47237] <= 16'b0000_0000_0000_0000;
array[47238] <= 16'b0000_0000_0000_0000;
array[47239] <= 16'b0000_0000_0000_0000;
array[47240] <= 16'b0000_0000_0000_0000;
array[47241] <= 16'b0000_0000_0000_0000;
array[47242] <= 16'b0000_0000_0000_0000;
array[47243] <= 16'b0000_0000_0000_0000;
array[47244] <= 16'b0000_0000_0000_0000;
array[47245] <= 16'b0000_0000_0000_0000;
array[47246] <= 16'b0000_0000_0000_0000;
array[47247] <= 16'b0000_0000_0000_0000;
array[47248] <= 16'b0000_0000_0000_0000;
array[47249] <= 16'b0000_0000_0000_0000;
array[47250] <= 16'b0000_0000_0000_0000;
array[47251] <= 16'b0000_0000_0000_0000;
array[47252] <= 16'b0000_0000_0000_0000;
array[47253] <= 16'b0000_0000_0000_0000;
array[47254] <= 16'b0000_0000_0000_0000;
array[47255] <= 16'b0000_0000_0000_0000;
array[47256] <= 16'b0000_0000_0000_0000;
array[47257] <= 16'b0000_0000_0000_0000;
array[47258] <= 16'b0000_0000_0000_0000;
array[47259] <= 16'b0000_0000_0000_0000;
array[47260] <= 16'b0000_0000_0000_0000;
array[47261] <= 16'b0000_0000_0000_0000;
array[47262] <= 16'b0000_0000_0000_0000;
array[47263] <= 16'b0000_0000_0000_0000;
array[47264] <= 16'b0000_0000_0000_0000;
array[47265] <= 16'b0000_0000_0000_0000;
array[47266] <= 16'b0000_0000_0000_0000;
array[47267] <= 16'b0000_0000_0000_0000;
array[47268] <= 16'b0000_0000_0000_0000;
array[47269] <= 16'b0000_0000_0000_0000;
array[47270] <= 16'b0000_0000_0000_0000;
array[47271] <= 16'b0000_0000_0000_0000;
array[47272] <= 16'b0000_0000_0000_0000;
array[47273] <= 16'b0000_0000_0000_0000;
array[47274] <= 16'b0000_0000_0000_0000;
array[47275] <= 16'b0000_0000_0000_0000;
array[47276] <= 16'b0000_0000_0000_0000;
array[47277] <= 16'b0000_0000_0000_0000;
array[47278] <= 16'b0000_0000_0000_0000;
array[47279] <= 16'b0000_0000_0000_0000;
array[47280] <= 16'b0000_0000_0000_0000;
array[47281] <= 16'b0000_0000_0000_0000;
array[47282] <= 16'b0000_0000_0000_0000;
array[47283] <= 16'b0000_0000_0000_0000;
array[47284] <= 16'b0000_0000_0000_0000;
array[47285] <= 16'b0000_0000_0000_0000;
array[47286] <= 16'b0000_0000_0000_0000;
array[47287] <= 16'b0000_0000_0000_0000;
array[47288] <= 16'b0000_0000_0000_0000;
array[47289] <= 16'b0000_0000_0000_0000;
array[47290] <= 16'b0000_0000_0000_0000;
array[47291] <= 16'b0000_0000_0000_0000;
array[47292] <= 16'b0000_0000_0000_0000;
array[47293] <= 16'b0000_0000_0000_0000;
array[47294] <= 16'b0000_0000_0000_0000;
array[47295] <= 16'b0000_0000_0000_0000;
array[47296] <= 16'b0000_0000_0000_0000;
array[47297] <= 16'b0000_0000_0000_0000;
array[47298] <= 16'b0000_0000_0000_0000;
array[47299] <= 16'b0000_0000_0000_0000;
array[47300] <= 16'b0000_0000_0000_0000;
array[47301] <= 16'b0000_0000_0000_0000;
array[47302] <= 16'b0000_0000_0000_0000;
array[47303] <= 16'b0000_0000_0000_0000;
array[47304] <= 16'b0000_0000_0000_0000;
array[47305] <= 16'b0000_0000_0000_0000;
array[47306] <= 16'b0000_0000_0000_0000;
array[47307] <= 16'b0000_0000_0000_0000;
array[47308] <= 16'b0000_0000_0000_0000;
array[47309] <= 16'b0000_0000_0000_0000;
array[47310] <= 16'b0000_0000_0000_0000;
array[47311] <= 16'b0000_0000_0000_0000;
array[47312] <= 16'b0000_0000_0000_0000;
array[47313] <= 16'b0000_0000_0000_0000;
array[47314] <= 16'b0000_0000_0000_0000;
array[47315] <= 16'b0000_0000_0000_0000;
array[47316] <= 16'b0000_0000_0000_0000;
array[47317] <= 16'b0000_0000_0000_0000;
array[47318] <= 16'b0000_0000_0000_0000;
array[47319] <= 16'b0000_0000_0000_0000;
array[47320] <= 16'b0000_0000_0000_0000;
array[47321] <= 16'b0000_0000_0000_0000;
array[47322] <= 16'b0000_0000_0000_0000;
array[47323] <= 16'b0000_0000_0000_0000;
array[47324] <= 16'b0000_0000_0000_0000;
array[47325] <= 16'b0000_0000_0000_0000;
array[47326] <= 16'b0000_0000_0000_0000;
array[47327] <= 16'b0000_0000_0000_0000;
array[47328] <= 16'b0000_0000_0000_0000;
array[47329] <= 16'b0000_0000_0000_0000;
array[47330] <= 16'b0000_0000_0000_0000;
array[47331] <= 16'b0000_0000_0000_0000;
array[47332] <= 16'b0000_0000_0000_0000;
array[47333] <= 16'b0000_0000_0000_0000;
array[47334] <= 16'b0000_0000_0000_0000;
array[47335] <= 16'b0000_0000_0000_0000;
array[47336] <= 16'b0000_0000_0000_0000;
array[47337] <= 16'b0000_0000_0000_0000;
array[47338] <= 16'b0000_0000_0000_0000;
array[47339] <= 16'b0000_0000_0000_0000;
array[47340] <= 16'b0000_0000_0000_0000;
array[47341] <= 16'b0000_0000_0000_0000;
array[47342] <= 16'b0000_0000_0000_0000;
array[47343] <= 16'b0000_0000_0000_0000;
array[47344] <= 16'b0000_0000_0000_0000;
array[47345] <= 16'b0000_0000_0000_0000;
array[47346] <= 16'b0000_0000_0000_0000;
array[47347] <= 16'b0000_0000_0000_0000;
array[47348] <= 16'b0000_0000_0000_0000;
array[47349] <= 16'b0000_0000_0000_0000;
array[47350] <= 16'b0000_0000_0000_0000;
array[47351] <= 16'b0000_0000_0000_0000;
array[47352] <= 16'b0000_0000_0000_0000;
array[47353] <= 16'b0000_0000_0000_0000;
array[47354] <= 16'b0000_0000_0000_0000;
array[47355] <= 16'b0000_0000_0000_0000;
array[47356] <= 16'b0000_0000_0000_0000;
array[47357] <= 16'b0000_0000_0000_0000;
array[47358] <= 16'b0000_0000_0000_0000;
array[47359] <= 16'b0000_0000_0000_0000;
array[47360] <= 16'b0000_0000_0000_0000;
array[47361] <= 16'b0000_0000_0000_0000;
array[47362] <= 16'b0000_0000_0000_0000;
array[47363] <= 16'b0000_0000_0000_0000;
array[47364] <= 16'b0000_0000_0000_0000;
array[47365] <= 16'b0000_0000_0000_0000;
array[47366] <= 16'b0000_0000_0000_0000;
array[47367] <= 16'b0000_0000_0000_0000;
array[47368] <= 16'b0000_0000_0000_0000;
array[47369] <= 16'b0000_0000_0000_0000;
array[47370] <= 16'b0000_0000_0000_0000;
array[47371] <= 16'b0000_0000_0000_0000;
array[47372] <= 16'b0000_0000_0000_0000;
array[47373] <= 16'b0000_0000_0000_0000;
array[47374] <= 16'b0000_0000_0000_0000;
array[47375] <= 16'b0000_0000_0000_0000;
array[47376] <= 16'b0000_0000_0000_0000;
array[47377] <= 16'b0000_0000_0000_0000;
array[47378] <= 16'b0000_0000_0000_0000;
array[47379] <= 16'b0000_0000_0000_0000;
array[47380] <= 16'b0000_0000_0000_0000;
array[47381] <= 16'b0000_0000_0000_0000;
array[47382] <= 16'b0000_0000_0000_0000;
array[47383] <= 16'b0000_0000_0000_0000;
array[47384] <= 16'b0000_0000_0000_0000;
array[47385] <= 16'b0000_0000_0000_0000;
array[47386] <= 16'b0000_0000_0000_0000;
array[47387] <= 16'b0000_0000_0000_0000;
array[47388] <= 16'b0000_0000_0000_0000;
array[47389] <= 16'b0000_0000_0000_0000;
array[47390] <= 16'b0000_0000_0000_0000;
array[47391] <= 16'b0000_0000_0000_0000;
array[47392] <= 16'b0000_0000_0000_0000;
array[47393] <= 16'b0000_0000_0000_0000;
array[47394] <= 16'b0000_0000_0000_0000;
array[47395] <= 16'b0000_0000_0000_0000;
array[47396] <= 16'b0000_0000_0000_0000;
array[47397] <= 16'b0000_0000_0000_0000;
array[47398] <= 16'b0000_0000_0000_0000;
array[47399] <= 16'b0000_0000_0000_0000;
array[47400] <= 16'b0000_0000_0000_0000;
array[47401] <= 16'b0000_0000_0000_0000;
array[47402] <= 16'b0000_0000_0000_0000;
array[47403] <= 16'b0000_0000_0000_0000;
array[47404] <= 16'b0000_0000_0000_0000;
array[47405] <= 16'b0000_0000_0000_0000;
array[47406] <= 16'b0000_0000_0000_0000;
array[47407] <= 16'b0000_0000_0000_0000;
array[47408] <= 16'b0000_0000_0000_0000;
array[47409] <= 16'b0000_0000_0000_0000;
array[47410] <= 16'b0000_0000_0000_0000;
array[47411] <= 16'b0000_0000_0000_0000;
array[47412] <= 16'b0000_0000_0000_0000;
array[47413] <= 16'b0000_0000_0000_0000;
array[47414] <= 16'b0000_0000_0000_0000;
array[47415] <= 16'b0000_0000_0000_0000;
array[47416] <= 16'b0000_0000_0000_0000;
array[47417] <= 16'b0000_0000_0000_0000;
array[47418] <= 16'b0000_0000_0000_0000;
array[47419] <= 16'b0000_0000_0000_0000;
array[47420] <= 16'b0000_0000_0000_0000;
array[47421] <= 16'b0000_0000_0000_0000;
array[47422] <= 16'b0000_0000_0000_0000;
array[47423] <= 16'b0000_0000_0000_0000;
array[47424] <= 16'b0000_0000_0000_0000;
array[47425] <= 16'b0000_0000_0000_0000;
array[47426] <= 16'b0000_0000_0000_0000;
array[47427] <= 16'b0000_0000_0000_0000;
array[47428] <= 16'b0000_0000_0000_0000;
array[47429] <= 16'b0000_0000_0000_0000;
array[47430] <= 16'b0000_0000_0000_0000;
array[47431] <= 16'b0000_0000_0000_0000;
array[47432] <= 16'b0000_0000_0000_0000;
array[47433] <= 16'b0000_0000_0000_0000;
array[47434] <= 16'b0000_0000_0000_0000;
array[47435] <= 16'b0000_0000_0000_0000;
array[47436] <= 16'b0000_0000_0000_0000;
array[47437] <= 16'b0000_0000_0000_0000;
array[47438] <= 16'b0000_0000_0000_0000;
array[47439] <= 16'b0000_0000_0000_0000;
array[47440] <= 16'b0000_0000_0000_0000;
array[47441] <= 16'b0000_0000_0000_0000;
array[47442] <= 16'b0000_0000_0000_0000;
array[47443] <= 16'b0000_0000_0000_0000;
array[47444] <= 16'b0000_0000_0000_0000;
array[47445] <= 16'b0000_0000_0000_0000;
array[47446] <= 16'b0000_0000_0000_0000;
array[47447] <= 16'b0000_0000_0000_0000;
array[47448] <= 16'b0000_0000_0000_0000;
array[47449] <= 16'b0000_0000_0000_0000;
array[47450] <= 16'b0000_0000_0000_0000;
array[47451] <= 16'b0000_0000_0000_0000;
array[47452] <= 16'b0000_0000_0000_0000;
array[47453] <= 16'b0000_0000_0000_0000;
array[47454] <= 16'b0000_0000_0000_0000;
array[47455] <= 16'b0000_0000_0000_0000;
array[47456] <= 16'b0000_0000_0000_0000;
array[47457] <= 16'b0000_0000_0000_0000;
array[47458] <= 16'b0000_0000_0000_0000;
array[47459] <= 16'b0000_0000_0000_0000;
array[47460] <= 16'b0000_0000_0000_0000;
array[47461] <= 16'b0000_0000_0000_0000;
array[47462] <= 16'b0000_0000_0000_0000;
array[47463] <= 16'b0000_0000_0000_0000;
array[47464] <= 16'b0000_0000_0000_0000;
array[47465] <= 16'b0000_0000_0000_0000;
array[47466] <= 16'b0000_0000_0000_0000;
array[47467] <= 16'b0000_0000_0000_0000;
array[47468] <= 16'b0000_0000_0000_0000;
array[47469] <= 16'b0000_0000_0000_0000;
array[47470] <= 16'b0000_0000_0000_0000;
array[47471] <= 16'b0000_0000_0000_0000;
array[47472] <= 16'b0000_0000_0000_0000;
array[47473] <= 16'b0000_0000_0000_0000;
array[47474] <= 16'b0000_0000_0000_0000;
array[47475] <= 16'b0000_0000_0000_0000;
array[47476] <= 16'b0000_0000_0000_0000;
array[47477] <= 16'b0000_0000_0000_0000;
array[47478] <= 16'b0000_0000_0000_0000;
array[47479] <= 16'b0000_0000_0000_0000;
array[47480] <= 16'b0000_0000_0000_0000;
array[47481] <= 16'b0000_0000_0000_0000;
array[47482] <= 16'b0000_0000_0000_0000;
array[47483] <= 16'b0000_0000_0000_0000;
array[47484] <= 16'b0000_0000_0000_0000;
array[47485] <= 16'b0000_0000_0000_0000;
array[47486] <= 16'b0000_0000_0000_0000;
array[47487] <= 16'b0000_0000_0000_0000;
array[47488] <= 16'b0000_0000_0000_0000;
array[47489] <= 16'b0000_0000_0000_0000;
array[47490] <= 16'b0000_0000_0000_0000;
array[47491] <= 16'b0000_0000_0000_0000;
array[47492] <= 16'b0000_0000_0000_0000;
array[47493] <= 16'b0000_0000_0000_0000;
array[47494] <= 16'b0000_0000_0000_0000;
array[47495] <= 16'b0000_0000_0000_0000;
array[47496] <= 16'b0000_0000_0000_0000;
array[47497] <= 16'b0000_0000_0000_0000;
array[47498] <= 16'b0000_0000_0000_0000;
array[47499] <= 16'b0000_0000_0000_0000;
array[47500] <= 16'b0000_0000_0000_0000;
array[47501] <= 16'b0000_0000_0000_0000;
array[47502] <= 16'b0000_0000_0000_0000;
array[47503] <= 16'b0000_0000_0000_0000;
array[47504] <= 16'b0000_0000_0000_0000;
array[47505] <= 16'b0000_0000_0000_0000;
array[47506] <= 16'b0000_0000_0000_0000;
array[47507] <= 16'b0000_0000_0000_0000;
array[47508] <= 16'b0000_0000_0000_0000;
array[47509] <= 16'b0000_0000_0000_0000;
array[47510] <= 16'b0000_0000_0000_0000;
array[47511] <= 16'b0000_0000_0000_0000;
array[47512] <= 16'b0000_0000_0000_0000;
array[47513] <= 16'b0000_0000_0000_0000;
array[47514] <= 16'b0000_0000_0000_0000;
array[47515] <= 16'b0000_0000_0000_0000;
array[47516] <= 16'b0000_0000_0000_0000;
array[47517] <= 16'b0000_0000_0000_0000;
array[47518] <= 16'b0000_0000_0000_0000;
array[47519] <= 16'b0000_0000_0000_0000;
array[47520] <= 16'b0000_0000_0000_0000;
array[47521] <= 16'b0000_0000_0000_0000;
array[47522] <= 16'b0000_0000_0000_0000;
array[47523] <= 16'b0000_0000_0000_0000;
array[47524] <= 16'b0000_0000_0000_0000;
array[47525] <= 16'b0000_0000_0000_0000;
array[47526] <= 16'b0000_0000_0000_0000;
array[47527] <= 16'b0000_0000_0000_0000;
array[47528] <= 16'b0000_0000_0000_0000;
array[47529] <= 16'b0000_0000_0000_0000;
array[47530] <= 16'b0000_0000_0000_0000;
array[47531] <= 16'b0000_0000_0000_0000;
array[47532] <= 16'b0000_0000_0000_0000;
array[47533] <= 16'b0000_0000_0000_0000;
array[47534] <= 16'b0000_0000_0000_0000;
array[47535] <= 16'b0000_0000_0000_0000;
array[47536] <= 16'b0000_0000_0000_0000;
array[47537] <= 16'b0000_0000_0000_0000;
array[47538] <= 16'b0000_0000_0000_0000;
array[47539] <= 16'b0000_0000_0000_0000;
array[47540] <= 16'b0000_0000_0000_0000;
array[47541] <= 16'b0000_0000_0000_0000;
array[47542] <= 16'b0000_0000_0000_0000;
array[47543] <= 16'b0000_0000_0000_0000;
array[47544] <= 16'b0000_0000_0000_0000;
array[47545] <= 16'b0000_0000_0000_0000;
array[47546] <= 16'b0000_0000_0000_0000;
array[47547] <= 16'b0000_0000_0000_0000;
array[47548] <= 16'b0000_0000_0000_0000;
array[47549] <= 16'b0000_0000_0000_0000;
array[47550] <= 16'b0000_0000_0000_0000;
array[47551] <= 16'b0000_0000_0000_0000;
array[47552] <= 16'b0000_0000_0000_0000;
array[47553] <= 16'b0000_0000_0000_0000;
array[47554] <= 16'b0000_0000_0000_0000;
array[47555] <= 16'b0000_0000_0000_0000;
array[47556] <= 16'b0000_0000_0000_0000;
array[47557] <= 16'b0000_0000_0000_0000;
array[47558] <= 16'b0000_0000_0000_0000;
array[47559] <= 16'b0000_0000_0000_0000;
array[47560] <= 16'b0000_0000_0000_0000;
array[47561] <= 16'b0000_0000_0000_0000;
array[47562] <= 16'b0000_0000_0000_0000;
array[47563] <= 16'b0000_0000_0000_0000;
array[47564] <= 16'b0000_0000_0000_0000;
array[47565] <= 16'b0000_0000_0000_0000;
array[47566] <= 16'b0000_0000_0000_0000;
array[47567] <= 16'b0000_0000_0000_0000;
array[47568] <= 16'b0000_0000_0000_0000;
array[47569] <= 16'b0000_0000_0000_0000;
array[47570] <= 16'b0000_0000_0000_0000;
array[47571] <= 16'b0000_0000_0000_0000;
array[47572] <= 16'b0000_0000_0000_0000;
array[47573] <= 16'b0000_0000_0000_0000;
array[47574] <= 16'b0000_0000_0000_0000;
array[47575] <= 16'b0000_0000_0000_0000;
array[47576] <= 16'b0000_0000_0000_0000;
array[47577] <= 16'b0000_0000_0000_0000;
array[47578] <= 16'b0000_0000_0000_0000;
array[47579] <= 16'b0000_0000_0000_0000;
array[47580] <= 16'b0000_0000_0000_0000;
array[47581] <= 16'b0000_0000_0000_0000;
array[47582] <= 16'b0000_0000_0000_0000;
array[47583] <= 16'b0000_0000_0000_0000;
array[47584] <= 16'b0000_0000_0000_0000;
array[47585] <= 16'b0000_0000_0000_0000;
array[47586] <= 16'b0000_0000_0000_0000;
array[47587] <= 16'b0000_0000_0000_0000;
array[47588] <= 16'b0000_0000_0000_0000;
array[47589] <= 16'b0000_0000_0000_0000;
array[47590] <= 16'b0000_0000_0000_0000;
array[47591] <= 16'b0000_0000_0000_0000;
array[47592] <= 16'b0000_0000_0000_0000;
array[47593] <= 16'b0000_0000_0000_0000;
array[47594] <= 16'b0000_0000_0000_0000;
array[47595] <= 16'b0000_0000_0000_0000;
array[47596] <= 16'b0000_0000_0000_0000;
array[47597] <= 16'b0000_0000_0000_0000;
array[47598] <= 16'b0000_0000_0000_0000;
array[47599] <= 16'b0000_0000_0000_0000;
array[47600] <= 16'b0000_0000_0000_0000;
array[47601] <= 16'b0000_0000_0000_0000;
array[47602] <= 16'b0000_0000_0000_0000;
array[47603] <= 16'b0000_0000_0000_0000;
array[47604] <= 16'b0000_0000_0000_0000;
array[47605] <= 16'b0000_0000_0000_0000;
array[47606] <= 16'b0000_0000_0000_0000;
array[47607] <= 16'b0000_0000_0000_0000;
array[47608] <= 16'b0000_0000_0000_0000;
array[47609] <= 16'b0000_0000_0000_0000;
array[47610] <= 16'b0000_0000_0000_0000;
array[47611] <= 16'b0000_0000_0000_0000;
array[47612] <= 16'b0000_0000_0000_0000;
array[47613] <= 16'b0000_0000_0000_0000;
array[47614] <= 16'b0000_0000_0000_0000;
array[47615] <= 16'b0000_0000_0000_0000;
array[47616] <= 16'b0000_0000_0000_0000;
array[47617] <= 16'b0000_0000_0000_0000;
array[47618] <= 16'b0000_0000_0000_0000;
array[47619] <= 16'b0000_0000_0000_0000;
array[47620] <= 16'b0000_0000_0000_0000;
array[47621] <= 16'b0000_0000_0000_0000;
array[47622] <= 16'b0000_0000_0000_0000;
array[47623] <= 16'b0000_0000_0000_0000;
array[47624] <= 16'b0000_0000_0000_0000;
array[47625] <= 16'b0000_0000_0000_0000;
array[47626] <= 16'b0000_0000_0000_0000;
array[47627] <= 16'b0000_0000_0000_0000;
array[47628] <= 16'b0000_0000_0000_0000;
array[47629] <= 16'b0000_0000_0000_0000;
array[47630] <= 16'b0000_0000_0000_0000;
array[47631] <= 16'b0000_0000_0000_0000;
array[47632] <= 16'b0000_0000_0000_0000;
array[47633] <= 16'b0000_0000_0000_0000;
array[47634] <= 16'b0000_0000_0000_0000;
array[47635] <= 16'b0000_0000_0000_0000;
array[47636] <= 16'b0000_0000_0000_0000;
array[47637] <= 16'b0000_0000_0000_0000;
array[47638] <= 16'b0000_0000_0000_0000;
array[47639] <= 16'b0000_0000_0000_0000;
array[47640] <= 16'b0000_0000_0000_0000;
array[47641] <= 16'b0000_0000_0000_0000;
array[47642] <= 16'b0000_0000_0000_0000;
array[47643] <= 16'b0000_0000_0000_0000;
array[47644] <= 16'b0000_0000_0000_0000;
array[47645] <= 16'b0000_0000_0000_0000;
array[47646] <= 16'b0000_0000_0000_0000;
array[47647] <= 16'b0000_0000_0000_0000;
array[47648] <= 16'b0000_0000_0000_0000;
array[47649] <= 16'b0000_0000_0000_0000;
array[47650] <= 16'b0000_0000_0000_0000;
array[47651] <= 16'b0000_0000_0000_0000;
array[47652] <= 16'b0000_0000_0000_0000;
array[47653] <= 16'b0000_0000_0000_0000;
array[47654] <= 16'b0000_0000_0000_0000;
array[47655] <= 16'b0000_0000_0000_0000;
array[47656] <= 16'b0000_0000_0000_0000;
array[47657] <= 16'b0000_0000_0000_0000;
array[47658] <= 16'b0000_0000_0000_0000;
array[47659] <= 16'b0000_0000_0000_0000;
array[47660] <= 16'b0000_0000_0000_0000;
array[47661] <= 16'b0000_0000_0000_0000;
array[47662] <= 16'b0000_0000_0000_0000;
array[47663] <= 16'b0000_0000_0000_0000;
array[47664] <= 16'b0000_0000_0000_0000;
array[47665] <= 16'b0000_0000_0000_0000;
array[47666] <= 16'b0000_0000_0000_0000;
array[47667] <= 16'b0000_0000_0000_0000;
array[47668] <= 16'b0000_0000_0000_0000;
array[47669] <= 16'b0000_0000_0000_0000;
array[47670] <= 16'b0000_0000_0000_0000;
array[47671] <= 16'b0000_0000_0000_0000;
array[47672] <= 16'b0000_0000_0000_0000;
array[47673] <= 16'b0000_0000_0000_0000;
array[47674] <= 16'b0000_0000_0000_0000;
array[47675] <= 16'b0000_0000_0000_0000;
array[47676] <= 16'b0000_0000_0000_0000;
array[47677] <= 16'b0000_0000_0000_0000;
array[47678] <= 16'b0000_0000_0000_0000;
array[47679] <= 16'b0000_0000_0000_0000;
array[47680] <= 16'b0000_0000_0000_0000;
array[47681] <= 16'b0000_0000_0000_0000;
array[47682] <= 16'b0000_0000_0000_0000;
array[47683] <= 16'b0000_0000_0000_0000;
array[47684] <= 16'b0000_0000_0000_0000;
array[47685] <= 16'b0000_0000_0000_0000;
array[47686] <= 16'b0000_0000_0000_0000;
array[47687] <= 16'b0000_0000_0000_0000;
array[47688] <= 16'b0000_0000_0000_0000;
array[47689] <= 16'b0000_0000_0000_0000;
array[47690] <= 16'b0000_0000_0000_0000;
array[47691] <= 16'b0000_0000_0000_0000;
array[47692] <= 16'b0000_0000_0000_0000;
array[47693] <= 16'b0000_0000_0000_0000;
array[47694] <= 16'b0000_0000_0000_0000;
array[47695] <= 16'b0000_0000_0000_0000;
array[47696] <= 16'b0000_0000_0000_0000;
array[47697] <= 16'b0000_0000_0000_0000;
array[47698] <= 16'b0000_0000_0000_0000;
array[47699] <= 16'b0000_0000_0000_0000;
array[47700] <= 16'b0000_0000_0000_0000;
array[47701] <= 16'b0000_0000_0000_0000;
array[47702] <= 16'b0000_0000_0000_0000;
array[47703] <= 16'b0000_0000_0000_0000;
array[47704] <= 16'b0000_0000_0000_0000;
array[47705] <= 16'b0000_0000_0000_0000;
array[47706] <= 16'b0000_0000_0000_0000;
array[47707] <= 16'b0000_0000_0000_0000;
array[47708] <= 16'b0000_0000_0000_0000;
array[47709] <= 16'b0000_0000_0000_0000;
array[47710] <= 16'b0000_0000_0000_0000;
array[47711] <= 16'b0000_0000_0000_0000;
array[47712] <= 16'b0000_0000_0000_0000;
array[47713] <= 16'b0000_0000_0000_0000;
array[47714] <= 16'b0000_0000_0000_0000;
array[47715] <= 16'b0000_0000_0000_0000;
array[47716] <= 16'b0000_0000_0000_0000;
array[47717] <= 16'b0000_0000_0000_0000;
array[47718] <= 16'b0000_0000_0000_0000;
array[47719] <= 16'b0000_0000_0000_0000;
array[47720] <= 16'b0000_0000_0000_0000;
array[47721] <= 16'b0000_0000_0000_0000;
array[47722] <= 16'b0000_0000_0000_0000;
array[47723] <= 16'b0000_0000_0000_0000;
array[47724] <= 16'b0000_0000_0000_0000;
array[47725] <= 16'b0000_0000_0000_0000;
array[47726] <= 16'b0000_0000_0000_0000;
array[47727] <= 16'b0000_0000_0000_0000;
array[47728] <= 16'b0000_0000_0000_0000;
array[47729] <= 16'b0000_0000_0000_0000;
array[47730] <= 16'b0000_0000_0000_0000;
array[47731] <= 16'b0000_0000_0000_0000;
array[47732] <= 16'b0000_0000_0000_0000;
array[47733] <= 16'b0000_0000_0000_0000;
array[47734] <= 16'b0000_0000_0000_0000;
array[47735] <= 16'b0000_0000_0000_0000;
array[47736] <= 16'b0000_0000_0000_0000;
array[47737] <= 16'b0000_0000_0000_0000;
array[47738] <= 16'b0000_0000_0000_0000;
array[47739] <= 16'b0000_0000_0000_0000;
array[47740] <= 16'b0000_0000_0000_0000;
array[47741] <= 16'b0000_0000_0000_0000;
array[47742] <= 16'b0000_0000_0000_0000;
array[47743] <= 16'b0000_0000_0000_0000;
array[47744] <= 16'b0000_0000_0000_0000;
array[47745] <= 16'b0000_0000_0000_0000;
array[47746] <= 16'b0000_0000_0000_0000;
array[47747] <= 16'b0000_0000_0000_0000;
array[47748] <= 16'b0000_0000_0000_0000;
array[47749] <= 16'b0000_0000_0000_0000;
array[47750] <= 16'b0000_0000_0000_0000;
array[47751] <= 16'b0000_0000_0000_0000;
array[47752] <= 16'b0000_0000_0000_0000;
array[47753] <= 16'b0000_0000_0000_0000;
array[47754] <= 16'b0000_0000_0000_0000;
array[47755] <= 16'b0000_0000_0000_0000;
array[47756] <= 16'b0000_0000_0000_0000;
array[47757] <= 16'b0000_0000_0000_0000;
array[47758] <= 16'b0000_0000_0000_0000;
array[47759] <= 16'b0000_0000_0000_0000;
array[47760] <= 16'b0000_0000_0000_0000;
array[47761] <= 16'b0000_0000_0000_0000;
array[47762] <= 16'b0000_0000_0000_0000;
array[47763] <= 16'b0000_0000_0000_0000;
array[47764] <= 16'b0000_0000_0000_0000;
array[47765] <= 16'b0000_0000_0000_0000;
array[47766] <= 16'b0000_0000_0000_0000;
array[47767] <= 16'b0000_0000_0000_0000;
array[47768] <= 16'b0000_0000_0000_0000;
array[47769] <= 16'b0000_0000_0000_0000;
array[47770] <= 16'b0000_0000_0000_0000;
array[47771] <= 16'b0000_0000_0000_0000;
array[47772] <= 16'b0000_0000_0000_0000;
array[47773] <= 16'b0000_0000_0000_0000;
array[47774] <= 16'b0000_0000_0000_0000;
array[47775] <= 16'b0000_0000_0000_0000;
array[47776] <= 16'b0000_0000_0000_0000;
array[47777] <= 16'b0000_0000_0000_0000;
array[47778] <= 16'b0000_0000_0000_0000;
array[47779] <= 16'b0000_0000_0000_0000;
array[47780] <= 16'b0000_0000_0000_0000;
array[47781] <= 16'b0000_0000_0000_0000;
array[47782] <= 16'b0000_0000_0000_0000;
array[47783] <= 16'b0000_0000_0000_0000;
array[47784] <= 16'b0000_0000_0000_0000;
array[47785] <= 16'b0000_0000_0000_0000;
array[47786] <= 16'b0000_0000_0000_0000;
array[47787] <= 16'b0000_0000_0000_0000;
array[47788] <= 16'b0000_0000_0000_0000;
array[47789] <= 16'b0000_0000_0000_0000;
array[47790] <= 16'b0000_0000_0000_0000;
array[47791] <= 16'b0000_0000_0000_0000;
array[47792] <= 16'b0000_0000_0000_0000;
array[47793] <= 16'b0000_0000_0000_0000;
array[47794] <= 16'b0000_0000_0000_0000;
array[47795] <= 16'b0000_0000_0000_0000;
array[47796] <= 16'b0000_0000_0000_0000;
array[47797] <= 16'b0000_0000_0000_0000;
array[47798] <= 16'b0000_0000_0000_0000;
array[47799] <= 16'b0000_0000_0000_0000;
array[47800] <= 16'b0000_0000_0000_0000;
array[47801] <= 16'b0000_0000_0000_0000;
array[47802] <= 16'b0000_0000_0000_0000;
array[47803] <= 16'b0000_0000_0000_0000;
array[47804] <= 16'b0000_0000_0000_0000;
array[47805] <= 16'b0000_0000_0000_0000;
array[47806] <= 16'b0000_0000_0000_0000;
array[47807] <= 16'b0000_0000_0000_0000;
array[47808] <= 16'b0000_0000_0000_0000;
array[47809] <= 16'b0000_0000_0000_0000;
array[47810] <= 16'b0000_0000_0000_0000;
array[47811] <= 16'b0000_0000_0000_0000;
array[47812] <= 16'b0000_0000_0000_0000;
array[47813] <= 16'b0000_0000_0000_0000;
array[47814] <= 16'b0000_0000_0000_0000;
array[47815] <= 16'b0000_0000_0000_0000;
array[47816] <= 16'b0000_0000_0000_0000;
array[47817] <= 16'b0000_0000_0000_0000;
array[47818] <= 16'b0000_0000_0000_0000;
array[47819] <= 16'b0000_0000_0000_0000;
array[47820] <= 16'b0000_0000_0000_0000;
array[47821] <= 16'b0000_0000_0000_0000;
array[47822] <= 16'b0000_0000_0000_0000;
array[47823] <= 16'b0000_0000_0000_0000;
array[47824] <= 16'b0000_0000_0000_0000;
array[47825] <= 16'b0000_0000_0000_0000;
array[47826] <= 16'b0000_0000_0000_0000;
array[47827] <= 16'b0000_0000_0000_0000;
array[47828] <= 16'b0000_0000_0000_0000;
array[47829] <= 16'b0000_0000_0000_0000;
array[47830] <= 16'b0000_0000_0000_0000;
array[47831] <= 16'b0000_0000_0000_0000;
array[47832] <= 16'b0000_0000_0000_0000;
array[47833] <= 16'b0000_0000_0000_0000;
array[47834] <= 16'b0000_0000_0000_0000;
array[47835] <= 16'b0000_0000_0000_0000;
array[47836] <= 16'b0000_0000_0000_0000;
array[47837] <= 16'b0000_0000_0000_0000;
array[47838] <= 16'b0000_0000_0000_0000;
array[47839] <= 16'b0000_0000_0000_0000;
array[47840] <= 16'b0000_0000_0000_0000;
array[47841] <= 16'b0000_0000_0000_0000;
array[47842] <= 16'b0000_0000_0000_0000;
array[47843] <= 16'b0000_0000_0000_0000;
array[47844] <= 16'b0000_0000_0000_0000;
array[47845] <= 16'b0000_0000_0000_0000;
array[47846] <= 16'b0000_0000_0000_0000;
array[47847] <= 16'b0000_0000_0000_0000;
array[47848] <= 16'b0000_0000_0000_0000;
array[47849] <= 16'b0000_0000_0000_0000;
array[47850] <= 16'b0000_0000_0000_0000;
array[47851] <= 16'b0000_0000_0000_0000;
array[47852] <= 16'b0000_0000_0000_0000;
array[47853] <= 16'b0000_0000_0000_0000;
array[47854] <= 16'b0000_0000_0000_0000;
array[47855] <= 16'b0000_0000_0000_0000;
array[47856] <= 16'b0000_0000_0000_0000;
array[47857] <= 16'b0000_0000_0000_0000;
array[47858] <= 16'b0000_0000_0000_0000;
array[47859] <= 16'b0000_0000_0000_0000;
array[47860] <= 16'b0000_0000_0000_0000;
array[47861] <= 16'b0000_0000_0000_0000;
array[47862] <= 16'b0000_0000_0000_0000;
array[47863] <= 16'b0000_0000_0000_0000;
array[47864] <= 16'b0000_0000_0000_0000;
array[47865] <= 16'b0000_0000_0000_0000;
array[47866] <= 16'b0000_0000_0000_0000;
array[47867] <= 16'b0000_0000_0000_0000;
array[47868] <= 16'b0000_0000_0000_0000;
array[47869] <= 16'b0000_0000_0000_0000;
array[47870] <= 16'b0000_0000_0000_0000;
array[47871] <= 16'b0000_0000_0000_0000;
array[47872] <= 16'b0000_0000_0000_0000;
array[47873] <= 16'b0000_0000_0000_0000;
array[47874] <= 16'b0000_0000_0000_0000;
array[47875] <= 16'b0000_0000_0000_0000;
array[47876] <= 16'b0000_0000_0000_0000;
array[47877] <= 16'b0000_0000_0000_0000;
array[47878] <= 16'b0000_0000_0000_0000;
array[47879] <= 16'b0000_0000_0000_0000;
array[47880] <= 16'b0000_0000_0000_0000;
array[47881] <= 16'b0000_0000_0000_0000;
array[47882] <= 16'b0000_0000_0000_0000;
array[47883] <= 16'b0000_0000_0000_0000;
array[47884] <= 16'b0000_0000_0000_0000;
array[47885] <= 16'b0000_0000_0000_0000;
array[47886] <= 16'b0000_0000_0000_0000;
array[47887] <= 16'b0000_0000_0000_0000;
array[47888] <= 16'b0000_0000_0000_0000;
array[47889] <= 16'b0000_0000_0000_0000;
array[47890] <= 16'b0000_0000_0000_0000;
array[47891] <= 16'b0000_0000_0000_0000;
array[47892] <= 16'b0000_0000_0000_0000;
array[47893] <= 16'b0000_0000_0000_0000;
array[47894] <= 16'b0000_0000_0000_0000;
array[47895] <= 16'b0000_0000_0000_0000;
array[47896] <= 16'b0000_0000_0000_0000;
array[47897] <= 16'b0000_0000_0000_0000;
array[47898] <= 16'b0000_0000_0000_0000;
array[47899] <= 16'b0000_0000_0000_0000;
array[47900] <= 16'b0000_0000_0000_0000;
array[47901] <= 16'b0000_0000_0000_0000;
array[47902] <= 16'b0000_0000_0000_0000;
array[47903] <= 16'b0000_0000_0000_0000;
array[47904] <= 16'b0000_0000_0000_0000;
array[47905] <= 16'b0000_0000_0000_0000;
array[47906] <= 16'b0000_0000_0000_0000;
array[47907] <= 16'b0000_0000_0000_0000;
array[47908] <= 16'b0000_0000_0000_0000;
array[47909] <= 16'b0000_0000_0000_0000;
array[47910] <= 16'b0000_0000_0000_0000;
array[47911] <= 16'b0000_0000_0000_0000;
array[47912] <= 16'b0000_0000_0000_0000;
array[47913] <= 16'b0000_0000_0000_0000;
array[47914] <= 16'b0000_0000_0000_0000;
array[47915] <= 16'b0000_0000_0000_0000;
array[47916] <= 16'b0000_0000_0000_0000;
array[47917] <= 16'b0000_0000_0000_0000;
array[47918] <= 16'b0000_0000_0000_0000;
array[47919] <= 16'b0000_0000_0000_0000;
array[47920] <= 16'b0000_0000_0000_0000;
array[47921] <= 16'b0000_0000_0000_0000;
array[47922] <= 16'b0000_0000_0000_0000;
array[47923] <= 16'b0000_0000_0000_0000;
array[47924] <= 16'b0000_0000_0000_0000;
array[47925] <= 16'b0000_0000_0000_0000;
array[47926] <= 16'b0000_0000_0000_0000;
array[47927] <= 16'b0000_0000_0000_0000;
array[47928] <= 16'b0000_0000_0000_0000;
array[47929] <= 16'b0000_0000_0000_0000;
array[47930] <= 16'b0000_0000_0000_0000;
array[47931] <= 16'b0000_0000_0000_0000;
array[47932] <= 16'b0000_0000_0000_0000;
array[47933] <= 16'b0000_0000_0000_0000;
array[47934] <= 16'b0000_0000_0000_0000;
array[47935] <= 16'b0000_0000_0000_0000;
array[47936] <= 16'b0000_0000_0000_0000;
array[47937] <= 16'b0000_0000_0000_0000;
array[47938] <= 16'b0000_0000_0000_0000;
array[47939] <= 16'b0000_0000_0000_0000;
array[47940] <= 16'b0000_0000_0000_0000;
array[47941] <= 16'b0000_0000_0000_0000;
array[47942] <= 16'b0000_0000_0000_0000;
array[47943] <= 16'b0000_0000_0000_0000;
array[47944] <= 16'b0000_0000_0000_0000;
array[47945] <= 16'b0000_0000_0000_0000;
array[47946] <= 16'b0000_0000_0000_0000;
array[47947] <= 16'b0000_0000_0000_0000;
array[47948] <= 16'b0000_0000_0000_0000;
array[47949] <= 16'b0000_0000_0000_0000;
array[47950] <= 16'b0000_0000_0000_0000;
array[47951] <= 16'b0000_0000_0000_0000;
array[47952] <= 16'b0000_0000_0000_0000;
array[47953] <= 16'b0000_0000_0000_0000;
array[47954] <= 16'b0000_0000_0000_0000;
array[47955] <= 16'b0000_0000_0000_0000;
array[47956] <= 16'b0000_0000_0000_0000;
array[47957] <= 16'b0000_0000_0000_0000;
array[47958] <= 16'b0000_0000_0000_0000;
array[47959] <= 16'b0000_0000_0000_0000;
array[47960] <= 16'b0000_0000_0000_0000;
array[47961] <= 16'b0000_0000_0000_0000;
array[47962] <= 16'b0000_0000_0000_0000;
array[47963] <= 16'b0000_0000_0000_0000;
array[47964] <= 16'b0000_0000_0000_0000;
array[47965] <= 16'b0000_0000_0000_0000;
array[47966] <= 16'b0000_0000_0000_0000;
array[47967] <= 16'b0000_0000_0000_0000;
array[47968] <= 16'b0000_0000_0000_0000;
array[47969] <= 16'b0000_0000_0000_0000;
array[47970] <= 16'b0000_0000_0000_0000;
array[47971] <= 16'b0000_0000_0000_0000;
array[47972] <= 16'b0000_0000_0000_0000;
array[47973] <= 16'b0000_0000_0000_0000;
array[47974] <= 16'b0000_0000_0000_0000;
array[47975] <= 16'b0000_0000_0000_0000;
array[47976] <= 16'b0000_0000_0000_0000;
array[47977] <= 16'b0000_0000_0000_0000;
array[47978] <= 16'b0000_0000_0000_0000;
array[47979] <= 16'b0000_0000_0000_0000;
array[47980] <= 16'b0000_0000_0000_0000;
array[47981] <= 16'b0000_0000_0000_0000;
array[47982] <= 16'b0000_0000_0000_0000;
array[47983] <= 16'b0000_0000_0000_0000;
array[47984] <= 16'b0000_0000_0000_0000;
array[47985] <= 16'b0000_0000_0000_0000;
array[47986] <= 16'b0000_0000_0000_0000;
array[47987] <= 16'b0000_0000_0000_0000;
array[47988] <= 16'b0000_0000_0000_0000;
array[47989] <= 16'b0000_0000_0000_0000;
array[47990] <= 16'b0000_0000_0000_0000;
array[47991] <= 16'b0000_0000_0000_0000;
array[47992] <= 16'b0000_0000_0000_0000;
array[47993] <= 16'b0000_0000_0000_0000;
array[47994] <= 16'b0000_0000_0000_0000;
array[47995] <= 16'b0000_0000_0000_0000;
array[47996] <= 16'b0000_0000_0000_0000;
array[47997] <= 16'b0000_0000_0000_0000;
array[47998] <= 16'b0000_0000_0000_0000;
array[47999] <= 16'b0000_0000_0000_0000;
array[48000] <= 16'b0000_0000_0000_0000;
array[48001] <= 16'b0000_0000_0000_0000;
array[48002] <= 16'b0000_0000_0000_0000;
array[48003] <= 16'b0000_0000_0000_0000;
array[48004] <= 16'b0000_0000_0000_0000;
array[48005] <= 16'b0000_0000_0000_0000;
array[48006] <= 16'b0000_0000_0000_0000;
array[48007] <= 16'b0000_0000_0000_0000;
array[48008] <= 16'b0000_0000_0000_0000;
array[48009] <= 16'b0000_0000_0000_0000;
array[48010] <= 16'b0000_0000_0000_0000;
array[48011] <= 16'b0000_0000_0000_0000;
array[48012] <= 16'b0000_0000_0000_0000;
array[48013] <= 16'b0000_0000_0000_0000;
array[48014] <= 16'b0000_0000_0000_0000;
array[48015] <= 16'b0000_0000_0000_0000;
array[48016] <= 16'b0000_0000_0000_0000;
array[48017] <= 16'b0000_0000_0000_0000;
array[48018] <= 16'b0000_0000_0000_0000;
array[48019] <= 16'b0000_0000_0000_0000;
array[48020] <= 16'b0000_0000_0000_0000;
array[48021] <= 16'b0000_0000_0000_0000;
array[48022] <= 16'b0000_0000_0000_0000;
array[48023] <= 16'b0000_0000_0000_0000;
array[48024] <= 16'b0000_0000_0000_0000;
array[48025] <= 16'b0000_0000_0000_0000;
array[48026] <= 16'b0000_0000_0000_0000;
array[48027] <= 16'b0000_0000_0000_0000;
array[48028] <= 16'b0000_0000_0000_0000;
array[48029] <= 16'b0000_0000_0000_0000;
array[48030] <= 16'b0000_0000_0000_0000;
array[48031] <= 16'b0000_0000_0000_0000;
array[48032] <= 16'b0000_0000_0000_0000;
array[48033] <= 16'b0000_0000_0000_0000;
array[48034] <= 16'b0000_0000_0000_0000;
array[48035] <= 16'b0000_0000_0000_0000;
array[48036] <= 16'b0000_0000_0000_0000;
array[48037] <= 16'b0000_0000_0000_0000;
array[48038] <= 16'b0000_0000_0000_0000;
array[48039] <= 16'b0000_0000_0000_0000;
array[48040] <= 16'b0000_0000_0000_0000;
array[48041] <= 16'b0000_0000_0000_0000;
array[48042] <= 16'b0000_0000_0000_0000;
array[48043] <= 16'b0000_0000_0000_0000;
array[48044] <= 16'b0000_0000_0000_0000;
array[48045] <= 16'b0000_0000_0000_0000;
array[48046] <= 16'b0000_0000_0000_0000;
array[48047] <= 16'b0000_0000_0000_0000;
array[48048] <= 16'b0000_0000_0000_0000;
array[48049] <= 16'b0000_0000_0000_0000;
array[48050] <= 16'b0000_0000_0000_0000;
array[48051] <= 16'b0000_0000_0000_0000;
array[48052] <= 16'b0000_0000_0000_0000;
array[48053] <= 16'b0000_0000_0000_0000;
array[48054] <= 16'b0000_0000_0000_0000;
array[48055] <= 16'b0000_0000_0000_0000;
array[48056] <= 16'b0000_0000_0000_0000;
array[48057] <= 16'b0000_0000_0000_0000;
array[48058] <= 16'b0000_0000_0000_0000;
array[48059] <= 16'b0000_0000_0000_0000;
array[48060] <= 16'b0000_0000_0000_0000;
array[48061] <= 16'b0000_0000_0000_0000;
array[48062] <= 16'b0000_0000_0000_0000;
array[48063] <= 16'b0000_0000_0000_0000;
array[48064] <= 16'b0000_0000_0000_0000;
array[48065] <= 16'b0000_0000_0000_0000;
array[48066] <= 16'b0000_0000_0000_0000;
array[48067] <= 16'b0000_0000_0000_0000;
array[48068] <= 16'b0000_0000_0000_0000;
array[48069] <= 16'b0000_0000_0000_0000;
array[48070] <= 16'b0000_0000_0000_0000;
array[48071] <= 16'b0000_0000_0000_0000;
array[48072] <= 16'b0000_0000_0000_0000;
array[48073] <= 16'b0000_0000_0000_0000;
array[48074] <= 16'b0000_0000_0000_0000;
array[48075] <= 16'b0000_0000_0000_0000;
array[48076] <= 16'b0000_0000_0000_0000;
array[48077] <= 16'b0000_0000_0000_0000;
array[48078] <= 16'b0000_0000_0000_0000;
array[48079] <= 16'b0000_0000_0000_0000;
array[48080] <= 16'b0000_0000_0000_0000;
array[48081] <= 16'b0000_0000_0000_0000;
array[48082] <= 16'b0000_0000_0000_0000;
array[48083] <= 16'b0000_0000_0000_0000;
array[48084] <= 16'b0000_0000_0000_0000;
array[48085] <= 16'b0000_0000_0000_0000;
array[48086] <= 16'b0000_0000_0000_0000;
array[48087] <= 16'b0000_0000_0000_0000;
array[48088] <= 16'b0000_0000_0000_0000;
array[48089] <= 16'b0000_0000_0000_0000;
array[48090] <= 16'b0000_0000_0000_0000;
array[48091] <= 16'b0000_0000_0000_0000;
array[48092] <= 16'b0000_0000_0000_0000;
array[48093] <= 16'b0000_0000_0000_0000;
array[48094] <= 16'b0000_0000_0000_0000;
array[48095] <= 16'b0000_0000_0000_0000;
array[48096] <= 16'b0000_0000_0000_0000;
array[48097] <= 16'b0000_0000_0000_0000;
array[48098] <= 16'b0000_0000_0000_0000;
array[48099] <= 16'b0000_0000_0000_0000;
array[48100] <= 16'b0000_0000_0000_0000;
array[48101] <= 16'b0000_0000_0000_0000;
array[48102] <= 16'b0000_0000_0000_0000;
array[48103] <= 16'b0000_0000_0000_0000;
array[48104] <= 16'b0000_0000_0000_0000;
array[48105] <= 16'b0000_0000_0000_0000;
array[48106] <= 16'b0000_0000_0000_0000;
array[48107] <= 16'b0000_0000_0000_0000;
array[48108] <= 16'b0000_0000_0000_0000;
array[48109] <= 16'b0000_0000_0000_0000;
array[48110] <= 16'b0000_0000_0000_0000;
array[48111] <= 16'b0000_0000_0000_0000;
array[48112] <= 16'b0000_0000_0000_0000;
array[48113] <= 16'b0000_0000_0000_0000;
array[48114] <= 16'b0000_0000_0000_0000;
array[48115] <= 16'b0000_0000_0000_0000;
array[48116] <= 16'b0000_0000_0000_0000;
array[48117] <= 16'b0000_0000_0000_0000;
array[48118] <= 16'b0000_0000_0000_0000;
array[48119] <= 16'b0000_0000_0000_0000;
array[48120] <= 16'b0000_0000_0000_0000;
array[48121] <= 16'b0000_0000_0000_0000;
array[48122] <= 16'b0000_0000_0000_0000;
array[48123] <= 16'b0000_0000_0000_0000;
array[48124] <= 16'b0000_0000_0000_0000;
array[48125] <= 16'b0000_0000_0000_0000;
array[48126] <= 16'b0000_0000_0000_0000;
array[48127] <= 16'b0000_0000_0000_0000;
array[48128] <= 16'b0000_0000_0000_0000;
array[48129] <= 16'b0000_0000_0000_0000;
array[48130] <= 16'b0000_0000_0000_0000;
array[48131] <= 16'b0000_0000_0000_0000;
array[48132] <= 16'b0000_0000_0000_0000;
array[48133] <= 16'b0000_0000_0000_0000;
array[48134] <= 16'b0000_0000_0000_0000;
array[48135] <= 16'b0000_0000_0000_0000;
array[48136] <= 16'b0000_0000_0000_0000;
array[48137] <= 16'b0000_0000_0000_0000;
array[48138] <= 16'b0000_0000_0000_0000;
array[48139] <= 16'b0000_0000_0000_0000;
array[48140] <= 16'b0000_0000_0000_0000;
array[48141] <= 16'b0000_0000_0000_0000;
array[48142] <= 16'b0000_0000_0000_0000;
array[48143] <= 16'b0000_0000_0000_0000;
array[48144] <= 16'b0000_0000_0000_0000;
array[48145] <= 16'b0000_0000_0000_0000;
array[48146] <= 16'b0000_0000_0000_0000;
array[48147] <= 16'b0000_0000_0000_0000;
array[48148] <= 16'b0000_0000_0000_0000;
array[48149] <= 16'b0000_0000_0000_0000;
array[48150] <= 16'b0000_0000_0000_0000;
array[48151] <= 16'b0000_0000_0000_0000;
array[48152] <= 16'b0000_0000_0000_0000;
array[48153] <= 16'b0000_0000_0000_0000;
array[48154] <= 16'b0000_0000_0000_0000;
array[48155] <= 16'b0000_0000_0000_0000;
array[48156] <= 16'b0000_0000_0000_0000;
array[48157] <= 16'b0000_0000_0000_0000;
array[48158] <= 16'b0000_0000_0000_0000;
array[48159] <= 16'b0000_0000_0000_0000;
array[48160] <= 16'b0000_0000_0000_0000;
array[48161] <= 16'b0000_0000_0000_0000;
array[48162] <= 16'b0000_0000_0000_0000;
array[48163] <= 16'b0000_0000_0000_0000;
array[48164] <= 16'b0000_0000_0000_0000;
array[48165] <= 16'b0000_0000_0000_0000;
array[48166] <= 16'b0000_0000_0000_0000;
array[48167] <= 16'b0000_0000_0000_0000;
array[48168] <= 16'b0000_0000_0000_0000;
array[48169] <= 16'b0000_0000_0000_0000;
array[48170] <= 16'b0000_0000_0000_0000;
array[48171] <= 16'b0000_0000_0000_0000;
array[48172] <= 16'b0000_0000_0000_0000;
array[48173] <= 16'b0000_0000_0000_0000;
array[48174] <= 16'b0000_0000_0000_0000;
array[48175] <= 16'b0000_0000_0000_0000;
array[48176] <= 16'b0000_0000_0000_0000;
array[48177] <= 16'b0000_0000_0000_0000;
array[48178] <= 16'b0000_0000_0000_0000;
array[48179] <= 16'b0000_0000_0000_0000;
array[48180] <= 16'b0000_0000_0000_0000;
array[48181] <= 16'b0000_0000_0000_0000;
array[48182] <= 16'b0000_0000_0000_0000;
array[48183] <= 16'b0000_0000_0000_0000;
array[48184] <= 16'b0000_0000_0000_0000;
array[48185] <= 16'b0000_0000_0000_0000;
array[48186] <= 16'b0000_0000_0000_0000;
array[48187] <= 16'b0000_0000_0000_0000;
array[48188] <= 16'b0000_0000_0000_0000;
array[48189] <= 16'b0000_0000_0000_0000;
array[48190] <= 16'b0000_0000_0000_0000;
array[48191] <= 16'b0000_0000_0000_0000;
array[48192] <= 16'b0000_0000_0000_0000;
array[48193] <= 16'b0000_0000_0000_0000;
array[48194] <= 16'b0000_0000_0000_0000;
array[48195] <= 16'b0000_0000_0000_0000;
array[48196] <= 16'b0000_0000_0000_0000;
array[48197] <= 16'b0000_0000_0000_0000;
array[48198] <= 16'b0000_0000_0000_0000;
array[48199] <= 16'b0000_0000_0000_0000;
array[48200] <= 16'b0000_0000_0000_0000;
array[48201] <= 16'b0000_0000_0000_0000;
array[48202] <= 16'b0000_0000_0000_0000;
array[48203] <= 16'b0000_0000_0000_0000;
array[48204] <= 16'b0000_0000_0000_0000;
array[48205] <= 16'b0000_0000_0000_0000;
array[48206] <= 16'b0000_0000_0000_0000;
array[48207] <= 16'b0000_0000_0000_0000;
array[48208] <= 16'b0000_0000_0000_0000;
array[48209] <= 16'b0000_0000_0000_0000;
array[48210] <= 16'b0000_0000_0000_0000;
array[48211] <= 16'b0000_0000_0000_0000;
array[48212] <= 16'b0000_0000_0000_0000;
array[48213] <= 16'b0000_0000_0000_0000;
array[48214] <= 16'b0000_0000_0000_0000;
array[48215] <= 16'b0000_0000_0000_0000;
array[48216] <= 16'b0000_0000_0000_0000;
array[48217] <= 16'b0000_0000_0000_0000;
array[48218] <= 16'b0000_0000_0000_0000;
array[48219] <= 16'b0000_0000_0000_0000;
array[48220] <= 16'b0000_0000_0000_0000;
array[48221] <= 16'b0000_0000_0000_0000;
array[48222] <= 16'b0000_0000_0000_0000;
array[48223] <= 16'b0000_0000_0000_0000;
array[48224] <= 16'b0000_0000_0000_0000;
array[48225] <= 16'b0000_0000_0000_0000;
array[48226] <= 16'b0000_0000_0000_0000;
array[48227] <= 16'b0000_0000_0000_0000;
array[48228] <= 16'b0000_0000_0000_0000;
array[48229] <= 16'b0000_0000_0000_0000;
array[48230] <= 16'b0000_0000_0000_0000;
array[48231] <= 16'b0000_0000_0000_0000;
array[48232] <= 16'b0000_0000_0000_0000;
array[48233] <= 16'b0000_0000_0000_0000;
array[48234] <= 16'b0000_0000_0000_0000;
array[48235] <= 16'b0000_0000_0000_0000;
array[48236] <= 16'b0000_0000_0000_0000;
array[48237] <= 16'b0000_0000_0000_0000;
array[48238] <= 16'b0000_0000_0000_0000;
array[48239] <= 16'b0000_0000_0000_0000;
array[48240] <= 16'b0000_0000_0000_0000;
array[48241] <= 16'b0000_0000_0000_0000;
array[48242] <= 16'b0000_0000_0000_0000;
array[48243] <= 16'b0000_0000_0000_0000;
array[48244] <= 16'b0000_0000_0000_0000;
array[48245] <= 16'b0000_0000_0000_0000;
array[48246] <= 16'b0000_0000_0000_0000;
array[48247] <= 16'b0000_0000_0000_0000;
array[48248] <= 16'b0000_0000_0000_0000;
array[48249] <= 16'b0000_0000_0000_0000;
array[48250] <= 16'b0000_0000_0000_0000;
array[48251] <= 16'b0000_0000_0000_0000;
array[48252] <= 16'b0000_0000_0000_0000;
array[48253] <= 16'b0000_0000_0000_0000;
array[48254] <= 16'b0000_0000_0000_0000;
array[48255] <= 16'b0000_0000_0000_0000;
array[48256] <= 16'b0000_0000_0000_0000;
array[48257] <= 16'b0000_0000_0000_0000;
array[48258] <= 16'b0000_0000_0000_0000;
array[48259] <= 16'b0000_0000_0000_0000;
array[48260] <= 16'b0000_0000_0000_0000;
array[48261] <= 16'b0000_0000_0000_0000;
array[48262] <= 16'b0000_0000_0000_0000;
array[48263] <= 16'b0000_0000_0000_0000;
array[48264] <= 16'b0000_0000_0000_0000;
array[48265] <= 16'b0000_0000_0000_0000;
array[48266] <= 16'b0000_0000_0000_0000;
array[48267] <= 16'b0000_0000_0000_0000;
array[48268] <= 16'b0000_0000_0000_0000;
array[48269] <= 16'b0000_0000_0000_0000;
array[48270] <= 16'b0000_0000_0000_0000;
array[48271] <= 16'b0000_0000_0000_0000;
array[48272] <= 16'b0000_0000_0000_0000;
array[48273] <= 16'b0000_0000_0000_0000;
array[48274] <= 16'b0000_0000_0000_0000;
array[48275] <= 16'b0000_0000_0000_0000;
array[48276] <= 16'b0000_0000_0000_0000;
array[48277] <= 16'b0000_0000_0000_0000;
array[48278] <= 16'b0000_0000_0000_0000;
array[48279] <= 16'b0000_0000_0000_0000;
array[48280] <= 16'b0000_0000_0000_0000;
array[48281] <= 16'b0000_0000_0000_0000;
array[48282] <= 16'b0000_0000_0000_0000;
array[48283] <= 16'b0000_0000_0000_0000;
array[48284] <= 16'b0000_0000_0000_0000;
array[48285] <= 16'b0000_0000_0000_0000;
array[48286] <= 16'b0000_0000_0000_0000;
array[48287] <= 16'b0000_0000_0000_0000;
array[48288] <= 16'b0000_0000_0000_0000;
array[48289] <= 16'b0000_0000_0000_0000;
array[48290] <= 16'b0000_0000_0000_0000;
array[48291] <= 16'b0000_0000_0000_0000;
array[48292] <= 16'b0000_0000_0000_0000;
array[48293] <= 16'b0000_0000_0000_0000;
array[48294] <= 16'b0000_0000_0000_0000;
array[48295] <= 16'b0000_0000_0000_0000;
array[48296] <= 16'b0000_0000_0000_0000;
array[48297] <= 16'b0000_0000_0000_0000;
array[48298] <= 16'b0000_0000_0000_0000;
array[48299] <= 16'b0000_0000_0000_0000;
array[48300] <= 16'b0000_0000_0000_0000;
array[48301] <= 16'b0000_0000_0000_0000;
array[48302] <= 16'b0000_0000_0000_0000;
array[48303] <= 16'b0000_0000_0000_0000;
array[48304] <= 16'b0000_0000_0000_0000;
array[48305] <= 16'b0000_0000_0000_0000;
array[48306] <= 16'b0000_0000_0000_0000;
array[48307] <= 16'b0000_0000_0000_0000;
array[48308] <= 16'b0000_0000_0000_0000;
array[48309] <= 16'b0000_0000_0000_0000;
array[48310] <= 16'b0000_0000_0000_0000;
array[48311] <= 16'b0000_0000_0000_0000;
array[48312] <= 16'b0000_0000_0000_0000;
array[48313] <= 16'b0000_0000_0000_0000;
array[48314] <= 16'b0000_0000_0000_0000;
array[48315] <= 16'b0000_0000_0000_0000;
array[48316] <= 16'b0000_0000_0000_0000;
array[48317] <= 16'b0000_0000_0000_0000;
array[48318] <= 16'b0000_0000_0000_0000;
array[48319] <= 16'b0000_0000_0000_0000;
array[48320] <= 16'b0000_0000_0000_0000;
array[48321] <= 16'b0000_0000_0000_0000;
array[48322] <= 16'b0000_0000_0000_0000;
array[48323] <= 16'b0000_0000_0000_0000;
array[48324] <= 16'b0000_0000_0000_0000;
array[48325] <= 16'b0000_0000_0000_0000;
array[48326] <= 16'b0000_0000_0000_0000;
array[48327] <= 16'b0000_0000_0000_0000;
array[48328] <= 16'b0000_0000_0000_0000;
array[48329] <= 16'b0000_0000_0000_0000;
array[48330] <= 16'b0000_0000_0000_0000;
array[48331] <= 16'b0000_0000_0000_0000;
array[48332] <= 16'b0000_0000_0000_0000;
array[48333] <= 16'b0000_0000_0000_0000;
array[48334] <= 16'b0000_0000_0000_0000;
array[48335] <= 16'b0000_0000_0000_0000;
array[48336] <= 16'b0000_0000_0000_0000;
array[48337] <= 16'b0000_0000_0000_0000;
array[48338] <= 16'b0000_0000_0000_0000;
array[48339] <= 16'b0000_0000_0000_0000;
array[48340] <= 16'b0000_0000_0000_0000;
array[48341] <= 16'b0000_0000_0000_0000;
array[48342] <= 16'b0000_0000_0000_0000;
array[48343] <= 16'b0000_0000_0000_0000;
array[48344] <= 16'b0000_0000_0000_0000;
array[48345] <= 16'b0000_0000_0000_0000;
array[48346] <= 16'b0000_0000_0000_0000;
array[48347] <= 16'b0000_0000_0000_0000;
array[48348] <= 16'b0000_0000_0000_0000;
array[48349] <= 16'b0000_0000_0000_0000;
array[48350] <= 16'b0000_0000_0000_0000;
array[48351] <= 16'b0000_0000_0000_0000;
array[48352] <= 16'b0000_0000_0000_0000;
array[48353] <= 16'b0000_0000_0000_0000;
array[48354] <= 16'b0000_0000_0000_0000;
array[48355] <= 16'b0000_0000_0000_0000;
array[48356] <= 16'b0000_0000_0000_0000;
array[48357] <= 16'b0000_0000_0000_0000;
array[48358] <= 16'b0000_0000_0000_0000;
array[48359] <= 16'b0000_0000_0000_0000;
array[48360] <= 16'b0000_0000_0000_0000;
array[48361] <= 16'b0000_0000_0000_0000;
array[48362] <= 16'b0000_0000_0000_0000;
array[48363] <= 16'b0000_0000_0000_0000;
array[48364] <= 16'b0000_0000_0000_0000;
array[48365] <= 16'b0000_0000_0000_0000;
array[48366] <= 16'b0000_0000_0000_0000;
array[48367] <= 16'b0000_0000_0000_0000;
array[48368] <= 16'b0000_0000_0000_0000;
array[48369] <= 16'b0000_0000_0000_0000;
array[48370] <= 16'b0000_0000_0000_0000;
array[48371] <= 16'b0000_0000_0000_0000;
array[48372] <= 16'b0000_0000_0000_0000;
array[48373] <= 16'b0000_0000_0000_0000;
array[48374] <= 16'b0000_0000_0000_0000;
array[48375] <= 16'b0000_0000_0000_0000;
array[48376] <= 16'b0000_0000_0000_0000;
array[48377] <= 16'b0000_0000_0000_0000;
array[48378] <= 16'b0000_0000_0000_0000;
array[48379] <= 16'b0000_0000_0000_0000;
array[48380] <= 16'b0000_0000_0000_0000;
array[48381] <= 16'b0000_0000_0000_0000;
array[48382] <= 16'b0000_0000_0000_0000;
array[48383] <= 16'b0000_0000_0000_0000;
array[48384] <= 16'b0000_0000_0000_0000;
array[48385] <= 16'b0000_0000_0000_0000;
array[48386] <= 16'b0000_0000_0000_0000;
array[48387] <= 16'b0000_0000_0000_0000;
array[48388] <= 16'b0000_0000_0000_0000;
array[48389] <= 16'b0000_0000_0000_0000;
array[48390] <= 16'b0000_0000_0000_0000;
array[48391] <= 16'b0000_0000_0000_0000;
array[48392] <= 16'b0000_0000_0000_0000;
array[48393] <= 16'b0000_0000_0000_0000;
array[48394] <= 16'b0000_0000_0000_0000;
array[48395] <= 16'b0000_0000_0000_0000;
array[48396] <= 16'b0000_0000_0000_0000;
array[48397] <= 16'b0000_0000_0000_0000;
array[48398] <= 16'b0000_0000_0000_0000;
array[48399] <= 16'b0000_0000_0000_0000;
array[48400] <= 16'b0000_0000_0000_0000;
array[48401] <= 16'b0000_0000_0000_0000;
array[48402] <= 16'b0000_0000_0000_0000;
array[48403] <= 16'b0000_0000_0000_0000;
array[48404] <= 16'b0000_0000_0000_0000;
array[48405] <= 16'b0000_0000_0000_0000;
array[48406] <= 16'b0000_0000_0000_0000;
array[48407] <= 16'b0000_0000_0000_0000;
array[48408] <= 16'b0000_0000_0000_0000;
array[48409] <= 16'b0000_0000_0000_0000;
array[48410] <= 16'b0000_0000_0000_0000;
array[48411] <= 16'b0000_0000_0000_0000;
array[48412] <= 16'b0000_0000_0000_0000;
array[48413] <= 16'b0000_0000_0000_0000;
array[48414] <= 16'b0000_0000_0000_0000;
array[48415] <= 16'b0000_0000_0000_0000;
array[48416] <= 16'b0000_0000_0000_0000;
array[48417] <= 16'b0000_0000_0000_0000;
array[48418] <= 16'b0000_0000_0000_0000;
array[48419] <= 16'b0000_0000_0000_0000;
array[48420] <= 16'b0000_0000_0000_0000;
array[48421] <= 16'b0000_0000_0000_0000;
array[48422] <= 16'b0000_0000_0000_0000;
array[48423] <= 16'b0000_0000_0000_0000;
array[48424] <= 16'b0000_0000_0000_0000;
array[48425] <= 16'b0000_0000_0000_0000;
array[48426] <= 16'b0000_0000_0000_0000;
array[48427] <= 16'b0000_0000_0000_0000;
array[48428] <= 16'b0000_0000_0000_0000;
array[48429] <= 16'b0000_0000_0000_0000;
array[48430] <= 16'b0000_0000_0000_0000;
array[48431] <= 16'b0000_0000_0000_0000;
array[48432] <= 16'b0000_0000_0000_0000;
array[48433] <= 16'b0000_0000_0000_0000;
array[48434] <= 16'b0000_0000_0000_0000;
array[48435] <= 16'b0000_0000_0000_0000;
array[48436] <= 16'b0000_0000_0000_0000;
array[48437] <= 16'b0000_0000_0000_0000;
array[48438] <= 16'b0000_0000_0000_0000;
array[48439] <= 16'b0000_0000_0000_0000;
array[48440] <= 16'b0000_0000_0000_0000;
array[48441] <= 16'b0000_0000_0000_0000;
array[48442] <= 16'b0000_0000_0000_0000;
array[48443] <= 16'b0000_0000_0000_0000;
array[48444] <= 16'b0000_0000_0000_0000;
array[48445] <= 16'b0000_0000_0000_0000;
array[48446] <= 16'b0000_0000_0000_0000;
array[48447] <= 16'b0000_0000_0000_0000;
array[48448] <= 16'b0000_0000_0000_0000;
array[48449] <= 16'b0000_0000_0000_0000;
array[48450] <= 16'b0000_0000_0000_0000;
array[48451] <= 16'b0000_0000_0000_0000;
array[48452] <= 16'b0000_0000_0000_0000;
array[48453] <= 16'b0000_0000_0000_0000;
array[48454] <= 16'b0000_0000_0000_0000;
array[48455] <= 16'b0000_0000_0000_0000;
array[48456] <= 16'b0000_0000_0000_0000;
array[48457] <= 16'b0000_0000_0000_0000;
array[48458] <= 16'b0000_0000_0000_0000;
array[48459] <= 16'b0000_0000_0000_0000;
array[48460] <= 16'b0000_0000_0000_0000;
array[48461] <= 16'b0000_0000_0000_0000;
array[48462] <= 16'b0000_0000_0000_0000;
array[48463] <= 16'b0000_0000_0000_0000;
array[48464] <= 16'b0000_0000_0000_0000;
array[48465] <= 16'b0000_0000_0000_0000;
array[48466] <= 16'b0000_0000_0000_0000;
array[48467] <= 16'b0000_0000_0000_0000;
array[48468] <= 16'b0000_0000_0000_0000;
array[48469] <= 16'b0000_0000_0000_0000;
array[48470] <= 16'b0000_0000_0000_0000;
array[48471] <= 16'b0000_0000_0000_0000;
array[48472] <= 16'b0000_0000_0000_0000;
array[48473] <= 16'b0000_0000_0000_0000;
array[48474] <= 16'b0000_0000_0000_0000;
array[48475] <= 16'b0000_0000_0000_0000;
array[48476] <= 16'b0000_0000_0000_0000;
array[48477] <= 16'b0000_0000_0000_0000;
array[48478] <= 16'b0000_0000_0000_0000;
array[48479] <= 16'b0000_0000_0000_0000;
array[48480] <= 16'b0000_0000_0000_0000;
array[48481] <= 16'b0000_0000_0000_0000;
array[48482] <= 16'b0000_0000_0000_0000;
array[48483] <= 16'b0000_0000_0000_0000;
array[48484] <= 16'b0000_0000_0000_0000;
array[48485] <= 16'b0000_0000_0000_0000;
array[48486] <= 16'b0000_0000_0000_0000;
array[48487] <= 16'b0000_0000_0000_0000;
array[48488] <= 16'b0000_0000_0000_0000;
array[48489] <= 16'b0000_0000_0000_0000;
array[48490] <= 16'b0000_0000_0000_0000;
array[48491] <= 16'b0000_0000_0000_0000;
array[48492] <= 16'b0000_0000_0000_0000;
array[48493] <= 16'b0000_0000_0000_0000;
array[48494] <= 16'b0000_0000_0000_0000;
array[48495] <= 16'b0000_0000_0000_0000;
array[48496] <= 16'b0000_0000_0000_0000;
array[48497] <= 16'b0000_0000_0000_0000;
array[48498] <= 16'b0000_0000_0000_0000;
array[48499] <= 16'b0000_0000_0000_0000;
array[48500] <= 16'b0000_0000_0000_0000;
array[48501] <= 16'b0000_0000_0000_0000;
array[48502] <= 16'b0000_0000_0000_0000;
array[48503] <= 16'b0000_0000_0000_0000;
array[48504] <= 16'b0000_0000_0000_0000;
array[48505] <= 16'b0000_0000_0000_0000;
array[48506] <= 16'b0000_0000_0000_0000;
array[48507] <= 16'b0000_0000_0000_0000;
array[48508] <= 16'b0000_0000_0000_0000;
array[48509] <= 16'b0000_0000_0000_0000;
array[48510] <= 16'b0000_0000_0000_0000;
array[48511] <= 16'b0000_0000_0000_0000;
array[48512] <= 16'b0000_0000_0000_0000;
array[48513] <= 16'b0000_0000_0000_0000;
array[48514] <= 16'b0000_0000_0000_0000;
array[48515] <= 16'b0000_0000_0000_0000;
array[48516] <= 16'b0000_0000_0000_0000;
array[48517] <= 16'b0000_0000_0000_0000;
array[48518] <= 16'b0000_0000_0000_0000;
array[48519] <= 16'b0000_0000_0000_0000;
array[48520] <= 16'b0000_0000_0000_0000;
array[48521] <= 16'b0000_0000_0000_0000;
array[48522] <= 16'b0000_0000_0000_0000;
array[48523] <= 16'b0000_0000_0000_0000;
array[48524] <= 16'b0000_0000_0000_0000;
array[48525] <= 16'b0000_0000_0000_0000;
array[48526] <= 16'b0000_0000_0000_0000;
array[48527] <= 16'b0000_0000_0000_0000;
array[48528] <= 16'b0000_0000_0000_0000;
array[48529] <= 16'b0000_0000_0000_0000;
array[48530] <= 16'b0000_0000_0000_0000;
array[48531] <= 16'b0000_0000_0000_0000;
array[48532] <= 16'b0000_0000_0000_0000;
array[48533] <= 16'b0000_0000_0000_0000;
array[48534] <= 16'b0000_0000_0000_0000;
array[48535] <= 16'b0000_0000_0000_0000;
array[48536] <= 16'b0000_0000_0000_0000;
array[48537] <= 16'b0000_0000_0000_0000;
array[48538] <= 16'b0000_0000_0000_0000;
array[48539] <= 16'b0000_0000_0000_0000;
array[48540] <= 16'b0000_0000_0000_0000;
array[48541] <= 16'b0000_0000_0000_0000;
array[48542] <= 16'b0000_0000_0000_0000;
array[48543] <= 16'b0000_0000_0000_0000;
array[48544] <= 16'b0000_0000_0000_0000;
array[48545] <= 16'b0000_0000_0000_0000;
array[48546] <= 16'b0000_0000_0000_0000;
array[48547] <= 16'b0000_0000_0000_0000;
array[48548] <= 16'b0000_0000_0000_0000;
array[48549] <= 16'b0000_0000_0000_0000;
array[48550] <= 16'b0000_0000_0000_0000;
array[48551] <= 16'b0000_0000_0000_0000;
array[48552] <= 16'b0000_0000_0000_0000;
array[48553] <= 16'b0000_0000_0000_0000;
array[48554] <= 16'b0000_0000_0000_0000;
array[48555] <= 16'b0000_0000_0000_0000;
array[48556] <= 16'b0000_0000_0000_0000;
array[48557] <= 16'b0000_0000_0000_0000;
array[48558] <= 16'b0000_0000_0000_0000;
array[48559] <= 16'b0000_0000_0000_0000;
array[48560] <= 16'b0000_0000_0000_0000;
array[48561] <= 16'b0000_0000_0000_0000;
array[48562] <= 16'b0000_0000_0000_0000;
array[48563] <= 16'b0000_0000_0000_0000;
array[48564] <= 16'b0000_0000_0000_0000;
array[48565] <= 16'b0000_0000_0000_0000;
array[48566] <= 16'b0000_0000_0000_0000;
array[48567] <= 16'b0000_0000_0000_0000;
array[48568] <= 16'b0000_0000_0000_0000;
array[48569] <= 16'b0000_0000_0000_0000;
array[48570] <= 16'b0000_0000_0000_0000;
array[48571] <= 16'b0000_0000_0000_0000;
array[48572] <= 16'b0000_0000_0000_0000;
array[48573] <= 16'b0000_0000_0000_0000;
array[48574] <= 16'b0000_0000_0000_0000;
array[48575] <= 16'b0000_0000_0000_0000;
array[48576] <= 16'b0000_0000_0000_0000;
array[48577] <= 16'b0000_0000_0000_0000;
array[48578] <= 16'b0000_0000_0000_0000;
array[48579] <= 16'b0000_0000_0000_0000;
array[48580] <= 16'b0000_0000_0000_0000;
array[48581] <= 16'b0000_0000_0000_0000;
array[48582] <= 16'b0000_0000_0000_0000;
array[48583] <= 16'b0000_0000_0000_0000;
array[48584] <= 16'b0000_0000_0000_0000;
array[48585] <= 16'b0000_0000_0000_0000;
array[48586] <= 16'b0000_0000_0000_0000;
array[48587] <= 16'b0000_0000_0000_0000;
array[48588] <= 16'b0000_0000_0000_0000;
array[48589] <= 16'b0000_0000_0000_0000;
array[48590] <= 16'b0000_0000_0000_0000;
array[48591] <= 16'b0000_0000_0000_0000;
array[48592] <= 16'b0000_0000_0000_0000;
array[48593] <= 16'b0000_0000_0000_0000;
array[48594] <= 16'b0000_0000_0000_0000;
array[48595] <= 16'b0000_0000_0000_0000;
array[48596] <= 16'b0000_0000_0000_0000;
array[48597] <= 16'b0000_0000_0000_0000;
array[48598] <= 16'b0000_0000_0000_0000;
array[48599] <= 16'b0000_0000_0000_0000;
array[48600] <= 16'b0000_0000_0000_0000;
array[48601] <= 16'b0000_0000_0000_0000;
array[48602] <= 16'b0000_0000_0000_0000;
array[48603] <= 16'b0000_0000_0000_0000;
array[48604] <= 16'b0000_0000_0000_0000;
array[48605] <= 16'b0000_0000_0000_0000;
array[48606] <= 16'b0000_0000_0000_0000;
array[48607] <= 16'b0000_0000_0000_0000;
array[48608] <= 16'b0000_0000_0000_0000;
array[48609] <= 16'b0000_0000_0000_0000;
array[48610] <= 16'b0000_0000_0000_0000;
array[48611] <= 16'b0000_0000_0000_0000;
array[48612] <= 16'b0000_0000_0000_0000;
array[48613] <= 16'b0000_0000_0000_0000;
array[48614] <= 16'b0000_0000_0000_0000;
array[48615] <= 16'b0000_0000_0000_0000;
array[48616] <= 16'b0000_0000_0000_0000;
array[48617] <= 16'b0000_0000_0000_0000;
array[48618] <= 16'b0000_0000_0000_0000;
array[48619] <= 16'b0000_0000_0000_0000;
array[48620] <= 16'b0000_0000_0000_0000;
array[48621] <= 16'b0000_0000_0000_0000;
array[48622] <= 16'b0000_0000_0000_0000;
array[48623] <= 16'b0000_0000_0000_0000;
array[48624] <= 16'b0000_0000_0000_0000;
array[48625] <= 16'b0000_0000_0000_0000;
array[48626] <= 16'b0000_0000_0000_0000;
array[48627] <= 16'b0000_0000_0000_0000;
array[48628] <= 16'b0000_0000_0000_0000;
array[48629] <= 16'b0000_0000_0000_0000;
array[48630] <= 16'b0000_0000_0000_0000;
array[48631] <= 16'b0000_0000_0000_0000;
array[48632] <= 16'b0000_0000_0000_0000;
array[48633] <= 16'b0000_0000_0000_0000;
array[48634] <= 16'b0000_0000_0000_0000;
array[48635] <= 16'b0000_0000_0000_0000;
array[48636] <= 16'b0000_0000_0000_0000;
array[48637] <= 16'b0000_0000_0000_0000;
array[48638] <= 16'b0000_0000_0000_0000;
array[48639] <= 16'b0000_0000_0000_0000;
array[48640] <= 16'b0000_0000_0000_0000;
array[48641] <= 16'b0000_0000_0000_0000;
array[48642] <= 16'b0000_0000_0000_0000;
array[48643] <= 16'b0000_0000_0000_0000;
array[48644] <= 16'b0000_0000_0000_0000;
array[48645] <= 16'b0000_0000_0000_0000;
array[48646] <= 16'b0000_0000_0000_0000;
array[48647] <= 16'b0000_0000_0000_0000;
array[48648] <= 16'b0000_0000_0000_0000;
array[48649] <= 16'b0000_0000_0000_0000;
array[48650] <= 16'b0000_0000_0000_0000;
array[48651] <= 16'b0000_0000_0000_0000;
array[48652] <= 16'b0000_0000_0000_0000;
array[48653] <= 16'b0000_0000_0000_0000;
array[48654] <= 16'b0000_0000_0000_0000;
array[48655] <= 16'b0000_0000_0000_0000;
array[48656] <= 16'b0000_0000_0000_0000;
array[48657] <= 16'b0000_0000_0000_0000;
array[48658] <= 16'b0000_0000_0000_0000;
array[48659] <= 16'b0000_0000_0000_0000;
array[48660] <= 16'b0000_0000_0000_0000;
array[48661] <= 16'b0000_0000_0000_0000;
array[48662] <= 16'b0000_0000_0000_0000;
array[48663] <= 16'b0000_0000_0000_0000;
array[48664] <= 16'b0000_0000_0000_0000;
array[48665] <= 16'b0000_0000_0000_0000;
array[48666] <= 16'b0000_0000_0000_0000;
array[48667] <= 16'b0000_0000_0000_0000;
array[48668] <= 16'b0000_0000_0000_0000;
array[48669] <= 16'b0000_0000_0000_0000;
array[48670] <= 16'b0000_0000_0000_0000;
array[48671] <= 16'b0000_0000_0000_0000;
array[48672] <= 16'b0000_0000_0000_0000;
array[48673] <= 16'b0000_0000_0000_0000;
array[48674] <= 16'b0000_0000_0000_0000;
array[48675] <= 16'b0000_0000_0000_0000;
array[48676] <= 16'b0000_0000_0000_0000;
array[48677] <= 16'b0000_0000_0000_0000;
array[48678] <= 16'b0000_0000_0000_0000;
array[48679] <= 16'b0000_0000_0000_0000;
array[48680] <= 16'b0000_0000_0000_0000;
array[48681] <= 16'b0000_0000_0000_0000;
array[48682] <= 16'b0000_0000_0000_0000;
array[48683] <= 16'b0000_0000_0000_0000;
array[48684] <= 16'b0000_0000_0000_0000;
array[48685] <= 16'b0000_0000_0000_0000;
array[48686] <= 16'b0000_0000_0000_0000;
array[48687] <= 16'b0000_0000_0000_0000;
array[48688] <= 16'b0000_0000_0000_0000;
array[48689] <= 16'b0000_0000_0000_0000;
array[48690] <= 16'b0000_0000_0000_0000;
array[48691] <= 16'b0000_0000_0000_0000;
array[48692] <= 16'b0000_0000_0000_0000;
array[48693] <= 16'b0000_0000_0000_0000;
array[48694] <= 16'b0000_0000_0000_0000;
array[48695] <= 16'b0000_0000_0000_0000;
array[48696] <= 16'b0000_0000_0000_0000;
array[48697] <= 16'b0000_0000_0000_0000;
array[48698] <= 16'b0000_0000_0000_0000;
array[48699] <= 16'b0000_0000_0000_0000;
array[48700] <= 16'b0000_0000_0000_0000;
array[48701] <= 16'b0000_0000_0000_0000;
array[48702] <= 16'b0000_0000_0000_0000;
array[48703] <= 16'b0000_0000_0000_0000;
array[48704] <= 16'b0000_0000_0000_0000;
array[48705] <= 16'b0000_0000_0000_0000;
array[48706] <= 16'b0000_0000_0000_0000;
array[48707] <= 16'b0000_0000_0000_0000;
array[48708] <= 16'b0000_0000_0000_0000;
array[48709] <= 16'b0000_0000_0000_0000;
array[48710] <= 16'b0000_0000_0000_0000;
array[48711] <= 16'b0000_0000_0000_0000;
array[48712] <= 16'b0000_0000_0000_0000;
array[48713] <= 16'b0000_0000_0000_0000;
array[48714] <= 16'b0000_0000_0000_0000;
array[48715] <= 16'b0000_0000_0000_0000;
array[48716] <= 16'b0000_0000_0000_0000;
array[48717] <= 16'b0000_0000_0000_0000;
array[48718] <= 16'b0000_0000_0000_0000;
array[48719] <= 16'b0000_0000_0000_0000;
array[48720] <= 16'b0000_0000_0000_0000;
array[48721] <= 16'b0000_0000_0000_0000;
array[48722] <= 16'b0000_0000_0000_0000;
array[48723] <= 16'b0000_0000_0000_0000;
array[48724] <= 16'b0000_0000_0000_0000;
array[48725] <= 16'b0000_0000_0000_0000;
array[48726] <= 16'b0000_0000_0000_0000;
array[48727] <= 16'b0000_0000_0000_0000;
array[48728] <= 16'b0000_0000_0000_0000;
array[48729] <= 16'b0000_0000_0000_0000;
array[48730] <= 16'b0000_0000_0000_0000;
array[48731] <= 16'b0000_0000_0000_0000;
array[48732] <= 16'b0000_0000_0000_0000;
array[48733] <= 16'b0000_0000_0000_0000;
array[48734] <= 16'b0000_0000_0000_0000;
array[48735] <= 16'b0000_0000_0000_0000;
array[48736] <= 16'b0000_0000_0000_0000;
array[48737] <= 16'b0000_0000_0000_0000;
array[48738] <= 16'b0000_0000_0000_0000;
array[48739] <= 16'b0000_0000_0000_0000;
array[48740] <= 16'b0000_0000_0000_0000;
array[48741] <= 16'b0000_0000_0000_0000;
array[48742] <= 16'b0000_0000_0000_0000;
array[48743] <= 16'b0000_0000_0000_0000;
array[48744] <= 16'b0000_0000_0000_0000;
array[48745] <= 16'b0000_0000_0000_0000;
array[48746] <= 16'b0000_0000_0000_0000;
array[48747] <= 16'b0000_0000_0000_0000;
array[48748] <= 16'b0000_0000_0000_0000;
array[48749] <= 16'b0000_0000_0000_0000;
array[48750] <= 16'b0000_0000_0000_0000;
array[48751] <= 16'b0000_0000_0000_0000;
array[48752] <= 16'b0000_0000_0000_0000;
array[48753] <= 16'b0000_0000_0000_0000;
array[48754] <= 16'b0000_0000_0000_0000;
array[48755] <= 16'b0000_0000_0000_0000;
array[48756] <= 16'b0000_0000_0000_0000;
array[48757] <= 16'b0000_0000_0000_0000;
array[48758] <= 16'b0000_0000_0000_0000;
array[48759] <= 16'b0000_0000_0000_0000;
array[48760] <= 16'b0000_0000_0000_0000;
array[48761] <= 16'b0000_0000_0000_0000;
array[48762] <= 16'b0000_0000_0000_0000;
array[48763] <= 16'b0000_0000_0000_0000;
array[48764] <= 16'b0000_0000_0000_0000;
array[48765] <= 16'b0000_0000_0000_0000;
array[48766] <= 16'b0000_0000_0000_0000;
array[48767] <= 16'b0000_0000_0000_0000;
array[48768] <= 16'b0000_0000_0000_0000;
array[48769] <= 16'b0000_0000_0000_0000;
array[48770] <= 16'b0000_0000_0000_0000;
array[48771] <= 16'b0000_0000_0000_0000;
array[48772] <= 16'b0000_0000_0000_0000;
array[48773] <= 16'b0000_0000_0000_0000;
array[48774] <= 16'b0000_0000_0000_0000;
array[48775] <= 16'b0000_0000_0000_0000;
array[48776] <= 16'b0000_0000_0000_0000;
array[48777] <= 16'b0000_0000_0000_0000;
array[48778] <= 16'b0000_0000_0000_0000;
array[48779] <= 16'b0000_0000_0000_0000;
array[48780] <= 16'b0000_0000_0000_0000;
array[48781] <= 16'b0000_0000_0000_0000;
array[48782] <= 16'b0000_0000_0000_0000;
array[48783] <= 16'b0000_0000_0000_0000;
array[48784] <= 16'b0000_0000_0000_0000;
array[48785] <= 16'b0000_0000_0000_0000;
array[48786] <= 16'b0000_0000_0000_0000;
array[48787] <= 16'b0000_0000_0000_0000;
array[48788] <= 16'b0000_0000_0000_0000;
array[48789] <= 16'b0000_0000_0000_0000;
array[48790] <= 16'b0000_0000_0000_0000;
array[48791] <= 16'b0000_0000_0000_0000;
array[48792] <= 16'b0000_0000_0000_0000;
array[48793] <= 16'b0000_0000_0000_0000;
array[48794] <= 16'b0000_0000_0000_0000;
array[48795] <= 16'b0000_0000_0000_0000;
array[48796] <= 16'b0000_0000_0000_0000;
array[48797] <= 16'b0000_0000_0000_0000;
array[48798] <= 16'b0000_0000_0000_0000;
array[48799] <= 16'b0000_0000_0000_0000;
array[48800] <= 16'b0000_0000_0000_0000;
array[48801] <= 16'b0000_0000_0000_0000;
array[48802] <= 16'b0000_0000_0000_0000;
array[48803] <= 16'b0000_0000_0000_0000;
array[48804] <= 16'b0000_0000_0000_0000;
array[48805] <= 16'b0000_0000_0000_0000;
array[48806] <= 16'b0000_0000_0000_0000;
array[48807] <= 16'b0000_0000_0000_0000;
array[48808] <= 16'b0000_0000_0000_0000;
array[48809] <= 16'b0000_0000_0000_0000;
array[48810] <= 16'b0000_0000_0000_0000;
array[48811] <= 16'b0000_0000_0000_0000;
array[48812] <= 16'b0000_0000_0000_0000;
array[48813] <= 16'b0000_0000_0000_0000;
array[48814] <= 16'b0000_0000_0000_0000;
array[48815] <= 16'b0000_0000_0000_0000;
array[48816] <= 16'b0000_0000_0000_0000;
array[48817] <= 16'b0000_0000_0000_0000;
array[48818] <= 16'b0000_0000_0000_0000;
array[48819] <= 16'b0000_0000_0000_0000;
array[48820] <= 16'b0000_0000_0000_0000;
array[48821] <= 16'b0000_0000_0000_0000;
array[48822] <= 16'b0000_0000_0000_0000;
array[48823] <= 16'b0000_0000_0000_0000;
array[48824] <= 16'b0000_0000_0000_0000;
array[48825] <= 16'b0000_0000_0000_0000;
array[48826] <= 16'b0000_0000_0000_0000;
array[48827] <= 16'b0000_0000_0000_0000;
array[48828] <= 16'b0000_0000_0000_0000;
array[48829] <= 16'b0000_0000_0000_0000;
array[48830] <= 16'b0000_0000_0000_0000;
array[48831] <= 16'b0000_0000_0000_0000;
array[48832] <= 16'b0000_0000_0000_0000;
array[48833] <= 16'b0000_0000_0000_0000;
array[48834] <= 16'b0000_0000_0000_0000;
array[48835] <= 16'b0000_0000_0000_0000;
array[48836] <= 16'b0000_0000_0000_0000;
array[48837] <= 16'b0000_0000_0000_0000;
array[48838] <= 16'b0000_0000_0000_0000;
array[48839] <= 16'b0000_0000_0000_0000;
array[48840] <= 16'b0000_0000_0000_0000;
array[48841] <= 16'b0000_0000_0000_0000;
array[48842] <= 16'b0000_0000_0000_0000;
array[48843] <= 16'b0000_0000_0000_0000;
array[48844] <= 16'b0000_0000_0000_0000;
array[48845] <= 16'b0000_0000_0000_0000;
array[48846] <= 16'b0000_0000_0000_0000;
array[48847] <= 16'b0000_0000_0000_0000;
array[48848] <= 16'b0000_0000_0000_0000;
array[48849] <= 16'b0000_0000_0000_0000;
array[48850] <= 16'b0000_0000_0000_0000;
array[48851] <= 16'b0000_0000_0000_0000;
array[48852] <= 16'b0000_0000_0000_0000;
array[48853] <= 16'b0000_0000_0000_0000;
array[48854] <= 16'b0000_0000_0000_0000;
array[48855] <= 16'b0000_0000_0000_0000;
array[48856] <= 16'b0000_0000_0000_0000;
array[48857] <= 16'b0000_0000_0000_0000;
array[48858] <= 16'b0000_0000_0000_0000;
array[48859] <= 16'b0000_0000_0000_0000;
array[48860] <= 16'b0000_0000_0000_0000;
array[48861] <= 16'b0000_0000_0000_0000;
array[48862] <= 16'b0000_0000_0000_0000;
array[48863] <= 16'b0000_0000_0000_0000;
array[48864] <= 16'b0000_0000_0000_0000;
array[48865] <= 16'b0000_0000_0000_0000;
array[48866] <= 16'b0000_0000_0000_0000;
array[48867] <= 16'b0000_0000_0000_0000;
array[48868] <= 16'b0000_0000_0000_0000;
array[48869] <= 16'b0000_0000_0000_0000;
array[48870] <= 16'b0000_0000_0000_0000;
array[48871] <= 16'b0000_0000_0000_0000;
array[48872] <= 16'b0000_0000_0000_0000;
array[48873] <= 16'b0000_0000_0000_0000;
array[48874] <= 16'b0000_0000_0000_0000;
array[48875] <= 16'b0000_0000_0000_0000;
array[48876] <= 16'b0000_0000_0000_0000;
array[48877] <= 16'b0000_0000_0000_0000;
array[48878] <= 16'b0000_0000_0000_0000;
array[48879] <= 16'b0000_0000_0000_0000;
array[48880] <= 16'b0000_0000_0000_0000;
array[48881] <= 16'b0000_0000_0000_0000;
array[48882] <= 16'b0000_0000_0000_0000;
array[48883] <= 16'b0000_0000_0000_0000;
array[48884] <= 16'b0000_0000_0000_0000;
array[48885] <= 16'b0000_0000_0000_0000;
array[48886] <= 16'b0000_0000_0000_0000;
array[48887] <= 16'b0000_0000_0000_0000;
array[48888] <= 16'b0000_0000_0000_0000;
array[48889] <= 16'b0000_0000_0000_0000;
array[48890] <= 16'b0000_0000_0000_0000;
array[48891] <= 16'b0000_0000_0000_0000;
array[48892] <= 16'b0000_0000_0000_0000;
array[48893] <= 16'b0000_0000_0000_0000;
array[48894] <= 16'b0000_0000_0000_0000;
array[48895] <= 16'b0000_0000_0000_0000;
array[48896] <= 16'b0000_0000_0000_0000;
array[48897] <= 16'b0000_0000_0000_0000;
array[48898] <= 16'b0000_0000_0000_0000;
array[48899] <= 16'b0000_0000_0000_0000;
array[48900] <= 16'b0000_0000_0000_0000;
array[48901] <= 16'b0000_0000_0000_0000;
array[48902] <= 16'b0000_0000_0000_0000;
array[48903] <= 16'b0000_0000_0000_0000;
array[48904] <= 16'b0000_0000_0000_0000;
array[48905] <= 16'b0000_0000_0000_0000;
array[48906] <= 16'b0000_0000_0000_0000;
array[48907] <= 16'b0000_0000_0000_0000;
array[48908] <= 16'b0000_0000_0000_0000;
array[48909] <= 16'b0000_0000_0000_0000;
array[48910] <= 16'b0000_0000_0000_0000;
array[48911] <= 16'b0000_0000_0000_0000;
array[48912] <= 16'b0000_0000_0000_0000;
array[48913] <= 16'b0000_0000_0000_0000;
array[48914] <= 16'b0000_0000_0000_0000;
array[48915] <= 16'b0000_0000_0000_0000;
array[48916] <= 16'b0000_0000_0000_0000;
array[48917] <= 16'b0000_0000_0000_0000;
array[48918] <= 16'b0000_0000_0000_0000;
array[48919] <= 16'b0000_0000_0000_0000;
array[48920] <= 16'b0000_0000_0000_0000;
array[48921] <= 16'b0000_0000_0000_0000;
array[48922] <= 16'b0000_0000_0000_0000;
array[48923] <= 16'b0000_0000_0000_0000;
array[48924] <= 16'b0000_0000_0000_0000;
array[48925] <= 16'b0000_0000_0000_0000;
array[48926] <= 16'b0000_0000_0000_0000;
array[48927] <= 16'b0000_0000_0000_0000;
array[48928] <= 16'b0000_0000_0000_0000;
array[48929] <= 16'b0000_0000_0000_0000;
array[48930] <= 16'b0000_0000_0000_0000;
array[48931] <= 16'b0000_0000_0000_0000;
array[48932] <= 16'b0000_0000_0000_0000;
array[48933] <= 16'b0000_0000_0000_0000;
array[48934] <= 16'b0000_0000_0000_0000;
array[48935] <= 16'b0000_0000_0000_0000;
array[48936] <= 16'b0000_0000_0000_0000;
array[48937] <= 16'b0000_0000_0000_0000;
array[48938] <= 16'b0000_0000_0000_0000;
array[48939] <= 16'b0000_0000_0000_0000;
array[48940] <= 16'b0000_0000_0000_0000;
array[48941] <= 16'b0000_0000_0000_0000;
array[48942] <= 16'b0000_0000_0000_0000;
array[48943] <= 16'b0000_0000_0000_0000;
array[48944] <= 16'b0000_0000_0000_0000;
array[48945] <= 16'b0000_0000_0000_0000;
array[48946] <= 16'b0000_0000_0000_0000;
array[48947] <= 16'b0000_0000_0000_0000;
array[48948] <= 16'b0000_0000_0000_0000;
array[48949] <= 16'b0000_0000_0000_0000;
array[48950] <= 16'b0000_0000_0000_0000;
array[48951] <= 16'b0000_0000_0000_0000;
array[48952] <= 16'b0000_0000_0000_0000;
array[48953] <= 16'b0000_0000_0000_0000;
array[48954] <= 16'b0000_0000_0000_0000;
array[48955] <= 16'b0000_0000_0000_0000;
array[48956] <= 16'b0000_0000_0000_0000;
array[48957] <= 16'b0000_0000_0000_0000;
array[48958] <= 16'b0000_0000_0000_0000;
array[48959] <= 16'b0000_0000_0000_0000;
array[48960] <= 16'b0000_0000_0000_0000;
array[48961] <= 16'b0000_0000_0000_0000;
array[48962] <= 16'b0000_0000_0000_0000;
array[48963] <= 16'b0000_0000_0000_0000;
array[48964] <= 16'b0000_0000_0000_0000;
array[48965] <= 16'b0000_0000_0000_0000;
array[48966] <= 16'b0000_0000_0000_0000;
array[48967] <= 16'b0000_0000_0000_0000;
array[48968] <= 16'b0000_0000_0000_0000;
array[48969] <= 16'b0000_0000_0000_0000;
array[48970] <= 16'b0000_0000_0000_0000;
array[48971] <= 16'b0000_0000_0000_0000;
array[48972] <= 16'b0000_0000_0000_0000;
array[48973] <= 16'b0000_0000_0000_0000;
array[48974] <= 16'b0000_0000_0000_0000;
array[48975] <= 16'b0000_0000_0000_0000;
array[48976] <= 16'b0000_0000_0000_0000;
array[48977] <= 16'b0000_0000_0000_0000;
array[48978] <= 16'b0000_0000_0000_0000;
array[48979] <= 16'b0000_0000_0000_0000;
array[48980] <= 16'b0000_0000_0000_0000;
array[48981] <= 16'b0000_0000_0000_0000;
array[48982] <= 16'b0000_0000_0000_0000;
array[48983] <= 16'b0000_0000_0000_0000;
array[48984] <= 16'b0000_0000_0000_0000;
array[48985] <= 16'b0000_0000_0000_0000;
array[48986] <= 16'b0000_0000_0000_0000;
array[48987] <= 16'b0000_0000_0000_0000;
array[48988] <= 16'b0000_0000_0000_0000;
array[48989] <= 16'b0000_0000_0000_0000;
array[48990] <= 16'b0000_0000_0000_0000;
array[48991] <= 16'b0000_0000_0000_0000;
array[48992] <= 16'b0000_0000_0000_0000;
array[48993] <= 16'b0000_0000_0000_0000;
array[48994] <= 16'b0000_0000_0000_0000;
array[48995] <= 16'b0000_0000_0000_0000;
array[48996] <= 16'b0000_0000_0000_0000;
array[48997] <= 16'b0000_0000_0000_0000;
array[48998] <= 16'b0000_0000_0000_0000;
array[48999] <= 16'b0000_0000_0000_0000;
array[49000] <= 16'b0000_0000_0000_0000;
array[49001] <= 16'b0000_0000_0000_0000;
array[49002] <= 16'b0000_0000_0000_0000;
array[49003] <= 16'b0000_0000_0000_0000;
array[49004] <= 16'b0000_0000_0000_0000;
array[49005] <= 16'b0000_0000_0000_0000;
array[49006] <= 16'b0000_0000_0000_0000;
array[49007] <= 16'b0000_0000_0000_0000;
array[49008] <= 16'b0000_0000_0000_0000;
array[49009] <= 16'b0000_0000_0000_0000;
array[49010] <= 16'b0000_0000_0000_0000;
array[49011] <= 16'b0000_0000_0000_0000;
array[49012] <= 16'b0000_0000_0000_0000;
array[49013] <= 16'b0000_0000_0000_0000;
array[49014] <= 16'b0000_0000_0000_0000;
array[49015] <= 16'b0000_0000_0000_0000;
array[49016] <= 16'b0000_0000_0000_0000;
array[49017] <= 16'b0000_0000_0000_0000;
array[49018] <= 16'b0000_0000_0000_0000;
array[49019] <= 16'b0000_0000_0000_0000;
array[49020] <= 16'b0000_0000_0000_0000;
array[49021] <= 16'b0000_0000_0000_0000;
array[49022] <= 16'b0000_0000_0000_0000;
array[49023] <= 16'b0000_0000_0000_0000;
array[49024] <= 16'b0000_0000_0000_0000;
array[49025] <= 16'b0000_0000_0000_0000;
array[49026] <= 16'b0000_0000_0000_0000;
array[49027] <= 16'b0000_0000_0000_0000;
array[49028] <= 16'b0000_0000_0000_0000;
array[49029] <= 16'b0000_0000_0000_0000;
array[49030] <= 16'b0000_0000_0000_0000;
array[49031] <= 16'b0000_0000_0000_0000;
array[49032] <= 16'b0000_0000_0000_0000;
array[49033] <= 16'b0000_0000_0000_0000;
array[49034] <= 16'b0000_0000_0000_0000;
array[49035] <= 16'b0000_0000_0000_0000;
array[49036] <= 16'b0000_0000_0000_0000;
array[49037] <= 16'b0000_0000_0000_0000;
array[49038] <= 16'b0000_0000_0000_0000;
array[49039] <= 16'b0000_0000_0000_0000;
array[49040] <= 16'b0000_0000_0000_0000;
array[49041] <= 16'b0000_0000_0000_0000;
array[49042] <= 16'b0000_0000_0000_0000;
array[49043] <= 16'b0000_0000_0000_0000;
array[49044] <= 16'b0000_0000_0000_0000;
array[49045] <= 16'b0000_0000_0000_0000;
array[49046] <= 16'b0000_0000_0000_0000;
array[49047] <= 16'b0000_0000_0000_0000;
array[49048] <= 16'b0000_0000_0000_0000;
array[49049] <= 16'b0000_0000_0000_0000;
array[49050] <= 16'b0000_0000_0000_0000;
array[49051] <= 16'b0000_0000_0000_0000;
array[49052] <= 16'b0000_0000_0000_0000;
array[49053] <= 16'b0000_0000_0000_0000;
array[49054] <= 16'b0000_0000_0000_0000;
array[49055] <= 16'b0000_0000_0000_0000;
array[49056] <= 16'b0000_0000_0000_0000;
array[49057] <= 16'b0000_0000_0000_0000;
array[49058] <= 16'b0000_0000_0000_0000;
array[49059] <= 16'b0000_0000_0000_0000;
array[49060] <= 16'b0000_0000_0000_0000;
array[49061] <= 16'b0000_0000_0000_0000;
array[49062] <= 16'b0000_0000_0000_0000;
array[49063] <= 16'b0000_0000_0000_0000;
array[49064] <= 16'b0000_0000_0000_0000;
array[49065] <= 16'b0000_0000_0000_0000;
array[49066] <= 16'b0000_0000_0000_0000;
array[49067] <= 16'b0000_0000_0000_0000;
array[49068] <= 16'b0000_0000_0000_0000;
array[49069] <= 16'b0000_0000_0000_0000;
array[49070] <= 16'b0000_0000_0000_0000;
array[49071] <= 16'b0000_0000_0000_0000;
array[49072] <= 16'b0000_0000_0000_0000;
array[49073] <= 16'b0000_0000_0000_0000;
array[49074] <= 16'b0000_0000_0000_0000;
array[49075] <= 16'b0000_0000_0000_0000;
array[49076] <= 16'b0000_0000_0000_0000;
array[49077] <= 16'b0000_0000_0000_0000;
array[49078] <= 16'b0000_0000_0000_0000;
array[49079] <= 16'b0000_0000_0000_0000;
array[49080] <= 16'b0000_0000_0000_0000;
array[49081] <= 16'b0000_0000_0000_0000;
array[49082] <= 16'b0000_0000_0000_0000;
array[49083] <= 16'b0000_0000_0000_0000;
array[49084] <= 16'b0000_0000_0000_0000;
array[49085] <= 16'b0000_0000_0000_0000;
array[49086] <= 16'b0000_0000_0000_0000;
array[49087] <= 16'b0000_0000_0000_0000;
array[49088] <= 16'b0000_0000_0000_0000;
array[49089] <= 16'b0000_0000_0000_0000;
array[49090] <= 16'b0000_0000_0000_0000;
array[49091] <= 16'b0000_0000_0000_0000;
array[49092] <= 16'b0000_0000_0000_0000;
array[49093] <= 16'b0000_0000_0000_0000;
array[49094] <= 16'b0000_0000_0000_0000;
array[49095] <= 16'b0000_0000_0000_0000;
array[49096] <= 16'b0000_0000_0000_0000;
array[49097] <= 16'b0000_0000_0000_0000;
array[49098] <= 16'b0000_0000_0000_0000;
array[49099] <= 16'b0000_0000_0000_0000;
array[49100] <= 16'b0000_0000_0000_0000;
array[49101] <= 16'b0000_0000_0000_0000;
array[49102] <= 16'b0000_0000_0000_0000;
array[49103] <= 16'b0000_0000_0000_0000;
array[49104] <= 16'b0000_0000_0000_0000;
array[49105] <= 16'b0000_0000_0000_0000;
array[49106] <= 16'b0000_0000_0000_0000;
array[49107] <= 16'b0000_0000_0000_0000;
array[49108] <= 16'b0000_0000_0000_0000;
array[49109] <= 16'b0000_0000_0000_0000;
array[49110] <= 16'b0000_0000_0000_0000;
array[49111] <= 16'b0000_0000_0000_0000;
array[49112] <= 16'b0000_0000_0000_0000;
array[49113] <= 16'b0000_0000_0000_0000;
array[49114] <= 16'b0000_0000_0000_0000;
array[49115] <= 16'b0000_0000_0000_0000;
array[49116] <= 16'b0000_0000_0000_0000;
array[49117] <= 16'b0000_0000_0000_0000;
array[49118] <= 16'b0000_0000_0000_0000;
array[49119] <= 16'b0000_0000_0000_0000;
array[49120] <= 16'b0000_0000_0000_0000;
array[49121] <= 16'b0000_0000_0000_0000;
array[49122] <= 16'b0000_0000_0000_0000;
array[49123] <= 16'b0000_0000_0000_0000;
array[49124] <= 16'b0000_0000_0000_0000;
array[49125] <= 16'b0000_0000_0000_0000;
array[49126] <= 16'b0000_0000_0000_0000;
array[49127] <= 16'b0000_0000_0000_0000;
array[49128] <= 16'b0000_0000_0000_0000;
array[49129] <= 16'b0000_0000_0000_0000;
array[49130] <= 16'b0000_0000_0000_0000;
array[49131] <= 16'b0000_0000_0000_0000;
array[49132] <= 16'b0000_0000_0000_0000;
array[49133] <= 16'b0000_0000_0000_0000;
array[49134] <= 16'b0000_0000_0000_0000;
array[49135] <= 16'b0000_0000_0000_0000;
array[49136] <= 16'b0000_0000_0000_0000;
array[49137] <= 16'b0000_0000_0000_0000;
array[49138] <= 16'b0000_0000_0000_0000;
array[49139] <= 16'b0000_0000_0000_0000;
array[49140] <= 16'b0000_0000_0000_0000;
array[49141] <= 16'b0000_0000_0000_0000;
array[49142] <= 16'b0000_0000_0000_0000;
array[49143] <= 16'b0000_0000_0000_0000;
array[49144] <= 16'b0000_0000_0000_0000;
array[49145] <= 16'b0000_0000_0000_0000;
array[49146] <= 16'b0000_0000_0000_0000;
array[49147] <= 16'b0000_0000_0000_0000;
array[49148] <= 16'b0000_0000_0000_0000;
array[49149] <= 16'b0000_0000_0000_0000;
array[49150] <= 16'b0000_0000_0000_0000;
array[49151] <= 16'b0000_0000_0000_0000;
array[49152] <= 16'b0000_0000_0000_0000;
array[49153] <= 16'b0000_0000_0000_0000;
array[49154] <= 16'b0000_0000_0000_0000;
array[49155] <= 16'b0000_0000_0000_0000;
array[49156] <= 16'b0000_0000_0000_0000;
array[49157] <= 16'b0000_0000_0000_0000;
array[49158] <= 16'b0000_0000_0000_0000;
array[49159] <= 16'b0000_0000_0000_0000;
array[49160] <= 16'b0000_0000_0000_0000;
array[49161] <= 16'b0000_0000_0000_0000;
array[49162] <= 16'b0000_0000_0000_0000;
array[49163] <= 16'b0000_0000_0000_0000;
array[49164] <= 16'b0000_0000_0000_0000;
array[49165] <= 16'b0000_0000_0000_0000;
array[49166] <= 16'b0000_0000_0000_0000;
array[49167] <= 16'b0000_0000_0000_0000;
array[49168] <= 16'b0000_0000_0000_0000;
array[49169] <= 16'b0000_0000_0000_0000;
array[49170] <= 16'b0000_0000_0000_0000;
array[49171] <= 16'b0000_0000_0000_0000;
array[49172] <= 16'b0000_0000_0000_0000;
array[49173] <= 16'b0000_0000_0000_0000;
array[49174] <= 16'b0000_0000_0000_0000;
array[49175] <= 16'b0000_0000_0000_0000;
array[49176] <= 16'b0000_0000_0000_0000;
array[49177] <= 16'b0000_0000_0000_0000;
array[49178] <= 16'b0000_0000_0000_0000;
array[49179] <= 16'b0000_0000_0000_0000;
array[49180] <= 16'b0000_0000_0000_0000;
array[49181] <= 16'b0000_0000_0000_0000;
array[49182] <= 16'b0000_0000_0000_0000;
array[49183] <= 16'b0000_0000_0000_0000;
array[49184] <= 16'b0000_0000_0000_0000;
array[49185] <= 16'b0000_0000_0000_0000;
array[49186] <= 16'b0000_0000_0000_0000;
array[49187] <= 16'b0000_0000_0000_0000;
array[49188] <= 16'b0000_0000_0000_0000;
array[49189] <= 16'b0000_0000_0000_0000;
array[49190] <= 16'b0000_0000_0000_0000;
array[49191] <= 16'b0000_0000_0000_0000;
array[49192] <= 16'b0000_0000_0000_0000;
array[49193] <= 16'b0000_0000_0000_0000;
array[49194] <= 16'b0000_0000_0000_0000;
array[49195] <= 16'b0000_0000_0000_0000;
array[49196] <= 16'b0000_0000_0000_0000;
array[49197] <= 16'b0000_0000_0000_0000;
array[49198] <= 16'b0000_0000_0000_0000;
array[49199] <= 16'b0000_0000_0000_0000;
array[49200] <= 16'b0000_0000_0000_0000;
array[49201] <= 16'b0000_0000_0000_0000;
array[49202] <= 16'b0000_0000_0000_0000;
array[49203] <= 16'b0000_0000_0000_0000;
array[49204] <= 16'b0000_0000_0000_0000;
array[49205] <= 16'b0000_0000_0000_0000;
array[49206] <= 16'b0000_0000_0000_0000;
array[49207] <= 16'b0000_0000_0000_0000;
array[49208] <= 16'b0000_0000_0000_0000;
array[49209] <= 16'b0000_0000_0000_0000;
array[49210] <= 16'b0000_0000_0000_0000;
array[49211] <= 16'b0000_0000_0000_0000;
array[49212] <= 16'b0000_0000_0000_0000;
array[49213] <= 16'b0000_0000_0000_0000;
array[49214] <= 16'b0000_0000_0000_0000;
array[49215] <= 16'b0000_0000_0000_0000;
array[49216] <= 16'b0000_0000_0000_0000;
array[49217] <= 16'b0000_0000_0000_0000;
array[49218] <= 16'b0000_0000_0000_0000;
array[49219] <= 16'b0000_0000_0000_0000;
array[49220] <= 16'b0000_0000_0000_0000;
array[49221] <= 16'b0000_0000_0000_0000;
array[49222] <= 16'b0000_0000_0000_0000;
array[49223] <= 16'b0000_0000_0000_0000;
array[49224] <= 16'b0000_0000_0000_0000;
array[49225] <= 16'b0000_0000_0000_0000;
array[49226] <= 16'b0000_0000_0000_0000;
array[49227] <= 16'b0000_0000_0000_0000;
array[49228] <= 16'b0000_0000_0000_0000;
array[49229] <= 16'b0000_0000_0000_0000;
array[49230] <= 16'b0000_0000_0000_0000;
array[49231] <= 16'b0000_0000_0000_0000;
array[49232] <= 16'b0000_0000_0000_0000;
array[49233] <= 16'b0000_0000_0000_0000;
array[49234] <= 16'b0000_0000_0000_0000;
array[49235] <= 16'b0000_0000_0000_0000;
array[49236] <= 16'b0000_0000_0000_0000;
array[49237] <= 16'b0000_0000_0000_0000;
array[49238] <= 16'b0000_0000_0000_0000;
array[49239] <= 16'b0000_0000_0000_0000;
array[49240] <= 16'b0000_0000_0000_0000;
array[49241] <= 16'b0000_0000_0000_0000;
array[49242] <= 16'b0000_0000_0000_0000;
array[49243] <= 16'b0000_0000_0000_0000;
array[49244] <= 16'b0000_0000_0000_0000;
array[49245] <= 16'b0000_0000_0000_0000;
array[49246] <= 16'b0000_0000_0000_0000;
array[49247] <= 16'b0000_0000_0000_0000;
array[49248] <= 16'b0000_0000_0000_0000;
array[49249] <= 16'b0000_0000_0000_0000;
array[49250] <= 16'b0000_0000_0000_0000;
array[49251] <= 16'b0000_0000_0000_0000;
array[49252] <= 16'b0000_0000_0000_0000;
array[49253] <= 16'b0000_0000_0000_0000;
array[49254] <= 16'b0000_0000_0000_0000;
array[49255] <= 16'b0000_0000_0000_0000;
array[49256] <= 16'b0000_0000_0000_0000;
array[49257] <= 16'b0000_0000_0000_0000;
array[49258] <= 16'b0000_0000_0000_0000;
array[49259] <= 16'b0000_0000_0000_0000;
array[49260] <= 16'b0000_0000_0000_0000;
array[49261] <= 16'b0000_0000_0000_0000;
array[49262] <= 16'b0000_0000_0000_0000;
array[49263] <= 16'b0000_0000_0000_0000;
array[49264] <= 16'b0000_0000_0000_0000;
array[49265] <= 16'b0000_0000_0000_0000;
array[49266] <= 16'b0000_0000_0000_0000;
array[49267] <= 16'b0000_0000_0000_0000;
array[49268] <= 16'b0000_0000_0000_0000;
array[49269] <= 16'b0000_0000_0000_0000;
array[49270] <= 16'b0000_0000_0000_0000;
array[49271] <= 16'b0000_0000_0000_0000;
array[49272] <= 16'b0000_0000_0000_0000;
array[49273] <= 16'b0000_0000_0000_0000;
array[49274] <= 16'b0000_0000_0000_0000;
array[49275] <= 16'b0000_0000_0000_0000;
array[49276] <= 16'b0000_0000_0000_0000;
array[49277] <= 16'b0000_0000_0000_0000;
array[49278] <= 16'b0000_0000_0000_0000;
array[49279] <= 16'b0000_0000_0000_0000;
array[49280] <= 16'b0000_0000_0000_0000;
array[49281] <= 16'b0000_0000_0000_0000;
array[49282] <= 16'b0000_0000_0000_0000;
array[49283] <= 16'b0000_0000_0000_0000;
array[49284] <= 16'b0000_0000_0000_0000;
array[49285] <= 16'b0000_0000_0000_0000;
array[49286] <= 16'b0000_0000_0000_0000;
array[49287] <= 16'b0000_0000_0000_0000;
array[49288] <= 16'b0000_0000_0000_0000;
array[49289] <= 16'b0000_0000_0000_0000;
array[49290] <= 16'b0000_0000_0000_0000;
array[49291] <= 16'b0000_0000_0000_0000;
array[49292] <= 16'b0000_0000_0000_0000;
array[49293] <= 16'b0000_0000_0000_0000;
array[49294] <= 16'b0000_0000_0000_0000;
array[49295] <= 16'b0000_0000_0000_0000;
array[49296] <= 16'b0000_0000_0000_0000;
array[49297] <= 16'b0000_0000_0000_0000;
array[49298] <= 16'b0000_0000_0000_0000;
array[49299] <= 16'b0000_0000_0000_0000;
array[49300] <= 16'b0000_0000_0000_0000;
array[49301] <= 16'b0000_0000_0000_0000;
array[49302] <= 16'b0000_0000_0000_0000;
array[49303] <= 16'b0000_0000_0000_0000;
array[49304] <= 16'b0000_0000_0000_0000;
array[49305] <= 16'b0000_0000_0000_0000;
array[49306] <= 16'b0000_0000_0000_0000;
array[49307] <= 16'b0000_0000_0000_0000;
array[49308] <= 16'b0000_0000_0000_0000;
array[49309] <= 16'b0000_0000_0000_0000;
array[49310] <= 16'b0000_0000_0000_0000;
array[49311] <= 16'b0000_0000_0000_0000;
array[49312] <= 16'b0000_0000_0000_0000;
array[49313] <= 16'b0000_0000_0000_0000;
array[49314] <= 16'b0000_0000_0000_0000;
array[49315] <= 16'b0000_0000_0000_0000;
array[49316] <= 16'b0000_0000_0000_0000;
array[49317] <= 16'b0000_0000_0000_0000;
array[49318] <= 16'b0000_0000_0000_0000;
array[49319] <= 16'b0000_0000_0000_0000;
array[49320] <= 16'b0000_0000_0000_0000;
array[49321] <= 16'b0000_0000_0000_0000;
array[49322] <= 16'b0000_0000_0000_0000;
array[49323] <= 16'b0000_0000_0000_0000;
array[49324] <= 16'b0000_0000_0000_0000;
array[49325] <= 16'b0000_0000_0000_0000;
array[49326] <= 16'b0000_0000_0000_0000;
array[49327] <= 16'b0000_0000_0000_0000;
array[49328] <= 16'b0000_0000_0000_0000;
array[49329] <= 16'b0000_0000_0000_0000;
array[49330] <= 16'b0000_0000_0000_0000;
array[49331] <= 16'b0000_0000_0000_0000;
array[49332] <= 16'b0000_0000_0000_0000;
array[49333] <= 16'b0000_0000_0000_0000;
array[49334] <= 16'b0000_0000_0000_0000;
array[49335] <= 16'b0000_0000_0000_0000;
array[49336] <= 16'b0000_0000_0000_0000;
array[49337] <= 16'b0000_0000_0000_0000;
array[49338] <= 16'b0000_0000_0000_0000;
array[49339] <= 16'b0000_0000_0000_0000;
array[49340] <= 16'b0000_0000_0000_0000;
array[49341] <= 16'b0000_0000_0000_0000;
array[49342] <= 16'b0000_0000_0000_0000;
array[49343] <= 16'b0000_0000_0000_0000;
array[49344] <= 16'b0000_0000_0000_0000;
array[49345] <= 16'b0000_0000_0000_0000;
array[49346] <= 16'b0000_0000_0000_0000;
array[49347] <= 16'b0000_0000_0000_0000;
array[49348] <= 16'b0000_0000_0000_0000;
array[49349] <= 16'b0000_0000_0000_0000;
array[49350] <= 16'b0000_0000_0000_0000;
array[49351] <= 16'b0000_0000_0000_0000;
array[49352] <= 16'b0000_0000_0000_0000;
array[49353] <= 16'b0000_0000_0000_0000;
array[49354] <= 16'b0000_0000_0000_0000;
array[49355] <= 16'b0000_0000_0000_0000;
array[49356] <= 16'b0000_0000_0000_0000;
array[49357] <= 16'b0000_0000_0000_0000;
array[49358] <= 16'b0000_0000_0000_0000;
array[49359] <= 16'b0000_0000_0000_0000;
array[49360] <= 16'b0000_0000_0000_0000;
array[49361] <= 16'b0000_0000_0000_0000;
array[49362] <= 16'b0000_0000_0000_0000;
array[49363] <= 16'b0000_0000_0000_0000;
array[49364] <= 16'b0000_0000_0000_0000;
array[49365] <= 16'b0000_0000_0000_0000;
array[49366] <= 16'b0000_0000_0000_0000;
array[49367] <= 16'b0000_0000_0000_0000;
array[49368] <= 16'b0000_0000_0000_0000;
array[49369] <= 16'b0000_0000_0000_0000;
array[49370] <= 16'b0000_0000_0000_0000;
array[49371] <= 16'b0000_0000_0000_0000;
array[49372] <= 16'b0000_0000_0000_0000;
array[49373] <= 16'b0000_0000_0000_0000;
array[49374] <= 16'b0000_0000_0000_0000;
array[49375] <= 16'b0000_0000_0000_0000;
array[49376] <= 16'b0000_0000_0000_0000;
array[49377] <= 16'b0000_0000_0000_0000;
array[49378] <= 16'b0000_0000_0000_0000;
array[49379] <= 16'b0000_0000_0000_0000;
array[49380] <= 16'b0000_0000_0000_0000;
array[49381] <= 16'b0000_0000_0000_0000;
array[49382] <= 16'b0000_0000_0000_0000;
array[49383] <= 16'b0000_0000_0000_0000;
array[49384] <= 16'b0000_0000_0000_0000;
array[49385] <= 16'b0000_0000_0000_0000;
array[49386] <= 16'b0000_0000_0000_0000;
array[49387] <= 16'b0000_0000_0000_0000;
array[49388] <= 16'b0000_0000_0000_0000;
array[49389] <= 16'b0000_0000_0000_0000;
array[49390] <= 16'b0000_0000_0000_0000;
array[49391] <= 16'b0000_0000_0000_0000;
array[49392] <= 16'b0000_0000_0000_0000;
array[49393] <= 16'b0000_0000_0000_0000;
array[49394] <= 16'b0000_0000_0000_0000;
array[49395] <= 16'b0000_0000_0000_0000;
array[49396] <= 16'b0000_0000_0000_0000;
array[49397] <= 16'b0000_0000_0000_0000;
array[49398] <= 16'b0000_0000_0000_0000;
array[49399] <= 16'b0000_0000_0000_0000;
array[49400] <= 16'b0000_0000_0000_0000;
array[49401] <= 16'b0000_0000_0000_0000;
array[49402] <= 16'b0000_0000_0000_0000;
array[49403] <= 16'b0000_0000_0000_0000;
array[49404] <= 16'b0000_0000_0000_0000;
array[49405] <= 16'b0000_0000_0000_0000;
array[49406] <= 16'b0000_0000_0000_0000;
array[49407] <= 16'b0000_0000_0000_0000;
array[49408] <= 16'b0000_0000_0000_0000;
array[49409] <= 16'b0000_0000_0000_0000;
array[49410] <= 16'b0000_0000_0000_0000;
array[49411] <= 16'b0000_0000_0000_0000;
array[49412] <= 16'b0000_0000_0000_0000;
array[49413] <= 16'b0000_0000_0000_0000;
array[49414] <= 16'b0000_0000_0000_0000;
array[49415] <= 16'b0000_0000_0000_0000;
array[49416] <= 16'b0000_0000_0000_0000;
array[49417] <= 16'b0000_0000_0000_0000;
array[49418] <= 16'b0000_0000_0000_0000;
array[49419] <= 16'b0000_0000_0000_0000;
array[49420] <= 16'b0000_0000_0000_0000;
array[49421] <= 16'b0000_0000_0000_0000;
array[49422] <= 16'b0000_0000_0000_0000;
array[49423] <= 16'b0000_0000_0000_0000;
array[49424] <= 16'b0000_0000_0000_0000;
array[49425] <= 16'b0000_0000_0000_0000;
array[49426] <= 16'b0000_0000_0000_0000;
array[49427] <= 16'b0000_0000_0000_0000;
array[49428] <= 16'b0000_0000_0000_0000;
array[49429] <= 16'b0000_0000_0000_0000;
array[49430] <= 16'b0000_0000_0000_0000;
array[49431] <= 16'b0000_0000_0000_0000;
array[49432] <= 16'b0000_0000_0000_0000;
array[49433] <= 16'b0000_0000_0000_0000;
array[49434] <= 16'b0000_0000_0000_0000;
array[49435] <= 16'b0000_0000_0000_0000;
array[49436] <= 16'b0000_0000_0000_0000;
array[49437] <= 16'b0000_0000_0000_0000;
array[49438] <= 16'b0000_0000_0000_0000;
array[49439] <= 16'b0000_0000_0000_0000;
array[49440] <= 16'b0000_0000_0000_0000;
array[49441] <= 16'b0000_0000_0000_0000;
array[49442] <= 16'b0000_0000_0000_0000;
array[49443] <= 16'b0000_0000_0000_0000;
array[49444] <= 16'b0000_0000_0000_0000;
array[49445] <= 16'b0000_0000_0000_0000;
array[49446] <= 16'b0000_0000_0000_0000;
array[49447] <= 16'b0000_0000_0000_0000;
array[49448] <= 16'b0000_0000_0000_0000;
array[49449] <= 16'b0000_0000_0000_0000;
array[49450] <= 16'b0000_0000_0000_0000;
array[49451] <= 16'b0000_0000_0000_0000;
array[49452] <= 16'b0000_0000_0000_0000;
array[49453] <= 16'b0000_0000_0000_0000;
array[49454] <= 16'b0000_0000_0000_0000;
array[49455] <= 16'b0000_0000_0000_0000;
array[49456] <= 16'b0000_0000_0000_0000;
array[49457] <= 16'b0000_0000_0000_0000;
array[49458] <= 16'b0000_0000_0000_0000;
array[49459] <= 16'b0000_0000_0000_0000;
array[49460] <= 16'b0000_0000_0000_0000;
array[49461] <= 16'b0000_0000_0000_0000;
array[49462] <= 16'b0000_0000_0000_0000;
array[49463] <= 16'b0000_0000_0000_0000;
array[49464] <= 16'b0000_0000_0000_0000;
array[49465] <= 16'b0000_0000_0000_0000;
array[49466] <= 16'b0000_0000_0000_0000;
array[49467] <= 16'b0000_0000_0000_0000;
array[49468] <= 16'b0000_0000_0000_0000;
array[49469] <= 16'b0000_0000_0000_0000;
array[49470] <= 16'b0000_0000_0000_0000;
array[49471] <= 16'b0000_0000_0000_0000;
array[49472] <= 16'b0000_0000_0000_0000;
array[49473] <= 16'b0000_0000_0000_0000;
array[49474] <= 16'b0000_0000_0000_0000;
array[49475] <= 16'b0000_0000_0000_0000;
array[49476] <= 16'b0000_0000_0000_0000;
array[49477] <= 16'b0000_0000_0000_0000;
array[49478] <= 16'b0000_0000_0000_0000;
array[49479] <= 16'b0000_0000_0000_0000;
array[49480] <= 16'b0000_0000_0000_0000;
array[49481] <= 16'b0000_0000_0000_0000;
array[49482] <= 16'b0000_0000_0000_0000;
array[49483] <= 16'b0000_0000_0000_0000;
array[49484] <= 16'b0000_0000_0000_0000;
array[49485] <= 16'b0000_0000_0000_0000;
array[49486] <= 16'b0000_0000_0000_0000;
array[49487] <= 16'b0000_0000_0000_0000;
array[49488] <= 16'b0000_0000_0000_0000;
array[49489] <= 16'b0000_0000_0000_0000;
array[49490] <= 16'b0000_0000_0000_0000;
array[49491] <= 16'b0000_0000_0000_0000;
array[49492] <= 16'b0000_0000_0000_0000;
array[49493] <= 16'b0000_0000_0000_0000;
array[49494] <= 16'b0000_0000_0000_0000;
array[49495] <= 16'b0000_0000_0000_0000;
array[49496] <= 16'b0000_0000_0000_0000;
array[49497] <= 16'b0000_0000_0000_0000;
array[49498] <= 16'b0000_0000_0000_0000;
array[49499] <= 16'b0000_0000_0000_0000;
array[49500] <= 16'b0000_0000_0000_0000;
array[49501] <= 16'b0000_0000_0000_0000;
array[49502] <= 16'b0000_0000_0000_0000;
array[49503] <= 16'b0000_0000_0000_0000;
array[49504] <= 16'b0000_0000_0000_0000;
array[49505] <= 16'b0000_0000_0000_0000;
array[49506] <= 16'b0000_0000_0000_0000;
array[49507] <= 16'b0000_0000_0000_0000;
array[49508] <= 16'b0000_0000_0000_0000;
array[49509] <= 16'b0000_0000_0000_0000;
array[49510] <= 16'b0000_0000_0000_0000;
array[49511] <= 16'b0000_0000_0000_0000;
array[49512] <= 16'b0000_0000_0000_0000;
array[49513] <= 16'b0000_0000_0000_0000;
array[49514] <= 16'b0000_0000_0000_0000;
array[49515] <= 16'b0000_0000_0000_0000;
array[49516] <= 16'b0000_0000_0000_0000;
array[49517] <= 16'b0000_0000_0000_0000;
array[49518] <= 16'b0000_0000_0000_0000;
array[49519] <= 16'b0000_0000_0000_0000;
array[49520] <= 16'b0000_0000_0000_0000;
array[49521] <= 16'b0000_0000_0000_0000;
array[49522] <= 16'b0000_0000_0000_0000;
array[49523] <= 16'b0000_0000_0000_0000;
array[49524] <= 16'b0000_0000_0000_0000;
array[49525] <= 16'b0000_0000_0000_0000;
array[49526] <= 16'b0000_0000_0000_0000;
array[49527] <= 16'b0000_0000_0000_0000;
array[49528] <= 16'b0000_0000_0000_0000;
array[49529] <= 16'b0000_0000_0000_0000;
array[49530] <= 16'b0000_0000_0000_0000;
array[49531] <= 16'b0000_0000_0000_0000;
array[49532] <= 16'b0000_0000_0000_0000;
array[49533] <= 16'b0000_0000_0000_0000;
array[49534] <= 16'b0000_0000_0000_0000;
array[49535] <= 16'b0000_0000_0000_0000;
array[49536] <= 16'b0000_0000_0000_0000;
array[49537] <= 16'b0000_0000_0000_0000;
array[49538] <= 16'b0000_0000_0000_0000;
array[49539] <= 16'b0000_0000_0000_0000;
array[49540] <= 16'b0000_0000_0000_0000;
array[49541] <= 16'b0000_0000_0000_0000;
array[49542] <= 16'b0000_0000_0000_0000;
array[49543] <= 16'b0000_0000_0000_0000;
array[49544] <= 16'b0000_0000_0000_0000;
array[49545] <= 16'b0000_0000_0000_0000;
array[49546] <= 16'b0000_0000_0000_0000;
array[49547] <= 16'b0000_0000_0000_0000;
array[49548] <= 16'b0000_0000_0000_0000;
array[49549] <= 16'b0000_0000_0000_0000;
array[49550] <= 16'b0000_0000_0000_0000;
array[49551] <= 16'b0000_0000_0000_0000;
array[49552] <= 16'b0000_0000_0000_0000;
array[49553] <= 16'b0000_0000_0000_0000;
array[49554] <= 16'b0000_0000_0000_0000;
array[49555] <= 16'b0000_0000_0000_0000;
array[49556] <= 16'b0000_0000_0000_0000;
array[49557] <= 16'b0000_0000_0000_0000;
array[49558] <= 16'b0000_0000_0000_0000;
array[49559] <= 16'b0000_0000_0000_0000;
array[49560] <= 16'b0000_0000_0000_0000;
array[49561] <= 16'b0000_0000_0000_0000;
array[49562] <= 16'b0000_0000_0000_0000;
array[49563] <= 16'b0000_0000_0000_0000;
array[49564] <= 16'b0000_0000_0000_0000;
array[49565] <= 16'b0000_0000_0000_0000;
array[49566] <= 16'b0000_0000_0000_0000;
array[49567] <= 16'b0000_0000_0000_0000;
array[49568] <= 16'b0000_0000_0000_0000;
array[49569] <= 16'b0000_0000_0000_0000;
array[49570] <= 16'b0000_0000_0000_0000;
array[49571] <= 16'b0000_0000_0000_0000;
array[49572] <= 16'b0000_0000_0000_0000;
array[49573] <= 16'b0000_0000_0000_0000;
array[49574] <= 16'b0000_0000_0000_0000;
array[49575] <= 16'b0000_0000_0000_0000;
array[49576] <= 16'b0000_0000_0000_0000;
array[49577] <= 16'b0000_0000_0000_0000;
array[49578] <= 16'b0000_0000_0000_0000;
array[49579] <= 16'b0000_0000_0000_0000;
array[49580] <= 16'b0000_0000_0000_0000;
array[49581] <= 16'b0000_0000_0000_0000;
array[49582] <= 16'b0000_0000_0000_0000;
array[49583] <= 16'b0000_0000_0000_0000;
array[49584] <= 16'b0000_0000_0000_0000;
array[49585] <= 16'b0000_0000_0000_0000;
array[49586] <= 16'b0000_0000_0000_0000;
array[49587] <= 16'b0000_0000_0000_0000;
array[49588] <= 16'b0000_0000_0000_0000;
array[49589] <= 16'b0000_0000_0000_0000;
array[49590] <= 16'b0000_0000_0000_0000;
array[49591] <= 16'b0000_0000_0000_0000;
array[49592] <= 16'b0000_0000_0000_0000;
array[49593] <= 16'b0000_0000_0000_0000;
array[49594] <= 16'b0000_0000_0000_0000;
array[49595] <= 16'b0000_0000_0000_0000;
array[49596] <= 16'b0000_0000_0000_0000;
array[49597] <= 16'b0000_0000_0000_0000;
array[49598] <= 16'b0000_0000_0000_0000;
array[49599] <= 16'b0000_0000_0000_0000;
array[49600] <= 16'b0000_0000_0000_0000;
array[49601] <= 16'b0000_0000_0000_0000;
array[49602] <= 16'b0000_0000_0000_0000;
array[49603] <= 16'b0000_0000_0000_0000;
array[49604] <= 16'b0000_0000_0000_0000;
array[49605] <= 16'b0000_0000_0000_0000;
array[49606] <= 16'b0000_0000_0000_0000;
array[49607] <= 16'b0000_0000_0000_0000;
array[49608] <= 16'b0000_0000_0000_0000;
array[49609] <= 16'b0000_0000_0000_0000;
array[49610] <= 16'b0000_0000_0000_0000;
array[49611] <= 16'b0000_0000_0000_0000;
array[49612] <= 16'b0000_0000_0000_0000;
array[49613] <= 16'b0000_0000_0000_0000;
array[49614] <= 16'b0000_0000_0000_0000;
array[49615] <= 16'b0000_0000_0000_0000;
array[49616] <= 16'b0000_0000_0000_0000;
array[49617] <= 16'b0000_0000_0000_0000;
array[49618] <= 16'b0000_0000_0000_0000;
array[49619] <= 16'b0000_0000_0000_0000;
array[49620] <= 16'b0000_0000_0000_0000;
array[49621] <= 16'b0000_0000_0000_0000;
array[49622] <= 16'b0000_0000_0000_0000;
array[49623] <= 16'b0000_0000_0000_0000;
array[49624] <= 16'b0000_0000_0000_0000;
array[49625] <= 16'b0000_0000_0000_0000;
array[49626] <= 16'b0000_0000_0000_0000;
array[49627] <= 16'b0000_0000_0000_0000;
array[49628] <= 16'b0000_0000_0000_0000;
array[49629] <= 16'b0000_0000_0000_0000;
array[49630] <= 16'b0000_0000_0000_0000;
array[49631] <= 16'b0000_0000_0000_0000;
array[49632] <= 16'b0000_0000_0000_0000;
array[49633] <= 16'b0000_0000_0000_0000;
array[49634] <= 16'b0000_0000_0000_0000;
array[49635] <= 16'b0000_0000_0000_0000;
array[49636] <= 16'b0000_0000_0000_0000;
array[49637] <= 16'b0000_0000_0000_0000;
array[49638] <= 16'b0000_0000_0000_0000;
array[49639] <= 16'b0000_0000_0000_0000;
array[49640] <= 16'b0000_0000_0000_0000;
array[49641] <= 16'b0000_0000_0000_0000;
array[49642] <= 16'b0000_0000_0000_0000;
array[49643] <= 16'b0000_0000_0000_0000;
array[49644] <= 16'b0000_0000_0000_0000;
array[49645] <= 16'b0000_0000_0000_0000;
array[49646] <= 16'b0000_0000_0000_0000;
array[49647] <= 16'b0000_0000_0000_0000;
array[49648] <= 16'b0000_0000_0000_0000;
array[49649] <= 16'b0000_0000_0000_0000;
array[49650] <= 16'b0000_0000_0000_0000;
array[49651] <= 16'b0000_0000_0000_0000;
array[49652] <= 16'b0000_0000_0000_0000;
array[49653] <= 16'b0000_0000_0000_0000;
array[49654] <= 16'b0000_0000_0000_0000;
array[49655] <= 16'b0000_0000_0000_0000;
array[49656] <= 16'b0000_0000_0000_0000;
array[49657] <= 16'b0000_0000_0000_0000;
array[49658] <= 16'b0000_0000_0000_0000;
array[49659] <= 16'b0000_0000_0000_0000;
array[49660] <= 16'b0000_0000_0000_0000;
array[49661] <= 16'b0000_0000_0000_0000;
array[49662] <= 16'b0000_0000_0000_0000;
array[49663] <= 16'b0000_0000_0000_0000;
array[49664] <= 16'b0000_0000_0000_0000;
array[49665] <= 16'b0000_0000_0000_0000;
array[49666] <= 16'b0000_0000_0000_0000;
array[49667] <= 16'b0000_0000_0000_0000;
array[49668] <= 16'b0000_0000_0000_0000;
array[49669] <= 16'b0000_0000_0000_0000;
array[49670] <= 16'b0000_0000_0000_0000;
array[49671] <= 16'b0000_0000_0000_0000;
array[49672] <= 16'b0000_0000_0000_0000;
array[49673] <= 16'b0000_0000_0000_0000;
array[49674] <= 16'b0000_0000_0000_0000;
array[49675] <= 16'b0000_0000_0000_0000;
array[49676] <= 16'b0000_0000_0000_0000;
array[49677] <= 16'b0000_0000_0000_0000;
array[49678] <= 16'b0000_0000_0000_0000;
array[49679] <= 16'b0000_0000_0000_0000;
array[49680] <= 16'b0000_0000_0000_0000;
array[49681] <= 16'b0000_0000_0000_0000;
array[49682] <= 16'b0000_0000_0000_0000;
array[49683] <= 16'b0000_0000_0000_0000;
array[49684] <= 16'b0000_0000_0000_0000;
array[49685] <= 16'b0000_0000_0000_0000;
array[49686] <= 16'b0000_0000_0000_0000;
array[49687] <= 16'b0000_0000_0000_0000;
array[49688] <= 16'b0000_0000_0000_0000;
array[49689] <= 16'b0000_0000_0000_0000;
array[49690] <= 16'b0000_0000_0000_0000;
array[49691] <= 16'b0000_0000_0000_0000;
array[49692] <= 16'b0000_0000_0000_0000;
array[49693] <= 16'b0000_0000_0000_0000;
array[49694] <= 16'b0000_0000_0000_0000;
array[49695] <= 16'b0000_0000_0000_0000;
array[49696] <= 16'b0000_0000_0000_0000;
array[49697] <= 16'b0000_0000_0000_0000;
array[49698] <= 16'b0000_0000_0000_0000;
array[49699] <= 16'b0000_0000_0000_0000;
array[49700] <= 16'b0000_0000_0000_0000;
array[49701] <= 16'b0000_0000_0000_0000;
array[49702] <= 16'b0000_0000_0000_0000;
array[49703] <= 16'b0000_0000_0000_0000;
array[49704] <= 16'b0000_0000_0000_0000;
array[49705] <= 16'b0000_0000_0000_0000;
array[49706] <= 16'b0000_0000_0000_0000;
array[49707] <= 16'b0000_0000_0000_0000;
array[49708] <= 16'b0000_0000_0000_0000;
array[49709] <= 16'b0000_0000_0000_0000;
array[49710] <= 16'b0000_0000_0000_0000;
array[49711] <= 16'b0000_0000_0000_0000;
array[49712] <= 16'b0000_0000_0000_0000;
array[49713] <= 16'b0000_0000_0000_0000;
array[49714] <= 16'b0000_0000_0000_0000;
array[49715] <= 16'b0000_0000_0000_0000;
array[49716] <= 16'b0000_0000_0000_0000;
array[49717] <= 16'b0000_0000_0000_0000;
array[49718] <= 16'b0000_0000_0000_0000;
array[49719] <= 16'b0000_0000_0000_0000;
array[49720] <= 16'b0000_0000_0000_0000;
array[49721] <= 16'b0000_0000_0000_0000;
array[49722] <= 16'b0000_0000_0000_0000;
array[49723] <= 16'b0000_0000_0000_0000;
array[49724] <= 16'b0000_0000_0000_0000;
array[49725] <= 16'b0000_0000_0000_0000;
array[49726] <= 16'b0000_0000_0000_0000;
array[49727] <= 16'b0000_0000_0000_0000;
array[49728] <= 16'b0000_0000_0000_0000;
array[49729] <= 16'b0000_0000_0000_0000;
array[49730] <= 16'b0000_0000_0000_0000;
array[49731] <= 16'b0000_0000_0000_0000;
array[49732] <= 16'b0000_0000_0000_0000;
array[49733] <= 16'b0000_0000_0000_0000;
array[49734] <= 16'b0000_0000_0000_0000;
array[49735] <= 16'b0000_0000_0000_0000;
array[49736] <= 16'b0000_0000_0000_0000;
array[49737] <= 16'b0000_0000_0000_0000;
array[49738] <= 16'b0000_0000_0000_0000;
array[49739] <= 16'b0000_0000_0000_0000;
array[49740] <= 16'b0000_0000_0000_0000;
array[49741] <= 16'b0000_0000_0000_0000;
array[49742] <= 16'b0000_0000_0000_0000;
array[49743] <= 16'b0000_0000_0000_0000;
array[49744] <= 16'b0000_0000_0000_0000;
array[49745] <= 16'b0000_0000_0000_0000;
array[49746] <= 16'b0000_0000_0000_0000;
array[49747] <= 16'b0000_0000_0000_0000;
array[49748] <= 16'b0000_0000_0000_0000;
array[49749] <= 16'b0000_0000_0000_0000;
array[49750] <= 16'b0000_0000_0000_0000;
array[49751] <= 16'b0000_0000_0000_0000;
array[49752] <= 16'b0000_0000_0000_0000;
array[49753] <= 16'b0000_0000_0000_0000;
array[49754] <= 16'b0000_0000_0000_0000;
array[49755] <= 16'b0000_0000_0000_0000;
array[49756] <= 16'b0000_0000_0000_0000;
array[49757] <= 16'b0000_0000_0000_0000;
array[49758] <= 16'b0000_0000_0000_0000;
array[49759] <= 16'b0000_0000_0000_0000;
array[49760] <= 16'b0000_0000_0000_0000;
array[49761] <= 16'b0000_0000_0000_0000;
array[49762] <= 16'b0000_0000_0000_0000;
array[49763] <= 16'b0000_0000_0000_0000;
array[49764] <= 16'b0000_0000_0000_0000;
array[49765] <= 16'b0000_0000_0000_0000;
array[49766] <= 16'b0000_0000_0000_0000;
array[49767] <= 16'b0000_0000_0000_0000;
array[49768] <= 16'b0000_0000_0000_0000;
array[49769] <= 16'b0000_0000_0000_0000;
array[49770] <= 16'b0000_0000_0000_0000;
array[49771] <= 16'b0000_0000_0000_0000;
array[49772] <= 16'b0000_0000_0000_0000;
array[49773] <= 16'b0000_0000_0000_0000;
array[49774] <= 16'b0000_0000_0000_0000;
array[49775] <= 16'b0000_0000_0000_0000;
array[49776] <= 16'b0000_0000_0000_0000;
array[49777] <= 16'b0000_0000_0000_0000;
array[49778] <= 16'b0000_0000_0000_0000;
array[49779] <= 16'b0000_0000_0000_0000;
array[49780] <= 16'b0000_0000_0000_0000;
array[49781] <= 16'b0000_0000_0000_0000;
array[49782] <= 16'b0000_0000_0000_0000;
array[49783] <= 16'b0000_0000_0000_0000;
array[49784] <= 16'b0000_0000_0000_0000;
array[49785] <= 16'b0000_0000_0000_0000;
array[49786] <= 16'b0000_0000_0000_0000;
array[49787] <= 16'b0000_0000_0000_0000;
array[49788] <= 16'b0000_0000_0000_0000;
array[49789] <= 16'b0000_0000_0000_0000;
array[49790] <= 16'b0000_0000_0000_0000;
array[49791] <= 16'b0000_0000_0000_0000;
array[49792] <= 16'b0000_0000_0000_0000;
array[49793] <= 16'b0000_0000_0000_0000;
array[49794] <= 16'b0000_0000_0000_0000;
array[49795] <= 16'b0000_0000_0000_0000;
array[49796] <= 16'b0000_0000_0000_0000;
array[49797] <= 16'b0000_0000_0000_0000;
array[49798] <= 16'b0000_0000_0000_0000;
array[49799] <= 16'b0000_0000_0000_0000;
array[49800] <= 16'b0000_0000_0000_0000;
array[49801] <= 16'b0000_0000_0000_0000;
array[49802] <= 16'b0000_0000_0000_0000;
array[49803] <= 16'b0000_0000_0000_0000;
array[49804] <= 16'b0000_0000_0000_0000;
array[49805] <= 16'b0000_0000_0000_0000;
array[49806] <= 16'b0000_0000_0000_0000;
array[49807] <= 16'b0000_0000_0000_0000;
array[49808] <= 16'b0000_0000_0000_0000;
array[49809] <= 16'b0000_0000_0000_0000;
array[49810] <= 16'b0000_0000_0000_0000;
array[49811] <= 16'b0000_0000_0000_0000;
array[49812] <= 16'b0000_0000_0000_0000;
array[49813] <= 16'b0000_0000_0000_0000;
array[49814] <= 16'b0000_0000_0000_0000;
array[49815] <= 16'b0000_0000_0000_0000;
array[49816] <= 16'b0000_0000_0000_0000;
array[49817] <= 16'b0000_0000_0000_0000;
array[49818] <= 16'b0000_0000_0000_0000;
array[49819] <= 16'b0000_0000_0000_0000;
array[49820] <= 16'b0000_0000_0000_0000;
array[49821] <= 16'b0000_0000_0000_0000;
array[49822] <= 16'b0000_0000_0000_0000;
array[49823] <= 16'b0000_0000_0000_0000;
array[49824] <= 16'b0000_0000_0000_0000;
array[49825] <= 16'b0000_0000_0000_0000;
array[49826] <= 16'b0000_0000_0000_0000;
array[49827] <= 16'b0000_0000_0000_0000;
array[49828] <= 16'b0000_0000_0000_0000;
array[49829] <= 16'b0000_0000_0000_0000;
array[49830] <= 16'b0000_0000_0000_0000;
array[49831] <= 16'b0000_0000_0000_0000;
array[49832] <= 16'b0000_0000_0000_0000;
array[49833] <= 16'b0000_0000_0000_0000;
array[49834] <= 16'b0000_0000_0000_0000;
array[49835] <= 16'b0000_0000_0000_0000;
array[49836] <= 16'b0000_0000_0000_0000;
array[49837] <= 16'b0000_0000_0000_0000;
array[49838] <= 16'b0000_0000_0000_0000;
array[49839] <= 16'b0000_0000_0000_0000;
array[49840] <= 16'b0000_0000_0000_0000;
array[49841] <= 16'b0000_0000_0000_0000;
array[49842] <= 16'b0000_0000_0000_0000;
array[49843] <= 16'b0000_0000_0000_0000;
array[49844] <= 16'b0000_0000_0000_0000;
array[49845] <= 16'b0000_0000_0000_0000;
array[49846] <= 16'b0000_0000_0000_0000;
array[49847] <= 16'b0000_0000_0000_0000;
array[49848] <= 16'b0000_0000_0000_0000;
array[49849] <= 16'b0000_0000_0000_0000;
array[49850] <= 16'b0000_0000_0000_0000;
array[49851] <= 16'b0000_0000_0000_0000;
array[49852] <= 16'b0000_0000_0000_0000;
array[49853] <= 16'b0000_0000_0000_0000;
array[49854] <= 16'b0000_0000_0000_0000;
array[49855] <= 16'b0000_0000_0000_0000;
array[49856] <= 16'b0000_0000_0000_0000;
array[49857] <= 16'b0000_0000_0000_0000;
array[49858] <= 16'b0000_0000_0000_0000;
array[49859] <= 16'b0000_0000_0000_0000;
array[49860] <= 16'b0000_0000_0000_0000;
array[49861] <= 16'b0000_0000_0000_0000;
array[49862] <= 16'b0000_0000_0000_0000;
array[49863] <= 16'b0000_0000_0000_0000;
array[49864] <= 16'b0000_0000_0000_0000;
array[49865] <= 16'b0000_0000_0000_0000;
array[49866] <= 16'b0000_0000_0000_0000;
array[49867] <= 16'b0000_0000_0000_0000;
array[49868] <= 16'b0000_0000_0000_0000;
array[49869] <= 16'b0000_0000_0000_0000;
array[49870] <= 16'b0000_0000_0000_0000;
array[49871] <= 16'b0000_0000_0000_0000;
array[49872] <= 16'b0000_0000_0000_0000;
array[49873] <= 16'b0000_0000_0000_0000;
array[49874] <= 16'b0000_0000_0000_0000;
array[49875] <= 16'b0000_0000_0000_0000;
array[49876] <= 16'b0000_0000_0000_0000;
array[49877] <= 16'b0000_0000_0000_0000;
array[49878] <= 16'b0000_0000_0000_0000;
array[49879] <= 16'b0000_0000_0000_0000;
array[49880] <= 16'b0000_0000_0000_0000;
array[49881] <= 16'b0000_0000_0000_0000;
array[49882] <= 16'b0000_0000_0000_0000;
array[49883] <= 16'b0000_0000_0000_0000;
array[49884] <= 16'b0000_0000_0000_0000;
array[49885] <= 16'b0000_0000_0000_0000;
array[49886] <= 16'b0000_0000_0000_0000;
array[49887] <= 16'b0000_0000_0000_0000;
array[49888] <= 16'b0000_0000_0000_0000;
array[49889] <= 16'b0000_0000_0000_0000;
array[49890] <= 16'b0000_0000_0000_0000;
array[49891] <= 16'b0000_0000_0000_0000;
array[49892] <= 16'b0000_0000_0000_0000;
array[49893] <= 16'b0000_0000_0000_0000;
array[49894] <= 16'b0000_0000_0000_0000;
array[49895] <= 16'b0000_0000_0000_0000;
array[49896] <= 16'b0000_0000_0000_0000;
array[49897] <= 16'b0000_0000_0000_0000;
array[49898] <= 16'b0000_0000_0000_0000;
array[49899] <= 16'b0000_0000_0000_0000;
array[49900] <= 16'b0000_0000_0000_0000;
array[49901] <= 16'b0000_0000_0000_0000;
array[49902] <= 16'b0000_0000_0000_0000;
array[49903] <= 16'b0000_0000_0000_0000;
array[49904] <= 16'b0000_0000_0000_0000;
array[49905] <= 16'b0000_0000_0000_0000;
array[49906] <= 16'b0000_0000_0000_0000;
array[49907] <= 16'b0000_0000_0000_0000;
array[49908] <= 16'b0000_0000_0000_0000;
array[49909] <= 16'b0000_0000_0000_0000;
array[49910] <= 16'b0000_0000_0000_0000;
array[49911] <= 16'b0000_0000_0000_0000;
array[49912] <= 16'b0000_0000_0000_0000;
array[49913] <= 16'b0000_0000_0000_0000;
array[49914] <= 16'b0000_0000_0000_0000;
array[49915] <= 16'b0000_0000_0000_0000;
array[49916] <= 16'b0000_0000_0000_0000;
array[49917] <= 16'b0000_0000_0000_0000;
array[49918] <= 16'b0000_0000_0000_0000;
array[49919] <= 16'b0000_0000_0000_0000;
array[49920] <= 16'b0000_0000_0000_0000;
array[49921] <= 16'b0000_0000_0000_0000;
array[49922] <= 16'b0000_0000_0000_0000;
array[49923] <= 16'b0000_0000_0000_0000;
array[49924] <= 16'b0000_0000_0000_0000;
array[49925] <= 16'b0000_0000_0000_0000;
array[49926] <= 16'b0000_0000_0000_0000;
array[49927] <= 16'b0000_0000_0000_0000;
array[49928] <= 16'b0000_0000_0000_0000;
array[49929] <= 16'b0000_0000_0000_0000;
array[49930] <= 16'b0000_0000_0000_0000;
array[49931] <= 16'b0000_0000_0000_0000;
array[49932] <= 16'b0000_0000_0000_0000;
array[49933] <= 16'b0000_0000_0000_0000;
array[49934] <= 16'b0000_0000_0000_0000;
array[49935] <= 16'b0000_0000_0000_0000;
array[49936] <= 16'b0000_0000_0000_0000;
array[49937] <= 16'b0000_0000_0000_0000;
array[49938] <= 16'b0000_0000_0000_0000;
array[49939] <= 16'b0000_0000_0000_0000;
array[49940] <= 16'b0000_0000_0000_0000;
array[49941] <= 16'b0000_0000_0000_0000;
array[49942] <= 16'b0000_0000_0000_0000;
array[49943] <= 16'b0000_0000_0000_0000;
array[49944] <= 16'b0000_0000_0000_0000;
array[49945] <= 16'b0000_0000_0000_0000;
array[49946] <= 16'b0000_0000_0000_0000;
array[49947] <= 16'b0000_0000_0000_0000;
array[49948] <= 16'b0000_0000_0000_0000;
array[49949] <= 16'b0000_0000_0000_0000;
array[49950] <= 16'b0000_0000_0000_0000;
array[49951] <= 16'b0000_0000_0000_0000;
array[49952] <= 16'b0000_0000_0000_0000;
array[49953] <= 16'b0000_0000_0000_0000;
array[49954] <= 16'b0000_0000_0000_0000;
array[49955] <= 16'b0000_0000_0000_0000;
array[49956] <= 16'b0000_0000_0000_0000;
array[49957] <= 16'b0000_0000_0000_0000;
array[49958] <= 16'b0000_0000_0000_0000;
array[49959] <= 16'b0000_0000_0000_0000;
array[49960] <= 16'b0000_0000_0000_0000;
array[49961] <= 16'b0000_0000_0000_0000;
array[49962] <= 16'b0000_0000_0000_0000;
array[49963] <= 16'b0000_0000_0000_0000;
array[49964] <= 16'b0000_0000_0000_0000;
array[49965] <= 16'b0000_0000_0000_0000;
array[49966] <= 16'b0000_0000_0000_0000;
array[49967] <= 16'b0000_0000_0000_0000;
array[49968] <= 16'b0000_0000_0000_0000;
array[49969] <= 16'b0000_0000_0000_0000;
array[49970] <= 16'b0000_0000_0000_0000;
array[49971] <= 16'b0000_0000_0000_0000;
array[49972] <= 16'b0000_0000_0000_0000;
array[49973] <= 16'b0000_0000_0000_0000;
array[49974] <= 16'b0000_0000_0000_0000;
array[49975] <= 16'b0000_0000_0000_0000;
array[49976] <= 16'b0000_0000_0000_0000;
array[49977] <= 16'b0000_0000_0000_0000;
array[49978] <= 16'b0000_0000_0000_0000;
array[49979] <= 16'b0000_0000_0000_0000;
array[49980] <= 16'b0000_0000_0000_0000;
array[49981] <= 16'b0000_0000_0000_0000;
array[49982] <= 16'b0000_0000_0000_0000;
array[49983] <= 16'b0000_0000_0000_0000;
array[49984] <= 16'b0000_0000_0000_0000;
array[49985] <= 16'b0000_0000_0000_0000;
array[49986] <= 16'b0000_0000_0000_0000;
array[49987] <= 16'b0000_0000_0000_0000;
array[49988] <= 16'b0000_0000_0000_0000;
array[49989] <= 16'b0000_0000_0000_0000;
array[49990] <= 16'b0000_0000_0000_0000;
array[49991] <= 16'b0000_0000_0000_0000;
array[49992] <= 16'b0000_0000_0000_0000;
array[49993] <= 16'b0000_0000_0000_0000;
array[49994] <= 16'b0000_0000_0000_0000;
array[49995] <= 16'b0000_0000_0000_0000;
array[49996] <= 16'b0000_0000_0000_0000;
array[49997] <= 16'b0000_0000_0000_0000;
array[49998] <= 16'b0000_0000_0000_0000;
array[49999] <= 16'b0000_0000_0000_0000;
array[50000] <= 16'b0000_0000_0000_0000;
array[50001] <= 16'b0000_0000_0000_0000;
array[50002] <= 16'b0000_0000_0000_0000;
array[50003] <= 16'b0000_0000_0000_0000;
array[50004] <= 16'b0000_0000_0000_0000;
array[50005] <= 16'b0000_0000_0000_0000;
array[50006] <= 16'b0000_0000_0000_0000;
array[50007] <= 16'b0000_0000_0000_0000;
array[50008] <= 16'b0000_0000_0000_0000;
array[50009] <= 16'b0000_0000_0000_0000;
array[50010] <= 16'b0000_0000_0000_0000;
array[50011] <= 16'b0000_0000_0000_0000;
array[50012] <= 16'b0000_0000_0000_0000;
array[50013] <= 16'b0000_0000_0000_0000;
array[50014] <= 16'b0000_0000_0000_0000;
array[50015] <= 16'b0000_0000_0000_0000;
array[50016] <= 16'b0000_0000_0000_0000;
array[50017] <= 16'b0000_0000_0000_0000;
array[50018] <= 16'b0000_0000_0000_0000;
array[50019] <= 16'b0000_0000_0000_0000;
array[50020] <= 16'b0000_0000_0000_0000;
array[50021] <= 16'b0000_0000_0000_0000;
array[50022] <= 16'b0000_0000_0000_0000;
array[50023] <= 16'b0000_0000_0000_0000;
array[50024] <= 16'b0000_0000_0000_0000;
array[50025] <= 16'b0000_0000_0000_0000;
array[50026] <= 16'b0000_0000_0000_0000;
array[50027] <= 16'b0000_0000_0000_0000;
array[50028] <= 16'b0000_0000_0000_0000;
array[50029] <= 16'b0000_0000_0000_0000;
array[50030] <= 16'b0000_0000_0000_0000;
array[50031] <= 16'b0000_0000_0000_0000;
array[50032] <= 16'b0000_0000_0000_0000;
array[50033] <= 16'b0000_0000_0000_0000;
array[50034] <= 16'b0000_0000_0000_0000;
array[50035] <= 16'b0000_0000_0000_0000;
array[50036] <= 16'b0000_0000_0000_0000;
array[50037] <= 16'b0000_0000_0000_0000;
array[50038] <= 16'b0000_0000_0000_0000;
array[50039] <= 16'b0000_0000_0000_0000;
array[50040] <= 16'b0000_0000_0000_0000;
array[50041] <= 16'b0000_0000_0000_0000;
array[50042] <= 16'b0000_0000_0000_0000;
array[50043] <= 16'b0000_0000_0000_0000;
array[50044] <= 16'b0000_0000_0000_0000;
array[50045] <= 16'b0000_0000_0000_0000;
array[50046] <= 16'b0000_0000_0000_0000;
array[50047] <= 16'b0000_0000_0000_0000;
array[50048] <= 16'b0000_0000_0000_0000;
array[50049] <= 16'b0000_0000_0000_0000;
array[50050] <= 16'b0000_0000_0000_0000;
array[50051] <= 16'b0000_0000_0000_0000;
array[50052] <= 16'b0000_0000_0000_0000;
array[50053] <= 16'b0000_0000_0000_0000;
array[50054] <= 16'b0000_0000_0000_0000;
array[50055] <= 16'b0000_0000_0000_0000;
array[50056] <= 16'b0000_0000_0000_0000;
array[50057] <= 16'b0000_0000_0000_0000;
array[50058] <= 16'b0000_0000_0000_0000;
array[50059] <= 16'b0000_0000_0000_0000;
array[50060] <= 16'b0000_0000_0000_0000;
array[50061] <= 16'b0000_0000_0000_0000;
array[50062] <= 16'b0000_0000_0000_0000;
array[50063] <= 16'b0000_0000_0000_0000;
array[50064] <= 16'b0000_0000_0000_0000;
array[50065] <= 16'b0000_0000_0000_0000;
array[50066] <= 16'b0000_0000_0000_0000;
array[50067] <= 16'b0000_0000_0000_0000;
array[50068] <= 16'b0000_0000_0000_0000;
array[50069] <= 16'b0000_0000_0000_0000;
array[50070] <= 16'b0000_0000_0000_0000;
array[50071] <= 16'b0000_0000_0000_0000;
array[50072] <= 16'b0000_0000_0000_0000;
array[50073] <= 16'b0000_0000_0000_0000;
array[50074] <= 16'b0000_0000_0000_0000;
array[50075] <= 16'b0000_0000_0000_0000;
array[50076] <= 16'b0000_0000_0000_0000;
array[50077] <= 16'b0000_0000_0000_0000;
array[50078] <= 16'b0000_0000_0000_0000;
array[50079] <= 16'b0000_0000_0000_0000;
array[50080] <= 16'b0000_0000_0000_0000;
array[50081] <= 16'b0000_0000_0000_0000;
array[50082] <= 16'b0000_0000_0000_0000;
array[50083] <= 16'b0000_0000_0000_0000;
array[50084] <= 16'b0000_0000_0000_0000;
array[50085] <= 16'b0000_0000_0000_0000;
array[50086] <= 16'b0000_0000_0000_0000;
array[50087] <= 16'b0000_0000_0000_0000;
array[50088] <= 16'b0000_0000_0000_0000;
array[50089] <= 16'b0000_0000_0000_0000;
array[50090] <= 16'b0000_0000_0000_0000;
array[50091] <= 16'b0000_0000_0000_0000;
array[50092] <= 16'b0000_0000_0000_0000;
array[50093] <= 16'b0000_0000_0000_0000;
array[50094] <= 16'b0000_0000_0000_0000;
array[50095] <= 16'b0000_0000_0000_0000;
array[50096] <= 16'b0000_0000_0000_0000;
array[50097] <= 16'b0000_0000_0000_0000;
array[50098] <= 16'b0000_0000_0000_0000;
array[50099] <= 16'b0000_0000_0000_0000;
array[50100] <= 16'b0000_0000_0000_0000;
array[50101] <= 16'b0000_0000_0000_0000;
array[50102] <= 16'b0000_0000_0000_0000;
array[50103] <= 16'b0000_0000_0000_0000;
array[50104] <= 16'b0000_0000_0000_0000;
array[50105] <= 16'b0000_0000_0000_0000;
array[50106] <= 16'b0000_0000_0000_0000;
array[50107] <= 16'b0000_0000_0000_0000;
array[50108] <= 16'b0000_0000_0000_0000;
array[50109] <= 16'b0000_0000_0000_0000;
array[50110] <= 16'b0000_0000_0000_0000;
array[50111] <= 16'b0000_0000_0000_0000;
array[50112] <= 16'b0000_0000_0000_0000;
array[50113] <= 16'b0000_0000_0000_0000;
array[50114] <= 16'b0000_0000_0000_0000;
array[50115] <= 16'b0000_0000_0000_0000;
array[50116] <= 16'b0000_0000_0000_0000;
array[50117] <= 16'b0000_0000_0000_0000;
array[50118] <= 16'b0000_0000_0000_0000;
array[50119] <= 16'b0000_0000_0000_0000;
array[50120] <= 16'b0000_0000_0000_0000;
array[50121] <= 16'b0000_0000_0000_0000;
array[50122] <= 16'b0000_0000_0000_0000;
array[50123] <= 16'b0000_0000_0000_0000;
array[50124] <= 16'b0000_0000_0000_0000;
array[50125] <= 16'b0000_0000_0000_0000;
array[50126] <= 16'b0000_0000_0000_0000;
array[50127] <= 16'b0000_0000_0000_0000;
array[50128] <= 16'b0000_0000_0000_0000;
array[50129] <= 16'b0000_0000_0000_0000;
array[50130] <= 16'b0000_0000_0000_0000;
array[50131] <= 16'b0000_0000_0000_0000;
array[50132] <= 16'b0000_0000_0000_0000;
array[50133] <= 16'b0000_0000_0000_0000;
array[50134] <= 16'b0000_0000_0000_0000;
array[50135] <= 16'b0000_0000_0000_0000;
array[50136] <= 16'b0000_0000_0000_0000;
array[50137] <= 16'b0000_0000_0000_0000;
array[50138] <= 16'b0000_0000_0000_0000;
array[50139] <= 16'b0000_0000_0000_0000;
array[50140] <= 16'b0000_0000_0000_0000;
array[50141] <= 16'b0000_0000_0000_0000;
array[50142] <= 16'b0000_0000_0000_0000;
array[50143] <= 16'b0000_0000_0000_0000;
array[50144] <= 16'b0000_0000_0000_0000;
array[50145] <= 16'b0000_0000_0000_0000;
array[50146] <= 16'b0000_0000_0000_0000;
array[50147] <= 16'b0000_0000_0000_0000;
array[50148] <= 16'b0000_0000_0000_0000;
array[50149] <= 16'b0000_0000_0000_0000;
array[50150] <= 16'b0000_0000_0000_0000;
array[50151] <= 16'b0000_0000_0000_0000;
array[50152] <= 16'b0000_0000_0000_0000;
array[50153] <= 16'b0000_0000_0000_0000;
array[50154] <= 16'b0000_0000_0000_0000;
array[50155] <= 16'b0000_0000_0000_0000;
array[50156] <= 16'b0000_0000_0000_0000;
array[50157] <= 16'b0000_0000_0000_0000;
array[50158] <= 16'b0000_0000_0000_0000;
array[50159] <= 16'b0000_0000_0000_0000;
array[50160] <= 16'b0000_0000_0000_0000;
array[50161] <= 16'b0000_0000_0000_0000;
array[50162] <= 16'b0000_0000_0000_0000;
array[50163] <= 16'b0000_0000_0000_0000;
array[50164] <= 16'b0000_0000_0000_0000;
array[50165] <= 16'b0000_0000_0000_0000;
array[50166] <= 16'b0000_0000_0000_0000;
array[50167] <= 16'b0000_0000_0000_0000;
array[50168] <= 16'b0000_0000_0000_0000;
array[50169] <= 16'b0000_0000_0000_0000;
array[50170] <= 16'b0000_0000_0000_0000;
array[50171] <= 16'b0000_0000_0000_0000;
array[50172] <= 16'b0000_0000_0000_0000;
array[50173] <= 16'b0000_0000_0000_0000;
array[50174] <= 16'b0000_0000_0000_0000;
array[50175] <= 16'b0000_0000_0000_0000;
array[50176] <= 16'b0000_0000_0000_0000;
array[50177] <= 16'b0000_0000_0000_0000;
array[50178] <= 16'b0000_0000_0000_0000;
array[50179] <= 16'b0000_0000_0000_0000;
array[50180] <= 16'b0000_0000_0000_0000;
array[50181] <= 16'b0000_0000_0000_0000;
array[50182] <= 16'b0000_0000_0000_0000;
array[50183] <= 16'b0000_0000_0000_0000;
array[50184] <= 16'b0000_0000_0000_0000;
array[50185] <= 16'b0000_0000_0000_0000;
array[50186] <= 16'b0000_0000_0000_0000;
array[50187] <= 16'b0000_0000_0000_0000;
array[50188] <= 16'b0000_0000_0000_0000;
array[50189] <= 16'b0000_0000_0000_0000;
array[50190] <= 16'b0000_0000_0000_0000;
array[50191] <= 16'b0000_0000_0000_0000;
array[50192] <= 16'b0000_0000_0000_0000;
array[50193] <= 16'b0000_0000_0000_0000;
array[50194] <= 16'b0000_0000_0000_0000;
array[50195] <= 16'b0000_0000_0000_0000;
array[50196] <= 16'b0000_0000_0000_0000;
array[50197] <= 16'b0000_0000_0000_0000;
array[50198] <= 16'b0000_0000_0000_0000;
array[50199] <= 16'b0000_0000_0000_0000;
array[50200] <= 16'b0000_0000_0000_0000;
array[50201] <= 16'b0000_0000_0000_0000;
array[50202] <= 16'b0000_0000_0000_0000;
array[50203] <= 16'b0000_0000_0000_0000;
array[50204] <= 16'b0000_0000_0000_0000;
array[50205] <= 16'b0000_0000_0000_0000;
array[50206] <= 16'b0000_0000_0000_0000;
array[50207] <= 16'b0000_0000_0000_0000;
array[50208] <= 16'b0000_0000_0000_0000;
array[50209] <= 16'b0000_0000_0000_0000;
array[50210] <= 16'b0000_0000_0000_0000;
array[50211] <= 16'b0000_0000_0000_0000;
array[50212] <= 16'b0000_0000_0000_0000;
array[50213] <= 16'b0000_0000_0000_0000;
array[50214] <= 16'b0000_0000_0000_0000;
array[50215] <= 16'b0000_0000_0000_0000;
array[50216] <= 16'b0000_0000_0000_0000;
array[50217] <= 16'b0000_0000_0000_0000;
array[50218] <= 16'b0000_0000_0000_0000;
array[50219] <= 16'b0000_0000_0000_0000;
array[50220] <= 16'b0000_0000_0000_0000;
array[50221] <= 16'b0000_0000_0000_0000;
array[50222] <= 16'b0000_0000_0000_0000;
array[50223] <= 16'b0000_0000_0000_0000;
array[50224] <= 16'b0000_0000_0000_0000;
array[50225] <= 16'b0000_0000_0000_0000;
array[50226] <= 16'b0000_0000_0000_0000;
array[50227] <= 16'b0000_0000_0000_0000;
array[50228] <= 16'b0000_0000_0000_0000;
array[50229] <= 16'b0000_0000_0000_0000;
array[50230] <= 16'b0000_0000_0000_0000;
array[50231] <= 16'b0000_0000_0000_0000;
array[50232] <= 16'b0000_0000_0000_0000;
array[50233] <= 16'b0000_0000_0000_0000;
array[50234] <= 16'b0000_0000_0000_0000;
array[50235] <= 16'b0000_0000_0000_0000;
array[50236] <= 16'b0000_0000_0000_0000;
array[50237] <= 16'b0000_0000_0000_0000;
array[50238] <= 16'b0000_0000_0000_0000;
array[50239] <= 16'b0000_0000_0000_0000;
array[50240] <= 16'b0000_0000_0000_0000;
array[50241] <= 16'b0000_0000_0000_0000;
array[50242] <= 16'b0000_0000_0000_0000;
array[50243] <= 16'b0000_0000_0000_0000;
array[50244] <= 16'b0000_0000_0000_0000;
array[50245] <= 16'b0000_0000_0000_0000;
array[50246] <= 16'b0000_0000_0000_0000;
array[50247] <= 16'b0000_0000_0000_0000;
array[50248] <= 16'b0000_0000_0000_0000;
array[50249] <= 16'b0000_0000_0000_0000;
array[50250] <= 16'b0000_0000_0000_0000;
array[50251] <= 16'b0000_0000_0000_0000;
array[50252] <= 16'b0000_0000_0000_0000;
array[50253] <= 16'b0000_0000_0000_0000;
array[50254] <= 16'b0000_0000_0000_0000;
array[50255] <= 16'b0000_0000_0000_0000;
array[50256] <= 16'b0000_0000_0000_0000;
array[50257] <= 16'b0000_0000_0000_0000;
array[50258] <= 16'b0000_0000_0000_0000;
array[50259] <= 16'b0000_0000_0000_0000;
array[50260] <= 16'b0000_0000_0000_0000;
array[50261] <= 16'b0000_0000_0000_0000;
array[50262] <= 16'b0000_0000_0000_0000;
array[50263] <= 16'b0000_0000_0000_0000;
array[50264] <= 16'b0000_0000_0000_0000;
array[50265] <= 16'b0000_0000_0000_0000;
array[50266] <= 16'b0000_0000_0000_0000;
array[50267] <= 16'b0000_0000_0000_0000;
array[50268] <= 16'b0000_0000_0000_0000;
array[50269] <= 16'b0000_0000_0000_0000;
array[50270] <= 16'b0000_0000_0000_0000;
array[50271] <= 16'b0000_0000_0000_0000;
array[50272] <= 16'b0000_0000_0000_0000;
array[50273] <= 16'b0000_0000_0000_0000;
array[50274] <= 16'b0000_0000_0000_0000;
array[50275] <= 16'b0000_0000_0000_0000;
array[50276] <= 16'b0000_0000_0000_0000;
array[50277] <= 16'b0000_0000_0000_0000;
array[50278] <= 16'b0000_0000_0000_0000;
array[50279] <= 16'b0000_0000_0000_0000;
array[50280] <= 16'b0000_0000_0000_0000;
array[50281] <= 16'b0000_0000_0000_0000;
array[50282] <= 16'b0000_0000_0000_0000;
array[50283] <= 16'b0000_0000_0000_0000;
array[50284] <= 16'b0000_0000_0000_0000;
array[50285] <= 16'b0000_0000_0000_0000;
array[50286] <= 16'b0000_0000_0000_0000;
array[50287] <= 16'b0000_0000_0000_0000;
array[50288] <= 16'b0000_0000_0000_0000;
array[50289] <= 16'b0000_0000_0000_0000;
array[50290] <= 16'b0000_0000_0000_0000;
array[50291] <= 16'b0000_0000_0000_0000;
array[50292] <= 16'b0000_0000_0000_0000;
array[50293] <= 16'b0000_0000_0000_0000;
array[50294] <= 16'b0000_0000_0000_0000;
array[50295] <= 16'b0000_0000_0000_0000;
array[50296] <= 16'b0000_0000_0000_0000;
array[50297] <= 16'b0000_0000_0000_0000;
array[50298] <= 16'b0000_0000_0000_0000;
array[50299] <= 16'b0000_0000_0000_0000;
array[50300] <= 16'b0000_0000_0000_0000;
array[50301] <= 16'b0000_0000_0000_0000;
array[50302] <= 16'b0000_0000_0000_0000;
array[50303] <= 16'b0000_0000_0000_0000;
array[50304] <= 16'b0000_0000_0000_0000;
array[50305] <= 16'b0000_0000_0000_0000;
array[50306] <= 16'b0000_0000_0000_0000;
array[50307] <= 16'b0000_0000_0000_0000;
array[50308] <= 16'b0000_0000_0000_0000;
array[50309] <= 16'b0000_0000_0000_0000;
array[50310] <= 16'b0000_0000_0000_0000;
array[50311] <= 16'b0000_0000_0000_0000;
array[50312] <= 16'b0000_0000_0000_0000;
array[50313] <= 16'b0000_0000_0000_0000;
array[50314] <= 16'b0000_0000_0000_0000;
array[50315] <= 16'b0000_0000_0000_0000;
array[50316] <= 16'b0000_0000_0000_0000;
array[50317] <= 16'b0000_0000_0000_0000;
array[50318] <= 16'b0000_0000_0000_0000;
array[50319] <= 16'b0000_0000_0000_0000;
array[50320] <= 16'b0000_0000_0000_0000;
array[50321] <= 16'b0000_0000_0000_0000;
array[50322] <= 16'b0000_0000_0000_0000;
array[50323] <= 16'b0000_0000_0000_0000;
array[50324] <= 16'b0000_0000_0000_0000;
array[50325] <= 16'b0000_0000_0000_0000;
array[50326] <= 16'b0000_0000_0000_0000;
array[50327] <= 16'b0000_0000_0000_0000;
array[50328] <= 16'b0000_0000_0000_0000;
array[50329] <= 16'b0000_0000_0000_0000;
array[50330] <= 16'b0000_0000_0000_0000;
array[50331] <= 16'b0000_0000_0000_0000;
array[50332] <= 16'b0000_0000_0000_0000;
array[50333] <= 16'b0000_0000_0000_0000;
array[50334] <= 16'b0000_0000_0000_0000;
array[50335] <= 16'b0000_0000_0000_0000;
array[50336] <= 16'b0000_0000_0000_0000;
array[50337] <= 16'b0000_0000_0000_0000;
array[50338] <= 16'b0000_0000_0000_0000;
array[50339] <= 16'b0000_0000_0000_0000;
array[50340] <= 16'b0000_0000_0000_0000;
array[50341] <= 16'b0000_0000_0000_0000;
array[50342] <= 16'b0000_0000_0000_0000;
array[50343] <= 16'b0000_0000_0000_0000;
array[50344] <= 16'b0000_0000_0000_0000;
array[50345] <= 16'b0000_0000_0000_0000;
array[50346] <= 16'b0000_0000_0000_0000;
array[50347] <= 16'b0000_0000_0000_0000;
array[50348] <= 16'b0000_0000_0000_0000;
array[50349] <= 16'b0000_0000_0000_0000;
array[50350] <= 16'b0000_0000_0000_0000;
array[50351] <= 16'b0000_0000_0000_0000;
array[50352] <= 16'b0000_0000_0000_0000;
array[50353] <= 16'b0000_0000_0000_0000;
array[50354] <= 16'b0000_0000_0000_0000;
array[50355] <= 16'b0000_0000_0000_0000;
array[50356] <= 16'b0000_0000_0000_0000;
array[50357] <= 16'b0000_0000_0000_0000;
array[50358] <= 16'b0000_0000_0000_0000;
array[50359] <= 16'b0000_0000_0000_0000;
array[50360] <= 16'b0000_0000_0000_0000;
array[50361] <= 16'b0000_0000_0000_0000;
array[50362] <= 16'b0000_0000_0000_0000;
array[50363] <= 16'b0000_0000_0000_0000;
array[50364] <= 16'b0000_0000_0000_0000;
array[50365] <= 16'b0000_0000_0000_0000;
array[50366] <= 16'b0000_0000_0000_0000;
array[50367] <= 16'b0000_0000_0000_0000;
array[50368] <= 16'b0000_0000_0000_0000;
array[50369] <= 16'b0000_0000_0000_0000;
array[50370] <= 16'b0000_0000_0000_0000;
array[50371] <= 16'b0000_0000_0000_0000;
array[50372] <= 16'b0000_0000_0000_0000;
array[50373] <= 16'b0000_0000_0000_0000;
array[50374] <= 16'b0000_0000_0000_0000;
array[50375] <= 16'b0000_0000_0000_0000;
array[50376] <= 16'b0000_0000_0000_0000;
array[50377] <= 16'b0000_0000_0000_0000;
array[50378] <= 16'b0000_0000_0000_0000;
array[50379] <= 16'b0000_0000_0000_0000;
array[50380] <= 16'b0000_0000_0000_0000;
array[50381] <= 16'b0000_0000_0000_0000;
array[50382] <= 16'b0000_0000_0000_0000;
array[50383] <= 16'b0000_0000_0000_0000;
array[50384] <= 16'b0000_0000_0000_0000;
array[50385] <= 16'b0000_0000_0000_0000;
array[50386] <= 16'b0000_0000_0000_0000;
array[50387] <= 16'b0000_0000_0000_0000;
array[50388] <= 16'b0000_0000_0000_0000;
array[50389] <= 16'b0000_0000_0000_0000;
array[50390] <= 16'b0000_0000_0000_0000;
array[50391] <= 16'b0000_0000_0000_0000;
array[50392] <= 16'b0000_0000_0000_0000;
array[50393] <= 16'b0000_0000_0000_0000;
array[50394] <= 16'b0000_0000_0000_0000;
array[50395] <= 16'b0000_0000_0000_0000;
array[50396] <= 16'b0000_0000_0000_0000;
array[50397] <= 16'b0000_0000_0000_0000;
array[50398] <= 16'b0000_0000_0000_0000;
array[50399] <= 16'b0000_0000_0000_0000;
array[50400] <= 16'b0000_0000_0000_0000;
array[50401] <= 16'b0000_0000_0000_0000;
array[50402] <= 16'b0000_0000_0000_0000;
array[50403] <= 16'b0000_0000_0000_0000;
array[50404] <= 16'b0000_0000_0000_0000;
array[50405] <= 16'b0000_0000_0000_0000;
array[50406] <= 16'b0000_0000_0000_0000;
array[50407] <= 16'b0000_0000_0000_0000;
array[50408] <= 16'b0000_0000_0000_0000;
array[50409] <= 16'b0000_0000_0000_0000;
array[50410] <= 16'b0000_0000_0000_0000;
array[50411] <= 16'b0000_0000_0000_0000;
array[50412] <= 16'b0000_0000_0000_0000;
array[50413] <= 16'b0000_0000_0000_0000;
array[50414] <= 16'b0000_0000_0000_0000;
array[50415] <= 16'b0000_0000_0000_0000;
array[50416] <= 16'b0000_0000_0000_0000;
array[50417] <= 16'b0000_0000_0000_0000;
array[50418] <= 16'b0000_0000_0000_0000;
array[50419] <= 16'b0000_0000_0000_0000;
array[50420] <= 16'b0000_0000_0000_0000;
array[50421] <= 16'b0000_0000_0000_0000;
array[50422] <= 16'b0000_0000_0000_0000;
array[50423] <= 16'b0000_0000_0000_0000;
array[50424] <= 16'b0000_0000_0000_0000;
array[50425] <= 16'b0000_0000_0000_0000;
array[50426] <= 16'b0000_0000_0000_0000;
array[50427] <= 16'b0000_0000_0000_0000;
array[50428] <= 16'b0000_0000_0000_0000;
array[50429] <= 16'b0000_0000_0000_0000;
array[50430] <= 16'b0000_0000_0000_0000;
array[50431] <= 16'b0000_0000_0000_0000;
array[50432] <= 16'b0000_0000_0000_0000;
array[50433] <= 16'b0000_0000_0000_0000;
array[50434] <= 16'b0000_0000_0000_0000;
array[50435] <= 16'b0000_0000_0000_0000;
array[50436] <= 16'b0000_0000_0000_0000;
array[50437] <= 16'b0000_0000_0000_0000;
array[50438] <= 16'b0000_0000_0000_0000;
array[50439] <= 16'b0000_0000_0000_0000;
array[50440] <= 16'b0000_0000_0000_0000;
array[50441] <= 16'b0000_0000_0000_0000;
array[50442] <= 16'b0000_0000_0000_0000;
array[50443] <= 16'b0000_0000_0000_0000;
array[50444] <= 16'b0000_0000_0000_0000;
array[50445] <= 16'b0000_0000_0000_0000;
array[50446] <= 16'b0000_0000_0000_0000;
array[50447] <= 16'b0000_0000_0000_0000;
array[50448] <= 16'b0000_0000_0000_0000;
array[50449] <= 16'b0000_0000_0000_0000;
array[50450] <= 16'b0000_0000_0000_0000;
array[50451] <= 16'b0000_0000_0000_0000;
array[50452] <= 16'b0000_0000_0000_0000;
array[50453] <= 16'b0000_0000_0000_0000;
array[50454] <= 16'b0000_0000_0000_0000;
array[50455] <= 16'b0000_0000_0000_0000;
array[50456] <= 16'b0000_0000_0000_0000;
array[50457] <= 16'b0000_0000_0000_0000;
array[50458] <= 16'b0000_0000_0000_0000;
array[50459] <= 16'b0000_0000_0000_0000;
array[50460] <= 16'b0000_0000_0000_0000;
array[50461] <= 16'b0000_0000_0000_0000;
array[50462] <= 16'b0000_0000_0000_0000;
array[50463] <= 16'b0000_0000_0000_0000;
array[50464] <= 16'b0000_0000_0000_0000;
array[50465] <= 16'b0000_0000_0000_0000;
array[50466] <= 16'b0000_0000_0000_0000;
array[50467] <= 16'b0000_0000_0000_0000;
array[50468] <= 16'b0000_0000_0000_0000;
array[50469] <= 16'b0000_0000_0000_0000;
array[50470] <= 16'b0000_0000_0000_0000;
array[50471] <= 16'b0000_0000_0000_0000;
array[50472] <= 16'b0000_0000_0000_0000;
array[50473] <= 16'b0000_0000_0000_0000;
array[50474] <= 16'b0000_0000_0000_0000;
array[50475] <= 16'b0000_0000_0000_0000;
array[50476] <= 16'b0000_0000_0000_0000;
array[50477] <= 16'b0000_0000_0000_0000;
array[50478] <= 16'b0000_0000_0000_0000;
array[50479] <= 16'b0000_0000_0000_0000;
array[50480] <= 16'b0000_0000_0000_0000;
array[50481] <= 16'b0000_0000_0000_0000;
array[50482] <= 16'b0000_0000_0000_0000;
array[50483] <= 16'b0000_0000_0000_0000;
array[50484] <= 16'b0000_0000_0000_0000;
array[50485] <= 16'b0000_0000_0000_0000;
array[50486] <= 16'b0000_0000_0000_0000;
array[50487] <= 16'b0000_0000_0000_0000;
array[50488] <= 16'b0000_0000_0000_0000;
array[50489] <= 16'b0000_0000_0000_0000;
array[50490] <= 16'b0000_0000_0000_0000;
array[50491] <= 16'b0000_0000_0000_0000;
array[50492] <= 16'b0000_0000_0000_0000;
array[50493] <= 16'b0000_0000_0000_0000;
array[50494] <= 16'b0000_0000_0000_0000;
array[50495] <= 16'b0000_0000_0000_0000;
array[50496] <= 16'b0000_0000_0000_0000;
array[50497] <= 16'b0000_0000_0000_0000;
array[50498] <= 16'b0000_0000_0000_0000;
array[50499] <= 16'b0000_0000_0000_0000;
array[50500] <= 16'b0000_0000_0000_0000;
array[50501] <= 16'b0000_0000_0000_0000;
array[50502] <= 16'b0000_0000_0000_0000;
array[50503] <= 16'b0000_0000_0000_0000;
array[50504] <= 16'b0000_0000_0000_0000;
array[50505] <= 16'b0000_0000_0000_0000;
array[50506] <= 16'b0000_0000_0000_0000;
array[50507] <= 16'b0000_0000_0000_0000;
array[50508] <= 16'b0000_0000_0000_0000;
array[50509] <= 16'b0000_0000_0000_0000;
array[50510] <= 16'b0000_0000_0000_0000;
array[50511] <= 16'b0000_0000_0000_0000;
array[50512] <= 16'b0000_0000_0000_0000;
array[50513] <= 16'b0000_0000_0000_0000;
array[50514] <= 16'b0000_0000_0000_0000;
array[50515] <= 16'b0000_0000_0000_0000;
array[50516] <= 16'b0000_0000_0000_0000;
array[50517] <= 16'b0000_0000_0000_0000;
array[50518] <= 16'b0000_0000_0000_0000;
array[50519] <= 16'b0000_0000_0000_0000;
array[50520] <= 16'b0000_0000_0000_0000;
array[50521] <= 16'b0000_0000_0000_0000;
array[50522] <= 16'b0000_0000_0000_0000;
array[50523] <= 16'b0000_0000_0000_0000;
array[50524] <= 16'b0000_0000_0000_0000;
array[50525] <= 16'b0000_0000_0000_0000;
array[50526] <= 16'b0000_0000_0000_0000;
array[50527] <= 16'b0000_0000_0000_0000;
array[50528] <= 16'b0000_0000_0000_0000;
array[50529] <= 16'b0000_0000_0000_0000;
array[50530] <= 16'b0000_0000_0000_0000;
array[50531] <= 16'b0000_0000_0000_0000;
array[50532] <= 16'b0000_0000_0000_0000;
array[50533] <= 16'b0000_0000_0000_0000;
array[50534] <= 16'b0000_0000_0000_0000;
array[50535] <= 16'b0000_0000_0000_0000;
array[50536] <= 16'b0000_0000_0000_0000;
array[50537] <= 16'b0000_0000_0000_0000;
array[50538] <= 16'b0000_0000_0000_0000;
array[50539] <= 16'b0000_0000_0000_0000;
array[50540] <= 16'b0000_0000_0000_0000;
array[50541] <= 16'b0000_0000_0000_0000;
array[50542] <= 16'b0000_0000_0000_0000;
array[50543] <= 16'b0000_0000_0000_0000;
array[50544] <= 16'b0000_0000_0000_0000;
array[50545] <= 16'b0000_0000_0000_0000;
array[50546] <= 16'b0000_0000_0000_0000;
array[50547] <= 16'b0000_0000_0000_0000;
array[50548] <= 16'b0000_0000_0000_0000;
array[50549] <= 16'b0000_0000_0000_0000;
array[50550] <= 16'b0000_0000_0000_0000;
array[50551] <= 16'b0000_0000_0000_0000;
array[50552] <= 16'b0000_0000_0000_0000;
array[50553] <= 16'b0000_0000_0000_0000;
array[50554] <= 16'b0000_0000_0000_0000;
array[50555] <= 16'b0000_0000_0000_0000;
array[50556] <= 16'b0000_0000_0000_0000;
array[50557] <= 16'b0000_0000_0000_0000;
array[50558] <= 16'b0000_0000_0000_0000;
array[50559] <= 16'b0000_0000_0000_0000;
array[50560] <= 16'b0000_0000_0000_0000;
array[50561] <= 16'b0000_0000_0000_0000;
array[50562] <= 16'b0000_0000_0000_0000;
array[50563] <= 16'b0000_0000_0000_0000;
array[50564] <= 16'b0000_0000_0000_0000;
array[50565] <= 16'b0000_0000_0000_0000;
array[50566] <= 16'b0000_0000_0000_0000;
array[50567] <= 16'b0000_0000_0000_0000;
array[50568] <= 16'b0000_0000_0000_0000;
array[50569] <= 16'b0000_0000_0000_0000;
array[50570] <= 16'b0000_0000_0000_0000;
array[50571] <= 16'b0000_0000_0000_0000;
array[50572] <= 16'b0000_0000_0000_0000;
array[50573] <= 16'b0000_0000_0000_0000;
array[50574] <= 16'b0000_0000_0000_0000;
array[50575] <= 16'b0000_0000_0000_0000;
array[50576] <= 16'b0000_0000_0000_0000;
array[50577] <= 16'b0000_0000_0000_0000;
array[50578] <= 16'b0000_0000_0000_0000;
array[50579] <= 16'b0000_0000_0000_0000;
array[50580] <= 16'b0000_0000_0000_0000;
array[50581] <= 16'b0000_0000_0000_0000;
array[50582] <= 16'b0000_0000_0000_0000;
array[50583] <= 16'b0000_0000_0000_0000;
array[50584] <= 16'b0000_0000_0000_0000;
array[50585] <= 16'b0000_0000_0000_0000;
array[50586] <= 16'b0000_0000_0000_0000;
array[50587] <= 16'b0000_0000_0000_0000;
array[50588] <= 16'b0000_0000_0000_0000;
array[50589] <= 16'b0000_0000_0000_0000;
array[50590] <= 16'b0000_0000_0000_0000;
array[50591] <= 16'b0000_0000_0000_0000;
array[50592] <= 16'b0000_0000_0000_0000;
array[50593] <= 16'b0000_0000_0000_0000;
array[50594] <= 16'b0000_0000_0000_0000;
array[50595] <= 16'b0000_0000_0000_0000;
array[50596] <= 16'b0000_0000_0000_0000;
array[50597] <= 16'b0000_0000_0000_0000;
array[50598] <= 16'b0000_0000_0000_0000;
array[50599] <= 16'b0000_0000_0000_0000;
array[50600] <= 16'b0000_0000_0000_0000;
array[50601] <= 16'b0000_0000_0000_0000;
array[50602] <= 16'b0000_0000_0000_0000;
array[50603] <= 16'b0000_0000_0000_0000;
array[50604] <= 16'b0000_0000_0000_0000;
array[50605] <= 16'b0000_0000_0000_0000;
array[50606] <= 16'b0000_0000_0000_0000;
array[50607] <= 16'b0000_0000_0000_0000;
array[50608] <= 16'b0000_0000_0000_0000;
array[50609] <= 16'b0000_0000_0000_0000;
array[50610] <= 16'b0000_0000_0000_0000;
array[50611] <= 16'b0000_0000_0000_0000;
array[50612] <= 16'b0000_0000_0000_0000;
array[50613] <= 16'b0000_0000_0000_0000;
array[50614] <= 16'b0000_0000_0000_0000;
array[50615] <= 16'b0000_0000_0000_0000;
array[50616] <= 16'b0000_0000_0000_0000;
array[50617] <= 16'b0000_0000_0000_0000;
array[50618] <= 16'b0000_0000_0000_0000;
array[50619] <= 16'b0000_0000_0000_0000;
array[50620] <= 16'b0000_0000_0000_0000;
array[50621] <= 16'b0000_0000_0000_0000;
array[50622] <= 16'b0000_0000_0000_0000;
array[50623] <= 16'b0000_0000_0000_0000;
array[50624] <= 16'b0000_0000_0000_0000;
array[50625] <= 16'b0000_0000_0000_0000;
array[50626] <= 16'b0000_0000_0000_0000;
array[50627] <= 16'b0000_0000_0000_0000;
array[50628] <= 16'b0000_0000_0000_0000;
array[50629] <= 16'b0000_0000_0000_0000;
array[50630] <= 16'b0000_0000_0000_0000;
array[50631] <= 16'b0000_0000_0000_0000;
array[50632] <= 16'b0000_0000_0000_0000;
array[50633] <= 16'b0000_0000_0000_0000;
array[50634] <= 16'b0000_0000_0000_0000;
array[50635] <= 16'b0000_0000_0000_0000;
array[50636] <= 16'b0000_0000_0000_0000;
array[50637] <= 16'b0000_0000_0000_0000;
array[50638] <= 16'b0000_0000_0000_0000;
array[50639] <= 16'b0000_0000_0000_0000;
array[50640] <= 16'b0000_0000_0000_0000;
array[50641] <= 16'b0000_0000_0000_0000;
array[50642] <= 16'b0000_0000_0000_0000;
array[50643] <= 16'b0000_0000_0000_0000;
array[50644] <= 16'b0000_0000_0000_0000;
array[50645] <= 16'b0000_0000_0000_0000;
array[50646] <= 16'b0000_0000_0000_0000;
array[50647] <= 16'b0000_0000_0000_0000;
array[50648] <= 16'b0000_0000_0000_0000;
array[50649] <= 16'b0000_0000_0000_0000;
array[50650] <= 16'b0000_0000_0000_0000;
array[50651] <= 16'b0000_0000_0000_0000;
array[50652] <= 16'b0000_0000_0000_0000;
array[50653] <= 16'b0000_0000_0000_0000;
array[50654] <= 16'b0000_0000_0000_0000;
array[50655] <= 16'b0000_0000_0000_0000;
array[50656] <= 16'b0000_0000_0000_0000;
array[50657] <= 16'b0000_0000_0000_0000;
array[50658] <= 16'b0000_0000_0000_0000;
array[50659] <= 16'b0000_0000_0000_0000;
array[50660] <= 16'b0000_0000_0000_0000;
array[50661] <= 16'b0000_0000_0000_0000;
array[50662] <= 16'b0000_0000_0000_0000;
array[50663] <= 16'b0000_0000_0000_0000;
array[50664] <= 16'b0000_0000_0000_0000;
array[50665] <= 16'b0000_0000_0000_0000;
array[50666] <= 16'b0000_0000_0000_0000;
array[50667] <= 16'b0000_0000_0000_0000;
array[50668] <= 16'b0000_0000_0000_0000;
array[50669] <= 16'b0000_0000_0000_0000;
array[50670] <= 16'b0000_0000_0000_0000;
array[50671] <= 16'b0000_0000_0000_0000;
array[50672] <= 16'b0000_0000_0000_0000;
array[50673] <= 16'b0000_0000_0000_0000;
array[50674] <= 16'b0000_0000_0000_0000;
array[50675] <= 16'b0000_0000_0000_0000;
array[50676] <= 16'b0000_0000_0000_0000;
array[50677] <= 16'b0000_0000_0000_0000;
array[50678] <= 16'b0000_0000_0000_0000;
array[50679] <= 16'b0000_0000_0000_0000;
array[50680] <= 16'b0000_0000_0000_0000;
array[50681] <= 16'b0000_0000_0000_0000;
array[50682] <= 16'b0000_0000_0000_0000;
array[50683] <= 16'b0000_0000_0000_0000;
array[50684] <= 16'b0000_0000_0000_0000;
array[50685] <= 16'b0000_0000_0000_0000;
array[50686] <= 16'b0000_0000_0000_0000;
array[50687] <= 16'b0000_0000_0000_0000;
array[50688] <= 16'b0000_0000_0000_0000;
array[50689] <= 16'b0000_0000_0000_0000;
array[50690] <= 16'b0000_0000_0000_0000;
array[50691] <= 16'b0000_0000_0000_0000;
array[50692] <= 16'b0000_0000_0000_0000;
array[50693] <= 16'b0000_0000_0000_0000;
array[50694] <= 16'b0000_0000_0000_0000;
array[50695] <= 16'b0000_0000_0000_0000;
array[50696] <= 16'b0000_0000_0000_0000;
array[50697] <= 16'b0000_0000_0000_0000;
array[50698] <= 16'b0000_0000_0000_0000;
array[50699] <= 16'b0000_0000_0000_0000;
array[50700] <= 16'b0000_0000_0000_0000;
array[50701] <= 16'b0000_0000_0000_0000;
array[50702] <= 16'b0000_0000_0000_0000;
array[50703] <= 16'b0000_0000_0000_0000;
array[50704] <= 16'b0000_0000_0000_0000;
array[50705] <= 16'b0000_0000_0000_0000;
array[50706] <= 16'b0000_0000_0000_0000;
array[50707] <= 16'b0000_0000_0000_0000;
array[50708] <= 16'b0000_0000_0000_0000;
array[50709] <= 16'b0000_0000_0000_0000;
array[50710] <= 16'b0000_0000_0000_0000;
array[50711] <= 16'b0000_0000_0000_0000;
array[50712] <= 16'b0000_0000_0000_0000;
array[50713] <= 16'b0000_0000_0000_0000;
array[50714] <= 16'b0000_0000_0000_0000;
array[50715] <= 16'b0000_0000_0000_0000;
array[50716] <= 16'b0000_0000_0000_0000;
array[50717] <= 16'b0000_0000_0000_0000;
array[50718] <= 16'b0000_0000_0000_0000;
array[50719] <= 16'b0000_0000_0000_0000;
array[50720] <= 16'b0000_0000_0000_0000;
array[50721] <= 16'b0000_0000_0000_0000;
array[50722] <= 16'b0000_0000_0000_0000;
array[50723] <= 16'b0000_0000_0000_0000;
array[50724] <= 16'b0000_0000_0000_0000;
array[50725] <= 16'b0000_0000_0000_0000;
array[50726] <= 16'b0000_0000_0000_0000;
array[50727] <= 16'b0000_0000_0000_0000;
array[50728] <= 16'b0000_0000_0000_0000;
array[50729] <= 16'b0000_0000_0000_0000;
array[50730] <= 16'b0000_0000_0000_0000;
array[50731] <= 16'b0000_0000_0000_0000;
array[50732] <= 16'b0000_0000_0000_0000;
array[50733] <= 16'b0000_0000_0000_0000;
array[50734] <= 16'b0000_0000_0000_0000;
array[50735] <= 16'b0000_0000_0000_0000;
array[50736] <= 16'b0000_0000_0000_0000;
array[50737] <= 16'b0000_0000_0000_0000;
array[50738] <= 16'b0000_0000_0000_0000;
array[50739] <= 16'b0000_0000_0000_0000;
array[50740] <= 16'b0000_0000_0000_0000;
array[50741] <= 16'b0000_0000_0000_0000;
array[50742] <= 16'b0000_0000_0000_0000;
array[50743] <= 16'b0000_0000_0000_0000;
array[50744] <= 16'b0000_0000_0000_0000;
array[50745] <= 16'b0000_0000_0000_0000;
array[50746] <= 16'b0000_0000_0000_0000;
array[50747] <= 16'b0000_0000_0000_0000;
array[50748] <= 16'b0000_0000_0000_0000;
array[50749] <= 16'b0000_0000_0000_0000;
array[50750] <= 16'b0000_0000_0000_0000;
array[50751] <= 16'b0000_0000_0000_0000;
array[50752] <= 16'b0000_0000_0000_0000;
array[50753] <= 16'b0000_0000_0000_0000;
array[50754] <= 16'b0000_0000_0000_0000;
array[50755] <= 16'b0000_0000_0000_0000;
array[50756] <= 16'b0000_0000_0000_0000;
array[50757] <= 16'b0000_0000_0000_0000;
array[50758] <= 16'b0000_0000_0000_0000;
array[50759] <= 16'b0000_0000_0000_0000;
array[50760] <= 16'b0000_0000_0000_0000;
array[50761] <= 16'b0000_0000_0000_0000;
array[50762] <= 16'b0000_0000_0000_0000;
array[50763] <= 16'b0000_0000_0000_0000;
array[50764] <= 16'b0000_0000_0000_0000;
array[50765] <= 16'b0000_0000_0000_0000;
array[50766] <= 16'b0000_0000_0000_0000;
array[50767] <= 16'b0000_0000_0000_0000;
array[50768] <= 16'b0000_0000_0000_0000;
array[50769] <= 16'b0000_0000_0000_0000;
array[50770] <= 16'b0000_0000_0000_0000;
array[50771] <= 16'b0000_0000_0000_0000;
array[50772] <= 16'b0000_0000_0000_0000;
array[50773] <= 16'b0000_0000_0000_0000;
array[50774] <= 16'b0000_0000_0000_0000;
array[50775] <= 16'b0000_0000_0000_0000;
array[50776] <= 16'b0000_0000_0000_0000;
array[50777] <= 16'b0000_0000_0000_0000;
array[50778] <= 16'b0000_0000_0000_0000;
array[50779] <= 16'b0000_0000_0000_0000;
array[50780] <= 16'b0000_0000_0000_0000;
array[50781] <= 16'b0000_0000_0000_0000;
array[50782] <= 16'b0000_0000_0000_0000;
array[50783] <= 16'b0000_0000_0000_0000;
array[50784] <= 16'b0000_0000_0000_0000;
array[50785] <= 16'b0000_0000_0000_0000;
array[50786] <= 16'b0000_0000_0000_0000;
array[50787] <= 16'b0000_0000_0000_0000;
array[50788] <= 16'b0000_0000_0000_0000;
array[50789] <= 16'b0000_0000_0000_0000;
array[50790] <= 16'b0000_0000_0000_0000;
array[50791] <= 16'b0000_0000_0000_0000;
array[50792] <= 16'b0000_0000_0000_0000;
array[50793] <= 16'b0000_0000_0000_0000;
array[50794] <= 16'b0000_0000_0000_0000;
array[50795] <= 16'b0000_0000_0000_0000;
array[50796] <= 16'b0000_0000_0000_0000;
array[50797] <= 16'b0000_0000_0000_0000;
array[50798] <= 16'b0000_0000_0000_0000;
array[50799] <= 16'b0000_0000_0000_0000;
array[50800] <= 16'b0000_0000_0000_0000;
array[50801] <= 16'b0000_0000_0000_0000;
array[50802] <= 16'b0000_0000_0000_0000;
array[50803] <= 16'b0000_0000_0000_0000;
array[50804] <= 16'b0000_0000_0000_0000;
array[50805] <= 16'b0000_0000_0000_0000;
array[50806] <= 16'b0000_0000_0000_0000;
array[50807] <= 16'b0000_0000_0000_0000;
array[50808] <= 16'b0000_0000_0000_0000;
array[50809] <= 16'b0000_0000_0000_0000;
array[50810] <= 16'b0000_0000_0000_0000;
array[50811] <= 16'b0000_0000_0000_0000;
array[50812] <= 16'b0000_0000_0000_0000;
array[50813] <= 16'b0000_0000_0000_0000;
array[50814] <= 16'b0000_0000_0000_0000;
array[50815] <= 16'b0000_0000_0000_0000;
array[50816] <= 16'b0000_0000_0000_0000;
array[50817] <= 16'b0000_0000_0000_0000;
array[50818] <= 16'b0000_0000_0000_0000;
array[50819] <= 16'b0000_0000_0000_0000;
array[50820] <= 16'b0000_0000_0000_0000;
array[50821] <= 16'b0000_0000_0000_0000;
array[50822] <= 16'b0000_0000_0000_0000;
array[50823] <= 16'b0000_0000_0000_0000;
array[50824] <= 16'b0000_0000_0000_0000;
array[50825] <= 16'b0000_0000_0000_0000;
array[50826] <= 16'b0000_0000_0000_0000;
array[50827] <= 16'b0000_0000_0000_0000;
array[50828] <= 16'b0000_0000_0000_0000;
array[50829] <= 16'b0000_0000_0000_0000;
array[50830] <= 16'b0000_0000_0000_0000;
array[50831] <= 16'b0000_0000_0000_0000;
array[50832] <= 16'b0000_0000_0000_0000;
array[50833] <= 16'b0000_0000_0000_0000;
array[50834] <= 16'b0000_0000_0000_0000;
array[50835] <= 16'b0000_0000_0000_0000;
array[50836] <= 16'b0000_0000_0000_0000;
array[50837] <= 16'b0000_0000_0000_0000;
array[50838] <= 16'b0000_0000_0000_0000;
array[50839] <= 16'b0000_0000_0000_0000;
array[50840] <= 16'b0000_0000_0000_0000;
array[50841] <= 16'b0000_0000_0000_0000;
array[50842] <= 16'b0000_0000_0000_0000;
array[50843] <= 16'b0000_0000_0000_0000;
array[50844] <= 16'b0000_0000_0000_0000;
array[50845] <= 16'b0000_0000_0000_0000;
array[50846] <= 16'b0000_0000_0000_0000;
array[50847] <= 16'b0000_0000_0000_0000;
array[50848] <= 16'b0000_0000_0000_0000;
array[50849] <= 16'b0000_0000_0000_0000;
array[50850] <= 16'b0000_0000_0000_0000;
array[50851] <= 16'b0000_0000_0000_0000;
array[50852] <= 16'b0000_0000_0000_0000;
array[50853] <= 16'b0000_0000_0000_0000;
array[50854] <= 16'b0000_0000_0000_0000;
array[50855] <= 16'b0000_0000_0000_0000;
array[50856] <= 16'b0000_0000_0000_0000;
array[50857] <= 16'b0000_0000_0000_0000;
array[50858] <= 16'b0000_0000_0000_0000;
array[50859] <= 16'b0000_0000_0000_0000;
array[50860] <= 16'b0000_0000_0000_0000;
array[50861] <= 16'b0000_0000_0000_0000;
array[50862] <= 16'b0000_0000_0000_0000;
array[50863] <= 16'b0000_0000_0000_0000;
array[50864] <= 16'b0000_0000_0000_0000;
array[50865] <= 16'b0000_0000_0000_0000;
array[50866] <= 16'b0000_0000_0000_0000;
array[50867] <= 16'b0000_0000_0000_0000;
array[50868] <= 16'b0000_0000_0000_0000;
array[50869] <= 16'b0000_0000_0000_0000;
array[50870] <= 16'b0000_0000_0000_0000;
array[50871] <= 16'b0000_0000_0000_0000;
array[50872] <= 16'b0000_0000_0000_0000;
array[50873] <= 16'b0000_0000_0000_0000;
array[50874] <= 16'b0000_0000_0000_0000;
array[50875] <= 16'b0000_0000_0000_0000;
array[50876] <= 16'b0000_0000_0000_0000;
array[50877] <= 16'b0000_0000_0000_0000;
array[50878] <= 16'b0000_0000_0000_0000;
array[50879] <= 16'b0000_0000_0000_0000;
array[50880] <= 16'b0000_0000_0000_0000;
array[50881] <= 16'b0000_0000_0000_0000;
array[50882] <= 16'b0000_0000_0000_0000;
array[50883] <= 16'b0000_0000_0000_0000;
array[50884] <= 16'b0000_0000_0000_0000;
array[50885] <= 16'b0000_0000_0000_0000;
array[50886] <= 16'b0000_0000_0000_0000;
array[50887] <= 16'b0000_0000_0000_0000;
array[50888] <= 16'b0000_0000_0000_0000;
array[50889] <= 16'b0000_0000_0000_0000;
array[50890] <= 16'b0000_0000_0000_0000;
array[50891] <= 16'b0000_0000_0000_0000;
array[50892] <= 16'b0000_0000_0000_0000;
array[50893] <= 16'b0000_0000_0000_0000;
array[50894] <= 16'b0000_0000_0000_0000;
array[50895] <= 16'b0000_0000_0000_0000;
array[50896] <= 16'b0000_0000_0000_0000;
array[50897] <= 16'b0000_0000_0000_0000;
array[50898] <= 16'b0000_0000_0000_0000;
array[50899] <= 16'b0000_0000_0000_0000;
array[50900] <= 16'b0000_0000_0000_0000;
array[50901] <= 16'b0000_0000_0000_0000;
array[50902] <= 16'b0000_0000_0000_0000;
array[50903] <= 16'b0000_0000_0000_0000;
array[50904] <= 16'b0000_0000_0000_0000;
array[50905] <= 16'b0000_0000_0000_0000;
array[50906] <= 16'b0000_0000_0000_0000;
array[50907] <= 16'b0000_0000_0000_0000;
array[50908] <= 16'b0000_0000_0000_0000;
array[50909] <= 16'b0000_0000_0000_0000;
array[50910] <= 16'b0000_0000_0000_0000;
array[50911] <= 16'b0000_0000_0000_0000;
array[50912] <= 16'b0000_0000_0000_0000;
array[50913] <= 16'b0000_0000_0000_0000;
array[50914] <= 16'b0000_0000_0000_0000;
array[50915] <= 16'b0000_0000_0000_0000;
array[50916] <= 16'b0000_0000_0000_0000;
array[50917] <= 16'b0000_0000_0000_0000;
array[50918] <= 16'b0000_0000_0000_0000;
array[50919] <= 16'b0000_0000_0000_0000;
array[50920] <= 16'b0000_0000_0000_0000;
array[50921] <= 16'b0000_0000_0000_0000;
array[50922] <= 16'b0000_0000_0000_0000;
array[50923] <= 16'b0000_0000_0000_0000;
array[50924] <= 16'b0000_0000_0000_0000;
array[50925] <= 16'b0000_0000_0000_0000;
array[50926] <= 16'b0000_0000_0000_0000;
array[50927] <= 16'b0000_0000_0000_0000;
array[50928] <= 16'b0000_0000_0000_0000;
array[50929] <= 16'b0000_0000_0000_0000;
array[50930] <= 16'b0000_0000_0000_0000;
array[50931] <= 16'b0000_0000_0000_0000;
array[50932] <= 16'b0000_0000_0000_0000;
array[50933] <= 16'b0000_0000_0000_0000;
array[50934] <= 16'b0000_0000_0000_0000;
array[50935] <= 16'b0000_0000_0000_0000;
array[50936] <= 16'b0000_0000_0000_0000;
array[50937] <= 16'b0000_0000_0000_0000;
array[50938] <= 16'b0000_0000_0000_0000;
array[50939] <= 16'b0000_0000_0000_0000;
array[50940] <= 16'b0000_0000_0000_0000;
array[50941] <= 16'b0000_0000_0000_0000;
array[50942] <= 16'b0000_0000_0000_0000;
array[50943] <= 16'b0000_0000_0000_0000;
array[50944] <= 16'b0000_0000_0000_0000;
array[50945] <= 16'b0000_0000_0000_0000;
array[50946] <= 16'b0000_0000_0000_0000;
array[50947] <= 16'b0000_0000_0000_0000;
array[50948] <= 16'b0000_0000_0000_0000;
array[50949] <= 16'b0000_0000_0000_0000;
array[50950] <= 16'b0000_0000_0000_0000;
array[50951] <= 16'b0000_0000_0000_0000;
array[50952] <= 16'b0000_0000_0000_0000;
array[50953] <= 16'b0000_0000_0000_0000;
array[50954] <= 16'b0000_0000_0000_0000;
array[50955] <= 16'b0000_0000_0000_0000;
array[50956] <= 16'b0000_0000_0000_0000;
array[50957] <= 16'b0000_0000_0000_0000;
array[50958] <= 16'b0000_0000_0000_0000;
array[50959] <= 16'b0000_0000_0000_0000;
array[50960] <= 16'b0000_0000_0000_0000;
array[50961] <= 16'b0000_0000_0000_0000;
array[50962] <= 16'b0000_0000_0000_0000;
array[50963] <= 16'b0000_0000_0000_0000;
array[50964] <= 16'b0000_0000_0000_0000;
array[50965] <= 16'b0000_0000_0000_0000;
array[50966] <= 16'b0000_0000_0000_0000;
array[50967] <= 16'b0000_0000_0000_0000;
array[50968] <= 16'b0000_0000_0000_0000;
array[50969] <= 16'b0000_0000_0000_0000;
array[50970] <= 16'b0000_0000_0000_0000;
array[50971] <= 16'b0000_0000_0000_0000;
array[50972] <= 16'b0000_0000_0000_0000;
array[50973] <= 16'b0000_0000_0000_0000;
array[50974] <= 16'b0000_0000_0000_0000;
array[50975] <= 16'b0000_0000_0000_0000;
array[50976] <= 16'b0000_0000_0000_0000;
array[50977] <= 16'b0000_0000_0000_0000;
array[50978] <= 16'b0000_0000_0000_0000;
array[50979] <= 16'b0000_0000_0000_0000;
array[50980] <= 16'b0000_0000_0000_0000;
array[50981] <= 16'b0000_0000_0000_0000;
array[50982] <= 16'b0000_0000_0000_0000;
array[50983] <= 16'b0000_0000_0000_0000;
array[50984] <= 16'b0000_0000_0000_0000;
array[50985] <= 16'b0000_0000_0000_0000;
array[50986] <= 16'b0000_0000_0000_0000;
array[50987] <= 16'b0000_0000_0000_0000;
array[50988] <= 16'b0000_0000_0000_0000;
array[50989] <= 16'b0000_0000_0000_0000;
array[50990] <= 16'b0000_0000_0000_0000;
array[50991] <= 16'b0000_0000_0000_0000;
array[50992] <= 16'b0000_0000_0000_0000;
array[50993] <= 16'b0000_0000_0000_0000;
array[50994] <= 16'b0000_0000_0000_0000;
array[50995] <= 16'b0000_0000_0000_0000;
array[50996] <= 16'b0000_0000_0000_0000;
array[50997] <= 16'b0000_0000_0000_0000;
array[50998] <= 16'b0000_0000_0000_0000;
array[50999] <= 16'b0000_0000_0000_0000;
array[51000] <= 16'b0000_0000_0000_0000;
array[51001] <= 16'b0000_0000_0000_0000;
array[51002] <= 16'b0000_0000_0000_0000;
array[51003] <= 16'b0000_0000_0000_0000;
array[51004] <= 16'b0000_0000_0000_0000;
array[51005] <= 16'b0000_0000_0000_0000;
array[51006] <= 16'b0000_0000_0000_0000;
array[51007] <= 16'b0000_0000_0000_0000;
array[51008] <= 16'b0000_0000_0000_0000;
array[51009] <= 16'b0000_0000_0000_0000;
array[51010] <= 16'b0000_0000_0000_0000;
array[51011] <= 16'b0000_0000_0000_0000;
array[51012] <= 16'b0000_0000_0000_0000;
array[51013] <= 16'b0000_0000_0000_0000;
array[51014] <= 16'b0000_0000_0000_0000;
array[51015] <= 16'b0000_0000_0000_0000;
array[51016] <= 16'b0000_0000_0000_0000;
array[51017] <= 16'b0000_0000_0000_0000;
array[51018] <= 16'b0000_0000_0000_0000;
array[51019] <= 16'b0000_0000_0000_0000;
array[51020] <= 16'b0000_0000_0000_0000;
array[51021] <= 16'b0000_0000_0000_0000;
array[51022] <= 16'b0000_0000_0000_0000;
array[51023] <= 16'b0000_0000_0000_0000;
array[51024] <= 16'b0000_0000_0000_0000;
array[51025] <= 16'b0000_0000_0000_0000;
array[51026] <= 16'b0000_0000_0000_0000;
array[51027] <= 16'b0000_0000_0000_0000;
array[51028] <= 16'b0000_0000_0000_0000;
array[51029] <= 16'b0000_0000_0000_0000;
array[51030] <= 16'b0000_0000_0000_0000;
array[51031] <= 16'b0000_0000_0000_0000;
array[51032] <= 16'b0000_0000_0000_0000;
array[51033] <= 16'b0000_0000_0000_0000;
array[51034] <= 16'b0000_0000_0000_0000;
array[51035] <= 16'b0000_0000_0000_0000;
array[51036] <= 16'b0000_0000_0000_0000;
array[51037] <= 16'b0000_0000_0000_0000;
array[51038] <= 16'b0000_0000_0000_0000;
array[51039] <= 16'b0000_0000_0000_0000;
array[51040] <= 16'b0000_0000_0000_0000;
array[51041] <= 16'b0000_0000_0000_0000;
array[51042] <= 16'b0000_0000_0000_0000;
array[51043] <= 16'b0000_0000_0000_0000;
array[51044] <= 16'b0000_0000_0000_0000;
array[51045] <= 16'b0000_0000_0000_0000;
array[51046] <= 16'b0000_0000_0000_0000;
array[51047] <= 16'b0000_0000_0000_0000;
array[51048] <= 16'b0000_0000_0000_0000;
array[51049] <= 16'b0000_0000_0000_0000;
array[51050] <= 16'b0000_0000_0000_0000;
array[51051] <= 16'b0000_0000_0000_0000;
array[51052] <= 16'b0000_0000_0000_0000;
array[51053] <= 16'b0000_0000_0000_0000;
array[51054] <= 16'b0000_0000_0000_0000;
array[51055] <= 16'b0000_0000_0000_0000;
array[51056] <= 16'b0000_0000_0000_0000;
array[51057] <= 16'b0000_0000_0000_0000;
array[51058] <= 16'b0000_0000_0000_0000;
array[51059] <= 16'b0000_0000_0000_0000;
array[51060] <= 16'b0000_0000_0000_0000;
array[51061] <= 16'b0000_0000_0000_0000;
array[51062] <= 16'b0000_0000_0000_0000;
array[51063] <= 16'b0000_0000_0000_0000;
array[51064] <= 16'b0000_0000_0000_0000;
array[51065] <= 16'b0000_0000_0000_0000;
array[51066] <= 16'b0000_0000_0000_0000;
array[51067] <= 16'b0000_0000_0000_0000;
array[51068] <= 16'b0000_0000_0000_0000;
array[51069] <= 16'b0000_0000_0000_0000;
array[51070] <= 16'b0000_0000_0000_0000;
array[51071] <= 16'b0000_0000_0000_0000;
array[51072] <= 16'b0000_0000_0000_0000;
array[51073] <= 16'b0000_0000_0000_0000;
array[51074] <= 16'b0000_0000_0000_0000;
array[51075] <= 16'b0000_0000_0000_0000;
array[51076] <= 16'b0000_0000_0000_0000;
array[51077] <= 16'b0000_0000_0000_0000;
array[51078] <= 16'b0000_0000_0000_0000;
array[51079] <= 16'b0000_0000_0000_0000;
array[51080] <= 16'b0000_0000_0000_0000;
array[51081] <= 16'b0000_0000_0000_0000;
array[51082] <= 16'b0000_0000_0000_0000;
array[51083] <= 16'b0000_0000_0000_0000;
array[51084] <= 16'b0000_0000_0000_0000;
array[51085] <= 16'b0000_0000_0000_0000;
array[51086] <= 16'b0000_0000_0000_0000;
array[51087] <= 16'b0000_0000_0000_0000;
array[51088] <= 16'b0000_0000_0000_0000;
array[51089] <= 16'b0000_0000_0000_0000;
array[51090] <= 16'b0000_0000_0000_0000;
array[51091] <= 16'b0000_0000_0000_0000;
array[51092] <= 16'b0000_0000_0000_0000;
array[51093] <= 16'b0000_0000_0000_0000;
array[51094] <= 16'b0000_0000_0000_0000;
array[51095] <= 16'b0000_0000_0000_0000;
array[51096] <= 16'b0000_0000_0000_0000;
array[51097] <= 16'b0000_0000_0000_0000;
array[51098] <= 16'b0000_0000_0000_0000;
array[51099] <= 16'b0000_0000_0000_0000;
array[51100] <= 16'b0000_0000_0000_0000;
array[51101] <= 16'b0000_0000_0000_0000;
array[51102] <= 16'b0000_0000_0000_0000;
array[51103] <= 16'b0000_0000_0000_0000;
array[51104] <= 16'b0000_0000_0000_0000;
array[51105] <= 16'b0000_0000_0000_0000;
array[51106] <= 16'b0000_0000_0000_0000;
array[51107] <= 16'b0000_0000_0000_0000;
array[51108] <= 16'b0000_0000_0000_0000;
array[51109] <= 16'b0000_0000_0000_0000;
array[51110] <= 16'b0000_0000_0000_0000;
array[51111] <= 16'b0000_0000_0000_0000;
array[51112] <= 16'b0000_0000_0000_0000;
array[51113] <= 16'b0000_0000_0000_0000;
array[51114] <= 16'b0000_0000_0000_0000;
array[51115] <= 16'b0000_0000_0000_0000;
array[51116] <= 16'b0000_0000_0000_0000;
array[51117] <= 16'b0000_0000_0000_0000;
array[51118] <= 16'b0000_0000_0000_0000;
array[51119] <= 16'b0000_0000_0000_0000;
array[51120] <= 16'b0000_0000_0000_0000;
array[51121] <= 16'b0000_0000_0000_0000;
array[51122] <= 16'b0000_0000_0000_0000;
array[51123] <= 16'b0000_0000_0000_0000;
array[51124] <= 16'b0000_0000_0000_0000;
array[51125] <= 16'b0000_0000_0000_0000;
array[51126] <= 16'b0000_0000_0000_0000;
array[51127] <= 16'b0000_0000_0000_0000;
array[51128] <= 16'b0000_0000_0000_0000;
array[51129] <= 16'b0000_0000_0000_0000;
array[51130] <= 16'b0000_0000_0000_0000;
array[51131] <= 16'b0000_0000_0000_0000;
array[51132] <= 16'b0000_0000_0000_0000;
array[51133] <= 16'b0000_0000_0000_0000;
array[51134] <= 16'b0000_0000_0000_0000;
array[51135] <= 16'b0000_0000_0000_0000;
array[51136] <= 16'b0000_0000_0000_0000;
array[51137] <= 16'b0000_0000_0000_0000;
array[51138] <= 16'b0000_0000_0000_0000;
array[51139] <= 16'b0000_0000_0000_0000;
array[51140] <= 16'b0000_0000_0000_0000;
array[51141] <= 16'b0000_0000_0000_0000;
array[51142] <= 16'b0000_0000_0000_0000;
array[51143] <= 16'b0000_0000_0000_0000;
array[51144] <= 16'b0000_0000_0000_0000;
array[51145] <= 16'b0000_0000_0000_0000;
array[51146] <= 16'b0000_0000_0000_0000;
array[51147] <= 16'b0000_0000_0000_0000;
array[51148] <= 16'b0000_0000_0000_0000;
array[51149] <= 16'b0000_0000_0000_0000;
array[51150] <= 16'b0000_0000_0000_0000;
array[51151] <= 16'b0000_0000_0000_0000;
array[51152] <= 16'b0000_0000_0000_0000;
array[51153] <= 16'b0000_0000_0000_0000;
array[51154] <= 16'b0000_0000_0000_0000;
array[51155] <= 16'b0000_0000_0000_0000;
array[51156] <= 16'b0000_0000_0000_0000;
array[51157] <= 16'b0000_0000_0000_0000;
array[51158] <= 16'b0000_0000_0000_0000;
array[51159] <= 16'b0000_0000_0000_0000;
array[51160] <= 16'b0000_0000_0000_0000;
array[51161] <= 16'b0000_0000_0000_0000;
array[51162] <= 16'b0000_0000_0000_0000;
array[51163] <= 16'b0000_0000_0000_0000;
array[51164] <= 16'b0000_0000_0000_0000;
array[51165] <= 16'b0000_0000_0000_0000;
array[51166] <= 16'b0000_0000_0000_0000;
array[51167] <= 16'b0000_0000_0000_0000;
array[51168] <= 16'b0000_0000_0000_0000;
array[51169] <= 16'b0000_0000_0000_0000;
array[51170] <= 16'b0000_0000_0000_0000;
array[51171] <= 16'b0000_0000_0000_0000;
array[51172] <= 16'b0000_0000_0000_0000;
array[51173] <= 16'b0000_0000_0000_0000;
array[51174] <= 16'b0000_0000_0000_0000;
array[51175] <= 16'b0000_0000_0000_0000;
array[51176] <= 16'b0000_0000_0000_0000;
array[51177] <= 16'b0000_0000_0000_0000;
array[51178] <= 16'b0000_0000_0000_0000;
array[51179] <= 16'b0000_0000_0000_0000;
array[51180] <= 16'b0000_0000_0000_0000;
array[51181] <= 16'b0000_0000_0000_0000;
array[51182] <= 16'b0000_0000_0000_0000;
array[51183] <= 16'b0000_0000_0000_0000;
array[51184] <= 16'b0000_0000_0000_0000;
array[51185] <= 16'b0000_0000_0000_0000;
array[51186] <= 16'b0000_0000_0000_0000;
array[51187] <= 16'b0000_0000_0000_0000;
array[51188] <= 16'b0000_0000_0000_0000;
array[51189] <= 16'b0000_0000_0000_0000;
array[51190] <= 16'b0000_0000_0000_0000;
array[51191] <= 16'b0000_0000_0000_0000;
array[51192] <= 16'b0000_0000_0000_0000;
array[51193] <= 16'b0000_0000_0000_0000;
array[51194] <= 16'b0000_0000_0000_0000;
array[51195] <= 16'b0000_0000_0000_0000;
array[51196] <= 16'b0000_0000_0000_0000;
array[51197] <= 16'b0000_0000_0000_0000;
array[51198] <= 16'b0000_0000_0000_0000;
array[51199] <= 16'b0000_0000_0000_0000;
array[51200] <= 16'b0000_0000_0000_0000;
array[51201] <= 16'b0000_0000_0000_0000;
array[51202] <= 16'b0000_0000_0000_0000;
array[51203] <= 16'b0000_0000_0000_0000;
array[51204] <= 16'b0000_0000_0000_0000;
array[51205] <= 16'b0000_0000_0000_0000;
array[51206] <= 16'b0000_0000_0000_0000;
array[51207] <= 16'b0000_0000_0000_0000;
array[51208] <= 16'b0000_0000_0000_0000;
array[51209] <= 16'b0000_0000_0000_0000;
array[51210] <= 16'b0000_0000_0000_0000;
array[51211] <= 16'b0000_0000_0000_0000;
array[51212] <= 16'b0000_0000_0000_0000;
array[51213] <= 16'b0000_0000_0000_0000;
array[51214] <= 16'b0000_0000_0000_0000;
array[51215] <= 16'b0000_0000_0000_0000;
array[51216] <= 16'b0000_0000_0000_0000;
array[51217] <= 16'b0000_0000_0000_0000;
array[51218] <= 16'b0000_0000_0000_0000;
array[51219] <= 16'b0000_0000_0000_0000;
array[51220] <= 16'b0000_0000_0000_0000;
array[51221] <= 16'b0000_0000_0000_0000;
array[51222] <= 16'b0000_0000_0000_0000;
array[51223] <= 16'b0000_0000_0000_0000;
array[51224] <= 16'b0000_0000_0000_0000;
array[51225] <= 16'b0000_0000_0000_0000;
array[51226] <= 16'b0000_0000_0000_0000;
array[51227] <= 16'b0000_0000_0000_0000;
array[51228] <= 16'b0000_0000_0000_0000;
array[51229] <= 16'b0000_0000_0000_0000;
array[51230] <= 16'b0000_0000_0000_0000;
array[51231] <= 16'b0000_0000_0000_0000;
array[51232] <= 16'b0000_0000_0000_0000;
array[51233] <= 16'b0000_0000_0000_0000;
array[51234] <= 16'b0000_0000_0000_0000;
array[51235] <= 16'b0000_0000_0000_0000;
array[51236] <= 16'b0000_0000_0000_0000;
array[51237] <= 16'b0000_0000_0000_0000;
array[51238] <= 16'b0000_0000_0000_0000;
array[51239] <= 16'b0000_0000_0000_0000;
array[51240] <= 16'b0000_0000_0000_0000;
array[51241] <= 16'b0000_0000_0000_0000;
array[51242] <= 16'b0000_0000_0000_0000;
array[51243] <= 16'b0000_0000_0000_0000;
array[51244] <= 16'b0000_0000_0000_0000;
array[51245] <= 16'b0000_0000_0000_0000;
array[51246] <= 16'b0000_0000_0000_0000;
array[51247] <= 16'b0000_0000_0000_0000;
array[51248] <= 16'b0000_0000_0000_0000;
array[51249] <= 16'b0000_0000_0000_0000;
array[51250] <= 16'b0000_0000_0000_0000;
array[51251] <= 16'b0000_0000_0000_0000;
array[51252] <= 16'b0000_0000_0000_0000;
array[51253] <= 16'b0000_0000_0000_0000;
array[51254] <= 16'b0000_0000_0000_0000;
array[51255] <= 16'b0000_0000_0000_0000;
array[51256] <= 16'b0000_0000_0000_0000;
array[51257] <= 16'b0000_0000_0000_0000;
array[51258] <= 16'b0000_0000_0000_0000;
array[51259] <= 16'b0000_0000_0000_0000;
array[51260] <= 16'b0000_0000_0000_0000;
array[51261] <= 16'b0000_0000_0000_0000;
array[51262] <= 16'b0000_0000_0000_0000;
array[51263] <= 16'b0000_0000_0000_0000;
array[51264] <= 16'b0000_0000_0000_0000;
array[51265] <= 16'b0000_0000_0000_0000;
array[51266] <= 16'b0000_0000_0000_0000;
array[51267] <= 16'b0000_0000_0000_0000;
array[51268] <= 16'b0000_0000_0000_0000;
array[51269] <= 16'b0000_0000_0000_0000;
array[51270] <= 16'b0000_0000_0000_0000;
array[51271] <= 16'b0000_0000_0000_0000;
array[51272] <= 16'b0000_0000_0000_0000;
array[51273] <= 16'b0000_0000_0000_0000;
array[51274] <= 16'b0000_0000_0000_0000;
array[51275] <= 16'b0000_0000_0000_0000;
array[51276] <= 16'b0000_0000_0000_0000;
array[51277] <= 16'b0000_0000_0000_0000;
array[51278] <= 16'b0000_0000_0000_0000;
array[51279] <= 16'b0000_0000_0000_0000;
array[51280] <= 16'b0000_0000_0000_0000;
array[51281] <= 16'b0000_0000_0000_0000;
array[51282] <= 16'b0000_0000_0000_0000;
array[51283] <= 16'b0000_0000_0000_0000;
array[51284] <= 16'b0000_0000_0000_0000;
array[51285] <= 16'b0000_0000_0000_0000;
array[51286] <= 16'b0000_0000_0000_0000;
array[51287] <= 16'b0000_0000_0000_0000;
array[51288] <= 16'b0000_0000_0000_0000;
array[51289] <= 16'b0000_0000_0000_0000;
array[51290] <= 16'b0000_0000_0000_0000;
array[51291] <= 16'b0000_0000_0000_0000;
array[51292] <= 16'b0000_0000_0000_0000;
array[51293] <= 16'b0000_0000_0000_0000;
array[51294] <= 16'b0000_0000_0000_0000;
array[51295] <= 16'b0000_0000_0000_0000;
array[51296] <= 16'b0000_0000_0000_0000;
array[51297] <= 16'b0000_0000_0000_0000;
array[51298] <= 16'b0000_0000_0000_0000;
array[51299] <= 16'b0000_0000_0000_0000;
array[51300] <= 16'b0000_0000_0000_0000;
array[51301] <= 16'b0000_0000_0000_0000;
array[51302] <= 16'b0000_0000_0000_0000;
array[51303] <= 16'b0000_0000_0000_0000;
array[51304] <= 16'b0000_0000_0000_0000;
array[51305] <= 16'b0000_0000_0000_0000;
array[51306] <= 16'b0000_0000_0000_0000;
array[51307] <= 16'b0000_0000_0000_0000;
array[51308] <= 16'b0000_0000_0000_0000;
array[51309] <= 16'b0000_0000_0000_0000;
array[51310] <= 16'b0000_0000_0000_0000;
array[51311] <= 16'b0000_0000_0000_0000;
array[51312] <= 16'b0000_0000_0000_0000;
array[51313] <= 16'b0000_0000_0000_0000;
array[51314] <= 16'b0000_0000_0000_0000;
array[51315] <= 16'b0000_0000_0000_0000;
array[51316] <= 16'b0000_0000_0000_0000;
array[51317] <= 16'b0000_0000_0000_0000;
array[51318] <= 16'b0000_0000_0000_0000;
array[51319] <= 16'b0000_0000_0000_0000;
array[51320] <= 16'b0000_0000_0000_0000;
array[51321] <= 16'b0000_0000_0000_0000;
array[51322] <= 16'b0000_0000_0000_0000;
array[51323] <= 16'b0000_0000_0000_0000;
array[51324] <= 16'b0000_0000_0000_0000;
array[51325] <= 16'b0000_0000_0000_0000;
array[51326] <= 16'b0000_0000_0000_0000;
array[51327] <= 16'b0000_0000_0000_0000;
array[51328] <= 16'b0000_0000_0000_0000;
array[51329] <= 16'b0000_0000_0000_0000;
array[51330] <= 16'b0000_0000_0000_0000;
array[51331] <= 16'b0000_0000_0000_0000;
array[51332] <= 16'b0000_0000_0000_0000;
array[51333] <= 16'b0000_0000_0000_0000;
array[51334] <= 16'b0000_0000_0000_0000;
array[51335] <= 16'b0000_0000_0000_0000;
array[51336] <= 16'b0000_0000_0000_0000;
array[51337] <= 16'b0000_0000_0000_0000;
array[51338] <= 16'b0000_0000_0000_0000;
array[51339] <= 16'b0000_0000_0000_0000;
array[51340] <= 16'b0000_0000_0000_0000;
array[51341] <= 16'b0000_0000_0000_0000;
array[51342] <= 16'b0000_0000_0000_0000;
array[51343] <= 16'b0000_0000_0000_0000;
array[51344] <= 16'b0000_0000_0000_0000;
array[51345] <= 16'b0000_0000_0000_0000;
array[51346] <= 16'b0000_0000_0000_0000;
array[51347] <= 16'b0000_0000_0000_0000;
array[51348] <= 16'b0000_0000_0000_0000;
array[51349] <= 16'b0000_0000_0000_0000;
array[51350] <= 16'b0000_0000_0000_0000;
array[51351] <= 16'b0000_0000_0000_0000;
array[51352] <= 16'b0000_0000_0000_0000;
array[51353] <= 16'b0000_0000_0000_0000;
array[51354] <= 16'b0000_0000_0000_0000;
array[51355] <= 16'b0000_0000_0000_0000;
array[51356] <= 16'b0000_0000_0000_0000;
array[51357] <= 16'b0000_0000_0000_0000;
array[51358] <= 16'b0000_0000_0000_0000;
array[51359] <= 16'b0000_0000_0000_0000;
array[51360] <= 16'b0000_0000_0000_0000;
array[51361] <= 16'b0000_0000_0000_0000;
array[51362] <= 16'b0000_0000_0000_0000;
array[51363] <= 16'b0000_0000_0000_0000;
array[51364] <= 16'b0000_0000_0000_0000;
array[51365] <= 16'b0000_0000_0000_0000;
array[51366] <= 16'b0000_0000_0000_0000;
array[51367] <= 16'b0000_0000_0000_0000;
array[51368] <= 16'b0000_0000_0000_0000;
array[51369] <= 16'b0000_0000_0000_0000;
array[51370] <= 16'b0000_0000_0000_0000;
array[51371] <= 16'b0000_0000_0000_0000;
array[51372] <= 16'b0000_0000_0000_0000;
array[51373] <= 16'b0000_0000_0000_0000;
array[51374] <= 16'b0000_0000_0000_0000;
array[51375] <= 16'b0000_0000_0000_0000;
array[51376] <= 16'b0000_0000_0000_0000;
array[51377] <= 16'b0000_0000_0000_0000;
array[51378] <= 16'b0000_0000_0000_0000;
array[51379] <= 16'b0000_0000_0000_0000;
array[51380] <= 16'b0000_0000_0000_0000;
array[51381] <= 16'b0000_0000_0000_0000;
array[51382] <= 16'b0000_0000_0000_0000;
array[51383] <= 16'b0000_0000_0000_0000;
array[51384] <= 16'b0000_0000_0000_0000;
array[51385] <= 16'b0000_0000_0000_0000;
array[51386] <= 16'b0000_0000_0000_0000;
array[51387] <= 16'b0000_0000_0000_0000;
array[51388] <= 16'b0000_0000_0000_0000;
array[51389] <= 16'b0000_0000_0000_0000;
array[51390] <= 16'b0000_0000_0000_0000;
array[51391] <= 16'b0000_0000_0000_0000;
array[51392] <= 16'b0000_0000_0000_0000;
array[51393] <= 16'b0000_0000_0000_0000;
array[51394] <= 16'b0000_0000_0000_0000;
array[51395] <= 16'b0000_0000_0000_0000;
array[51396] <= 16'b0000_0000_0000_0000;
array[51397] <= 16'b0000_0000_0000_0000;
array[51398] <= 16'b0000_0000_0000_0000;
array[51399] <= 16'b0000_0000_0000_0000;
array[51400] <= 16'b0000_0000_0000_0000;
array[51401] <= 16'b0000_0000_0000_0000;
array[51402] <= 16'b0000_0000_0000_0000;
array[51403] <= 16'b0000_0000_0000_0000;
array[51404] <= 16'b0000_0000_0000_0000;
array[51405] <= 16'b0000_0000_0000_0000;
array[51406] <= 16'b0000_0000_0000_0000;
array[51407] <= 16'b0000_0000_0000_0000;
array[51408] <= 16'b0000_0000_0000_0000;
array[51409] <= 16'b0000_0000_0000_0000;
array[51410] <= 16'b0000_0000_0000_0000;
array[51411] <= 16'b0000_0000_0000_0000;
array[51412] <= 16'b0000_0000_0000_0000;
array[51413] <= 16'b0000_0000_0000_0000;
array[51414] <= 16'b0000_0000_0000_0000;
array[51415] <= 16'b0000_0000_0000_0000;
array[51416] <= 16'b0000_0000_0000_0000;
array[51417] <= 16'b0000_0000_0000_0000;
array[51418] <= 16'b0000_0000_0000_0000;
array[51419] <= 16'b0000_0000_0000_0000;
array[51420] <= 16'b0000_0000_0000_0000;
array[51421] <= 16'b0000_0000_0000_0000;
array[51422] <= 16'b0000_0000_0000_0000;
array[51423] <= 16'b0000_0000_0000_0000;
array[51424] <= 16'b0000_0000_0000_0000;
array[51425] <= 16'b0000_0000_0000_0000;
array[51426] <= 16'b0000_0000_0000_0000;
array[51427] <= 16'b0000_0000_0000_0000;
array[51428] <= 16'b0000_0000_0000_0000;
array[51429] <= 16'b0000_0000_0000_0000;
array[51430] <= 16'b0000_0000_0000_0000;
array[51431] <= 16'b0000_0000_0000_0000;
array[51432] <= 16'b0000_0000_0000_0000;
array[51433] <= 16'b0000_0000_0000_0000;
array[51434] <= 16'b0000_0000_0000_0000;
array[51435] <= 16'b0000_0000_0000_0000;
array[51436] <= 16'b0000_0000_0000_0000;
array[51437] <= 16'b0000_0000_0000_0000;
array[51438] <= 16'b0000_0000_0000_0000;
array[51439] <= 16'b0000_0000_0000_0000;
array[51440] <= 16'b0000_0000_0000_0000;
array[51441] <= 16'b0000_0000_0000_0000;
array[51442] <= 16'b0000_0000_0000_0000;
array[51443] <= 16'b0000_0000_0000_0000;
array[51444] <= 16'b0000_0000_0000_0000;
array[51445] <= 16'b0000_0000_0000_0000;
array[51446] <= 16'b0000_0000_0000_0000;
array[51447] <= 16'b0000_0000_0000_0000;
array[51448] <= 16'b0000_0000_0000_0000;
array[51449] <= 16'b0000_0000_0000_0000;
array[51450] <= 16'b0000_0000_0000_0000;
array[51451] <= 16'b0000_0000_0000_0000;
array[51452] <= 16'b0000_0000_0000_0000;
array[51453] <= 16'b0000_0000_0000_0000;
array[51454] <= 16'b0000_0000_0000_0000;
array[51455] <= 16'b0000_0000_0000_0000;
array[51456] <= 16'b0000_0000_0000_0000;
array[51457] <= 16'b0000_0000_0000_0000;
array[51458] <= 16'b0000_0000_0000_0000;
array[51459] <= 16'b0000_0000_0000_0000;
array[51460] <= 16'b0000_0000_0000_0000;
array[51461] <= 16'b0000_0000_0000_0000;
array[51462] <= 16'b0000_0000_0000_0000;
array[51463] <= 16'b0000_0000_0000_0000;
array[51464] <= 16'b0000_0000_0000_0000;
array[51465] <= 16'b0000_0000_0000_0000;
array[51466] <= 16'b0000_0000_0000_0000;
array[51467] <= 16'b0000_0000_0000_0000;
array[51468] <= 16'b0000_0000_0000_0000;
array[51469] <= 16'b0000_0000_0000_0000;
array[51470] <= 16'b0000_0000_0000_0000;
array[51471] <= 16'b0000_0000_0000_0000;
array[51472] <= 16'b0000_0000_0000_0000;
array[51473] <= 16'b0000_0000_0000_0000;
array[51474] <= 16'b0000_0000_0000_0000;
array[51475] <= 16'b0000_0000_0000_0000;
array[51476] <= 16'b0000_0000_0000_0000;
array[51477] <= 16'b0000_0000_0000_0000;
array[51478] <= 16'b0000_0000_0000_0000;
array[51479] <= 16'b0000_0000_0000_0000;
array[51480] <= 16'b0000_0000_0000_0000;
array[51481] <= 16'b0000_0000_0000_0000;
array[51482] <= 16'b0000_0000_0000_0000;
array[51483] <= 16'b0000_0000_0000_0000;
array[51484] <= 16'b0000_0000_0000_0000;
array[51485] <= 16'b0000_0000_0000_0000;
array[51486] <= 16'b0000_0000_0000_0000;
array[51487] <= 16'b0000_0000_0000_0000;
array[51488] <= 16'b0000_0000_0000_0000;
array[51489] <= 16'b0000_0000_0000_0000;
array[51490] <= 16'b0000_0000_0000_0000;
array[51491] <= 16'b0000_0000_0000_0000;
array[51492] <= 16'b0000_0000_0000_0000;
array[51493] <= 16'b0000_0000_0000_0000;
array[51494] <= 16'b0000_0000_0000_0000;
array[51495] <= 16'b0000_0000_0000_0000;
array[51496] <= 16'b0000_0000_0000_0000;
array[51497] <= 16'b0000_0000_0000_0000;
array[51498] <= 16'b0000_0000_0000_0000;
array[51499] <= 16'b0000_0000_0000_0000;
array[51500] <= 16'b0000_0000_0000_0000;
array[51501] <= 16'b0000_0000_0000_0000;
array[51502] <= 16'b0000_0000_0000_0000;
array[51503] <= 16'b0000_0000_0000_0000;
array[51504] <= 16'b0000_0000_0000_0000;
array[51505] <= 16'b0000_0000_0000_0000;
array[51506] <= 16'b0000_0000_0000_0000;
array[51507] <= 16'b0000_0000_0000_0000;
array[51508] <= 16'b0000_0000_0000_0000;
array[51509] <= 16'b0000_0000_0000_0000;
array[51510] <= 16'b0000_0000_0000_0000;
array[51511] <= 16'b0000_0000_0000_0000;
array[51512] <= 16'b0000_0000_0000_0000;
array[51513] <= 16'b0000_0000_0000_0000;
array[51514] <= 16'b0000_0000_0000_0000;
array[51515] <= 16'b0000_0000_0000_0000;
array[51516] <= 16'b0000_0000_0000_0000;
array[51517] <= 16'b0000_0000_0000_0000;
array[51518] <= 16'b0000_0000_0000_0000;
array[51519] <= 16'b0000_0000_0000_0000;
array[51520] <= 16'b0000_0000_0000_0000;
array[51521] <= 16'b0000_0000_0000_0000;
array[51522] <= 16'b0000_0000_0000_0000;
array[51523] <= 16'b0000_0000_0000_0000;
array[51524] <= 16'b0000_0000_0000_0000;
array[51525] <= 16'b0000_0000_0000_0000;
array[51526] <= 16'b0000_0000_0000_0000;
array[51527] <= 16'b0000_0000_0000_0000;
array[51528] <= 16'b0000_0000_0000_0000;
array[51529] <= 16'b0000_0000_0000_0000;
array[51530] <= 16'b0000_0000_0000_0000;
array[51531] <= 16'b0000_0000_0000_0000;
array[51532] <= 16'b0000_0000_0000_0000;
array[51533] <= 16'b0000_0000_0000_0000;
array[51534] <= 16'b0000_0000_0000_0000;
array[51535] <= 16'b0000_0000_0000_0000;
array[51536] <= 16'b0000_0000_0000_0000;
array[51537] <= 16'b0000_0000_0000_0000;
array[51538] <= 16'b0000_0000_0000_0000;
array[51539] <= 16'b0000_0000_0000_0000;
array[51540] <= 16'b0000_0000_0000_0000;
array[51541] <= 16'b0000_0000_0000_0000;
array[51542] <= 16'b0000_0000_0000_0000;
array[51543] <= 16'b0000_0000_0000_0000;
array[51544] <= 16'b0000_0000_0000_0000;
array[51545] <= 16'b0000_0000_0000_0000;
array[51546] <= 16'b0000_0000_0000_0000;
array[51547] <= 16'b0000_0000_0000_0000;
array[51548] <= 16'b0000_0000_0000_0000;
array[51549] <= 16'b0000_0000_0000_0000;
array[51550] <= 16'b0000_0000_0000_0000;
array[51551] <= 16'b0000_0000_0000_0000;
array[51552] <= 16'b0000_0000_0000_0000;
array[51553] <= 16'b0000_0000_0000_0000;
array[51554] <= 16'b0000_0000_0000_0000;
array[51555] <= 16'b0000_0000_0000_0000;
array[51556] <= 16'b0000_0000_0000_0000;
array[51557] <= 16'b0000_0000_0000_0000;
array[51558] <= 16'b0000_0000_0000_0000;
array[51559] <= 16'b0000_0000_0000_0000;
array[51560] <= 16'b0000_0000_0000_0000;
array[51561] <= 16'b0000_0000_0000_0000;
array[51562] <= 16'b0000_0000_0000_0000;
array[51563] <= 16'b0000_0000_0000_0000;
array[51564] <= 16'b0000_0000_0000_0000;
array[51565] <= 16'b0000_0000_0000_0000;
array[51566] <= 16'b0000_0000_0000_0000;
array[51567] <= 16'b0000_0000_0000_0000;
array[51568] <= 16'b0000_0000_0000_0000;
array[51569] <= 16'b0000_0000_0000_0000;
array[51570] <= 16'b0000_0000_0000_0000;
array[51571] <= 16'b0000_0000_0000_0000;
array[51572] <= 16'b0000_0000_0000_0000;
array[51573] <= 16'b0000_0000_0000_0000;
array[51574] <= 16'b0000_0000_0000_0000;
array[51575] <= 16'b0000_0000_0000_0000;
array[51576] <= 16'b0000_0000_0000_0000;
array[51577] <= 16'b0000_0000_0000_0000;
array[51578] <= 16'b0000_0000_0000_0000;
array[51579] <= 16'b0000_0000_0000_0000;
array[51580] <= 16'b0000_0000_0000_0000;
array[51581] <= 16'b0000_0000_0000_0000;
array[51582] <= 16'b0000_0000_0000_0000;
array[51583] <= 16'b0000_0000_0000_0000;
array[51584] <= 16'b0000_0000_0000_0000;
array[51585] <= 16'b0000_0000_0000_0000;
array[51586] <= 16'b0000_0000_0000_0000;
array[51587] <= 16'b0000_0000_0000_0000;
array[51588] <= 16'b0000_0000_0000_0000;
array[51589] <= 16'b0000_0000_0000_0000;
array[51590] <= 16'b0000_0000_0000_0000;
array[51591] <= 16'b0000_0000_0000_0000;
array[51592] <= 16'b0000_0000_0000_0000;
array[51593] <= 16'b0000_0000_0000_0000;
array[51594] <= 16'b0000_0000_0000_0000;
array[51595] <= 16'b0000_0000_0000_0000;
array[51596] <= 16'b0000_0000_0000_0000;
array[51597] <= 16'b0000_0000_0000_0000;
array[51598] <= 16'b0000_0000_0000_0000;
array[51599] <= 16'b0000_0000_0000_0000;
array[51600] <= 16'b0000_0000_0000_0000;
array[51601] <= 16'b0000_0000_0000_0000;
array[51602] <= 16'b0000_0000_0000_0000;
array[51603] <= 16'b0000_0000_0000_0000;
array[51604] <= 16'b0000_0000_0000_0000;
array[51605] <= 16'b0000_0000_0000_0000;
array[51606] <= 16'b0000_0000_0000_0000;
array[51607] <= 16'b0000_0000_0000_0000;
array[51608] <= 16'b0000_0000_0000_0000;
array[51609] <= 16'b0000_0000_0000_0000;
array[51610] <= 16'b0000_0000_0000_0000;
array[51611] <= 16'b0000_0000_0000_0000;
array[51612] <= 16'b0000_0000_0000_0000;
array[51613] <= 16'b0000_0000_0000_0000;
array[51614] <= 16'b0000_0000_0000_0000;
array[51615] <= 16'b0000_0000_0000_0000;
array[51616] <= 16'b0000_0000_0000_0000;
array[51617] <= 16'b0000_0000_0000_0000;
array[51618] <= 16'b0000_0000_0000_0000;
array[51619] <= 16'b0000_0000_0000_0000;
array[51620] <= 16'b0000_0000_0000_0000;
array[51621] <= 16'b0000_0000_0000_0000;
array[51622] <= 16'b0000_0000_0000_0000;
array[51623] <= 16'b0000_0000_0000_0000;
array[51624] <= 16'b0000_0000_0000_0000;
array[51625] <= 16'b0000_0000_0000_0000;
array[51626] <= 16'b0000_0000_0000_0000;
array[51627] <= 16'b0000_0000_0000_0000;
array[51628] <= 16'b0000_0000_0000_0000;
array[51629] <= 16'b0000_0000_0000_0000;
array[51630] <= 16'b0000_0000_0000_0000;
array[51631] <= 16'b0000_0000_0000_0000;
array[51632] <= 16'b0000_0000_0000_0000;
array[51633] <= 16'b0000_0000_0000_0000;
array[51634] <= 16'b0000_0000_0000_0000;
array[51635] <= 16'b0000_0000_0000_0000;
array[51636] <= 16'b0000_0000_0000_0000;
array[51637] <= 16'b0000_0000_0000_0000;
array[51638] <= 16'b0000_0000_0000_0000;
array[51639] <= 16'b0000_0000_0000_0000;
array[51640] <= 16'b0000_0000_0000_0000;
array[51641] <= 16'b0000_0000_0000_0000;
array[51642] <= 16'b0000_0000_0000_0000;
array[51643] <= 16'b0000_0000_0000_0000;
array[51644] <= 16'b0000_0000_0000_0000;
array[51645] <= 16'b0000_0000_0000_0000;
array[51646] <= 16'b0000_0000_0000_0000;
array[51647] <= 16'b0000_0000_0000_0000;
array[51648] <= 16'b0000_0000_0000_0000;
array[51649] <= 16'b0000_0000_0000_0000;
array[51650] <= 16'b0000_0000_0000_0000;
array[51651] <= 16'b0000_0000_0000_0000;
array[51652] <= 16'b0000_0000_0000_0000;
array[51653] <= 16'b0000_0000_0000_0000;
array[51654] <= 16'b0000_0000_0000_0000;
array[51655] <= 16'b0000_0000_0000_0000;
array[51656] <= 16'b0000_0000_0000_0000;
array[51657] <= 16'b0000_0000_0000_0000;
array[51658] <= 16'b0000_0000_0000_0000;
array[51659] <= 16'b0000_0000_0000_0000;
array[51660] <= 16'b0000_0000_0000_0000;
array[51661] <= 16'b0000_0000_0000_0000;
array[51662] <= 16'b0000_0000_0000_0000;
array[51663] <= 16'b0000_0000_0000_0000;
array[51664] <= 16'b0000_0000_0000_0000;
array[51665] <= 16'b0000_0000_0000_0000;
array[51666] <= 16'b0000_0000_0000_0000;
array[51667] <= 16'b0000_0000_0000_0000;
array[51668] <= 16'b0000_0000_0000_0000;
array[51669] <= 16'b0000_0000_0000_0000;
array[51670] <= 16'b0000_0000_0000_0000;
array[51671] <= 16'b0000_0000_0000_0000;
array[51672] <= 16'b0000_0000_0000_0000;
array[51673] <= 16'b0000_0000_0000_0000;
array[51674] <= 16'b0000_0000_0000_0000;
array[51675] <= 16'b0000_0000_0000_0000;
array[51676] <= 16'b0000_0000_0000_0000;
array[51677] <= 16'b0000_0000_0000_0000;
array[51678] <= 16'b0000_0000_0000_0000;
array[51679] <= 16'b0000_0000_0000_0000;
array[51680] <= 16'b0000_0000_0000_0000;
array[51681] <= 16'b0000_0000_0000_0000;
array[51682] <= 16'b0000_0000_0000_0000;
array[51683] <= 16'b0000_0000_0000_0000;
array[51684] <= 16'b0000_0000_0000_0000;
array[51685] <= 16'b0000_0000_0000_0000;
array[51686] <= 16'b0000_0000_0000_0000;
array[51687] <= 16'b0000_0000_0000_0000;
array[51688] <= 16'b0000_0000_0000_0000;
array[51689] <= 16'b0000_0000_0000_0000;
array[51690] <= 16'b0000_0000_0000_0000;
array[51691] <= 16'b0000_0000_0000_0000;
array[51692] <= 16'b0000_0000_0000_0000;
array[51693] <= 16'b0000_0000_0000_0000;
array[51694] <= 16'b0000_0000_0000_0000;
array[51695] <= 16'b0000_0000_0000_0000;
array[51696] <= 16'b0000_0000_0000_0000;
array[51697] <= 16'b0000_0000_0000_0000;
array[51698] <= 16'b0000_0000_0000_0000;
array[51699] <= 16'b0000_0000_0000_0000;
array[51700] <= 16'b0000_0000_0000_0000;
array[51701] <= 16'b0000_0000_0000_0000;
array[51702] <= 16'b0000_0000_0000_0000;
array[51703] <= 16'b0000_0000_0000_0000;
array[51704] <= 16'b0000_0000_0000_0000;
array[51705] <= 16'b0000_0000_0000_0000;
array[51706] <= 16'b0000_0000_0000_0000;
array[51707] <= 16'b0000_0000_0000_0000;
array[51708] <= 16'b0000_0000_0000_0000;
array[51709] <= 16'b0000_0000_0000_0000;
array[51710] <= 16'b0000_0000_0000_0000;
array[51711] <= 16'b0000_0000_0000_0000;
array[51712] <= 16'b0000_0000_0000_0000;
array[51713] <= 16'b0000_0000_0000_0000;
array[51714] <= 16'b0000_0000_0000_0000;
array[51715] <= 16'b0000_0000_0000_0000;
array[51716] <= 16'b0000_0000_0000_0000;
array[51717] <= 16'b0000_0000_0000_0000;
array[51718] <= 16'b0000_0000_0000_0000;
array[51719] <= 16'b0000_0000_0000_0000;
array[51720] <= 16'b0000_0000_0000_0000;
array[51721] <= 16'b0000_0000_0000_0000;
array[51722] <= 16'b0000_0000_0000_0000;
array[51723] <= 16'b0000_0000_0000_0000;
array[51724] <= 16'b0000_0000_0000_0000;
array[51725] <= 16'b0000_0000_0000_0000;
array[51726] <= 16'b0000_0000_0000_0000;
array[51727] <= 16'b0000_0000_0000_0000;
array[51728] <= 16'b0000_0000_0000_0000;
array[51729] <= 16'b0000_0000_0000_0000;
array[51730] <= 16'b0000_0000_0000_0000;
array[51731] <= 16'b0000_0000_0000_0000;
array[51732] <= 16'b0000_0000_0000_0000;
array[51733] <= 16'b0000_0000_0000_0000;
array[51734] <= 16'b0000_0000_0000_0000;
array[51735] <= 16'b0000_0000_0000_0000;
array[51736] <= 16'b0000_0000_0000_0000;
array[51737] <= 16'b0000_0000_0000_0000;
array[51738] <= 16'b0000_0000_0000_0000;
array[51739] <= 16'b0000_0000_0000_0000;
array[51740] <= 16'b0000_0000_0000_0000;
array[51741] <= 16'b0000_0000_0000_0000;
array[51742] <= 16'b0000_0000_0000_0000;
array[51743] <= 16'b0000_0000_0000_0000;
array[51744] <= 16'b0000_0000_0000_0000;
array[51745] <= 16'b0000_0000_0000_0000;
array[51746] <= 16'b0000_0000_0000_0000;
array[51747] <= 16'b0000_0000_0000_0000;
array[51748] <= 16'b0000_0000_0000_0000;
array[51749] <= 16'b0000_0000_0000_0000;
array[51750] <= 16'b0000_0000_0000_0000;
array[51751] <= 16'b0000_0000_0000_0000;
array[51752] <= 16'b0000_0000_0000_0000;
array[51753] <= 16'b0000_0000_0000_0000;
array[51754] <= 16'b0000_0000_0000_0000;
array[51755] <= 16'b0000_0000_0000_0000;
array[51756] <= 16'b0000_0000_0000_0000;
array[51757] <= 16'b0000_0000_0000_0000;
array[51758] <= 16'b0000_0000_0000_0000;
array[51759] <= 16'b0000_0000_0000_0000;
array[51760] <= 16'b0000_0000_0000_0000;
array[51761] <= 16'b0000_0000_0000_0000;
array[51762] <= 16'b0000_0000_0000_0000;
array[51763] <= 16'b0000_0000_0000_0000;
array[51764] <= 16'b0000_0000_0000_0000;
array[51765] <= 16'b0000_0000_0000_0000;
array[51766] <= 16'b0000_0000_0000_0000;
array[51767] <= 16'b0000_0000_0000_0000;
array[51768] <= 16'b0000_0000_0000_0000;
array[51769] <= 16'b0000_0000_0000_0000;
array[51770] <= 16'b0000_0000_0000_0000;
array[51771] <= 16'b0000_0000_0000_0000;
array[51772] <= 16'b0000_0000_0000_0000;
array[51773] <= 16'b0000_0000_0000_0000;
array[51774] <= 16'b0000_0000_0000_0000;
array[51775] <= 16'b0000_0000_0000_0000;
array[51776] <= 16'b0000_0000_0000_0000;
array[51777] <= 16'b0000_0000_0000_0000;
array[51778] <= 16'b0000_0000_0000_0000;
array[51779] <= 16'b0000_0000_0000_0000;
array[51780] <= 16'b0000_0000_0000_0000;
array[51781] <= 16'b0000_0000_0000_0000;
array[51782] <= 16'b0000_0000_0000_0000;
array[51783] <= 16'b0000_0000_0000_0000;
array[51784] <= 16'b0000_0000_0000_0000;
array[51785] <= 16'b0000_0000_0000_0000;
array[51786] <= 16'b0000_0000_0000_0000;
array[51787] <= 16'b0000_0000_0000_0000;
array[51788] <= 16'b0000_0000_0000_0000;
array[51789] <= 16'b0000_0000_0000_0000;
array[51790] <= 16'b0000_0000_0000_0000;
array[51791] <= 16'b0000_0000_0000_0000;
array[51792] <= 16'b0000_0000_0000_0000;
array[51793] <= 16'b0000_0000_0000_0000;
array[51794] <= 16'b0000_0000_0000_0000;
array[51795] <= 16'b0000_0000_0000_0000;
array[51796] <= 16'b0000_0000_0000_0000;
array[51797] <= 16'b0000_0000_0000_0000;
array[51798] <= 16'b0000_0000_0000_0000;
array[51799] <= 16'b0000_0000_0000_0000;
array[51800] <= 16'b0000_0000_0000_0000;
array[51801] <= 16'b0000_0000_0000_0000;
array[51802] <= 16'b0000_0000_0000_0000;
array[51803] <= 16'b0000_0000_0000_0000;
array[51804] <= 16'b0000_0000_0000_0000;
array[51805] <= 16'b0000_0000_0000_0000;
array[51806] <= 16'b0000_0000_0000_0000;
array[51807] <= 16'b0000_0000_0000_0000;
array[51808] <= 16'b0000_0000_0000_0000;
array[51809] <= 16'b0000_0000_0000_0000;
array[51810] <= 16'b0000_0000_0000_0000;
array[51811] <= 16'b0000_0000_0000_0000;
array[51812] <= 16'b0000_0000_0000_0000;
array[51813] <= 16'b0000_0000_0000_0000;
array[51814] <= 16'b0000_0000_0000_0000;
array[51815] <= 16'b0000_0000_0000_0000;
array[51816] <= 16'b0000_0000_0000_0000;
array[51817] <= 16'b0000_0000_0000_0000;
array[51818] <= 16'b0000_0000_0000_0000;
array[51819] <= 16'b0000_0000_0000_0000;
array[51820] <= 16'b0000_0000_0000_0000;
array[51821] <= 16'b0000_0000_0000_0000;
array[51822] <= 16'b0000_0000_0000_0000;
array[51823] <= 16'b0000_0000_0000_0000;
array[51824] <= 16'b0000_0000_0000_0000;
array[51825] <= 16'b0000_0000_0000_0000;
array[51826] <= 16'b0000_0000_0000_0000;
array[51827] <= 16'b0000_0000_0000_0000;
array[51828] <= 16'b0000_0000_0000_0000;
array[51829] <= 16'b0000_0000_0000_0000;
array[51830] <= 16'b0000_0000_0000_0000;
array[51831] <= 16'b0000_0000_0000_0000;
array[51832] <= 16'b0000_0000_0000_0000;
array[51833] <= 16'b0000_0000_0000_0000;
array[51834] <= 16'b0000_0000_0000_0000;
array[51835] <= 16'b0000_0000_0000_0000;
array[51836] <= 16'b0000_0000_0000_0000;
array[51837] <= 16'b0000_0000_0000_0000;
array[51838] <= 16'b0000_0000_0000_0000;
array[51839] <= 16'b0000_0000_0000_0000;
array[51840] <= 16'b0000_0000_0000_0000;
array[51841] <= 16'b0000_0000_0000_0000;
array[51842] <= 16'b0000_0000_0000_0000;
array[51843] <= 16'b0000_0000_0000_0000;
array[51844] <= 16'b0000_0000_0000_0000;
array[51845] <= 16'b0000_0000_0000_0000;
array[51846] <= 16'b0000_0000_0000_0000;
array[51847] <= 16'b0000_0000_0000_0000;
array[51848] <= 16'b0000_0000_0000_0000;
array[51849] <= 16'b0000_0000_0000_0000;
array[51850] <= 16'b0000_0000_0000_0000;
array[51851] <= 16'b0000_0000_0000_0000;
array[51852] <= 16'b0000_0000_0000_0000;
array[51853] <= 16'b0000_0000_0000_0000;
array[51854] <= 16'b0000_0000_0000_0000;
array[51855] <= 16'b0000_0000_0000_0000;
array[51856] <= 16'b0000_0000_0000_0000;
array[51857] <= 16'b0000_0000_0000_0000;
array[51858] <= 16'b0000_0000_0000_0000;
array[51859] <= 16'b0000_0000_0000_0000;
array[51860] <= 16'b0000_0000_0000_0000;
array[51861] <= 16'b0000_0000_0000_0000;
array[51862] <= 16'b0000_0000_0000_0000;
array[51863] <= 16'b0000_0000_0000_0000;
array[51864] <= 16'b0000_0000_0000_0000;
array[51865] <= 16'b0000_0000_0000_0000;
array[51866] <= 16'b0000_0000_0000_0000;
array[51867] <= 16'b0000_0000_0000_0000;
array[51868] <= 16'b0000_0000_0000_0000;
array[51869] <= 16'b0000_0000_0000_0000;
array[51870] <= 16'b0000_0000_0000_0000;
array[51871] <= 16'b0000_0000_0000_0000;
array[51872] <= 16'b0000_0000_0000_0000;
array[51873] <= 16'b0000_0000_0000_0000;
array[51874] <= 16'b0000_0000_0000_0000;
array[51875] <= 16'b0000_0000_0000_0000;
array[51876] <= 16'b0000_0000_0000_0000;
array[51877] <= 16'b0000_0000_0000_0000;
array[51878] <= 16'b0000_0000_0000_0000;
array[51879] <= 16'b0000_0000_0000_0000;
array[51880] <= 16'b0000_0000_0000_0000;
array[51881] <= 16'b0000_0000_0000_0000;
array[51882] <= 16'b0000_0000_0000_0000;
array[51883] <= 16'b0000_0000_0000_0000;
array[51884] <= 16'b0000_0000_0000_0000;
array[51885] <= 16'b0000_0000_0000_0000;
array[51886] <= 16'b0000_0000_0000_0000;
array[51887] <= 16'b0000_0000_0000_0000;
array[51888] <= 16'b0000_0000_0000_0000;
array[51889] <= 16'b0000_0000_0000_0000;
array[51890] <= 16'b0000_0000_0000_0000;
array[51891] <= 16'b0000_0000_0000_0000;
array[51892] <= 16'b0000_0000_0000_0000;
array[51893] <= 16'b0000_0000_0000_0000;
array[51894] <= 16'b0000_0000_0000_0000;
array[51895] <= 16'b0000_0000_0000_0000;
array[51896] <= 16'b0000_0000_0000_0000;
array[51897] <= 16'b0000_0000_0000_0000;
array[51898] <= 16'b0000_0000_0000_0000;
array[51899] <= 16'b0000_0000_0000_0000;
array[51900] <= 16'b0000_0000_0000_0000;
array[51901] <= 16'b0000_0000_0000_0000;
array[51902] <= 16'b0000_0000_0000_0000;
array[51903] <= 16'b0000_0000_0000_0000;
array[51904] <= 16'b0000_0000_0000_0000;
array[51905] <= 16'b0000_0000_0000_0000;
array[51906] <= 16'b0000_0000_0000_0000;
array[51907] <= 16'b0000_0000_0000_0000;
array[51908] <= 16'b0000_0000_0000_0000;
array[51909] <= 16'b0000_0000_0000_0000;
array[51910] <= 16'b0000_0000_0000_0000;
array[51911] <= 16'b0000_0000_0000_0000;
array[51912] <= 16'b0000_0000_0000_0000;
array[51913] <= 16'b0000_0000_0000_0000;
array[51914] <= 16'b0000_0000_0000_0000;
array[51915] <= 16'b0000_0000_0000_0000;
array[51916] <= 16'b0000_0000_0000_0000;
array[51917] <= 16'b0000_0000_0000_0000;
array[51918] <= 16'b0000_0000_0000_0000;
array[51919] <= 16'b0000_0000_0000_0000;
array[51920] <= 16'b0000_0000_0000_0000;
array[51921] <= 16'b0000_0000_0000_0000;
array[51922] <= 16'b0000_0000_0000_0000;
array[51923] <= 16'b0000_0000_0000_0000;
array[51924] <= 16'b0000_0000_0000_0000;
array[51925] <= 16'b0000_0000_0000_0000;
array[51926] <= 16'b0000_0000_0000_0000;
array[51927] <= 16'b0000_0000_0000_0000;
array[51928] <= 16'b0000_0000_0000_0000;
array[51929] <= 16'b0000_0000_0000_0000;
array[51930] <= 16'b0000_0000_0000_0000;
array[51931] <= 16'b0000_0000_0000_0000;
array[51932] <= 16'b0000_0000_0000_0000;
array[51933] <= 16'b0000_0000_0000_0000;
array[51934] <= 16'b0000_0000_0000_0000;
array[51935] <= 16'b0000_0000_0000_0000;
array[51936] <= 16'b0000_0000_0000_0000;
array[51937] <= 16'b0000_0000_0000_0000;
array[51938] <= 16'b0000_0000_0000_0000;
array[51939] <= 16'b0000_0000_0000_0000;
array[51940] <= 16'b0000_0000_0000_0000;
array[51941] <= 16'b0000_0000_0000_0000;
array[51942] <= 16'b0000_0000_0000_0000;
array[51943] <= 16'b0000_0000_0000_0000;
array[51944] <= 16'b0000_0000_0000_0000;
array[51945] <= 16'b0000_0000_0000_0000;
array[51946] <= 16'b0000_0000_0000_0000;
array[51947] <= 16'b0000_0000_0000_0000;
array[51948] <= 16'b0000_0000_0000_0000;
array[51949] <= 16'b0000_0000_0000_0000;
array[51950] <= 16'b0000_0000_0000_0000;
array[51951] <= 16'b0000_0000_0000_0000;
array[51952] <= 16'b0000_0000_0000_0000;
array[51953] <= 16'b0000_0000_0000_0000;
array[51954] <= 16'b0000_0000_0000_0000;
array[51955] <= 16'b0000_0000_0000_0000;
array[51956] <= 16'b0000_0000_0000_0000;
array[51957] <= 16'b0000_0000_0000_0000;
array[51958] <= 16'b0000_0000_0000_0000;
array[51959] <= 16'b0000_0000_0000_0000;
array[51960] <= 16'b0000_0000_0000_0000;
array[51961] <= 16'b0000_0000_0000_0000;
array[51962] <= 16'b0000_0000_0000_0000;
array[51963] <= 16'b0000_0000_0000_0000;
array[51964] <= 16'b0000_0000_0000_0000;
array[51965] <= 16'b0000_0000_0000_0000;
array[51966] <= 16'b0000_0000_0000_0000;
array[51967] <= 16'b0000_0000_0000_0000;
array[51968] <= 16'b0000_0000_0000_0000;
array[51969] <= 16'b0000_0000_0000_0000;
array[51970] <= 16'b0000_0000_0000_0000;
array[51971] <= 16'b0000_0000_0000_0000;
array[51972] <= 16'b0000_0000_0000_0000;
array[51973] <= 16'b0000_0000_0000_0000;
array[51974] <= 16'b0000_0000_0000_0000;
array[51975] <= 16'b0000_0000_0000_0000;
array[51976] <= 16'b0000_0000_0000_0000;
array[51977] <= 16'b0000_0000_0000_0000;
array[51978] <= 16'b0000_0000_0000_0000;
array[51979] <= 16'b0000_0000_0000_0000;
array[51980] <= 16'b0000_0000_0000_0000;
array[51981] <= 16'b0000_0000_0000_0000;
array[51982] <= 16'b0000_0000_0000_0000;
array[51983] <= 16'b0000_0000_0000_0000;
array[51984] <= 16'b0000_0000_0000_0000;
array[51985] <= 16'b0000_0000_0000_0000;
array[51986] <= 16'b0000_0000_0000_0000;
array[51987] <= 16'b0000_0000_0000_0000;
array[51988] <= 16'b0000_0000_0000_0000;
array[51989] <= 16'b0000_0000_0000_0000;
array[51990] <= 16'b0000_0000_0000_0000;
array[51991] <= 16'b0000_0000_0000_0000;
array[51992] <= 16'b0000_0000_0000_0000;
array[51993] <= 16'b0000_0000_0000_0000;
array[51994] <= 16'b0000_0000_0000_0000;
array[51995] <= 16'b0000_0000_0000_0000;
array[51996] <= 16'b0000_0000_0000_0000;
array[51997] <= 16'b0000_0000_0000_0000;
array[51998] <= 16'b0000_0000_0000_0000;
array[51999] <= 16'b0000_0000_0000_0000;
array[52000] <= 16'b0000_0000_0000_0000;
array[52001] <= 16'b0000_0000_0000_0000;
array[52002] <= 16'b0000_0000_0000_0000;
array[52003] <= 16'b0000_0000_0000_0000;
array[52004] <= 16'b0000_0000_0000_0000;
array[52005] <= 16'b0000_0000_0000_0000;
array[52006] <= 16'b0000_0000_0000_0000;
array[52007] <= 16'b0000_0000_0000_0000;
array[52008] <= 16'b0000_0000_0000_0000;
array[52009] <= 16'b0000_0000_0000_0000;
array[52010] <= 16'b0000_0000_0000_0000;
array[52011] <= 16'b0000_0000_0000_0000;
array[52012] <= 16'b0000_0000_0000_0000;
array[52013] <= 16'b0000_0000_0000_0000;
array[52014] <= 16'b0000_0000_0000_0000;
array[52015] <= 16'b0000_0000_0000_0000;
array[52016] <= 16'b0000_0000_0000_0000;
array[52017] <= 16'b0000_0000_0000_0000;
array[52018] <= 16'b0000_0000_0000_0000;
array[52019] <= 16'b0000_0000_0000_0000;
array[52020] <= 16'b0000_0000_0000_0000;
array[52021] <= 16'b0000_0000_0000_0000;
array[52022] <= 16'b0000_0000_0000_0000;
array[52023] <= 16'b0000_0000_0000_0000;
array[52024] <= 16'b0000_0000_0000_0000;
array[52025] <= 16'b0000_0000_0000_0000;
array[52026] <= 16'b0000_0000_0000_0000;
array[52027] <= 16'b0000_0000_0000_0000;
array[52028] <= 16'b0000_0000_0000_0000;
array[52029] <= 16'b0000_0000_0000_0000;
array[52030] <= 16'b0000_0000_0000_0000;
array[52031] <= 16'b0000_0000_0000_0000;
array[52032] <= 16'b0000_0000_0000_0000;
array[52033] <= 16'b0000_0000_0000_0000;
array[52034] <= 16'b0000_0000_0000_0000;
array[52035] <= 16'b0000_0000_0000_0000;
array[52036] <= 16'b0000_0000_0000_0000;
array[52037] <= 16'b0000_0000_0000_0000;
array[52038] <= 16'b0000_0000_0000_0000;
array[52039] <= 16'b0000_0000_0000_0000;
array[52040] <= 16'b0000_0000_0000_0000;
array[52041] <= 16'b0000_0000_0000_0000;
array[52042] <= 16'b0000_0000_0000_0000;
array[52043] <= 16'b0000_0000_0000_0000;
array[52044] <= 16'b0000_0000_0000_0000;
array[52045] <= 16'b0000_0000_0000_0000;
array[52046] <= 16'b0000_0000_0000_0000;
array[52047] <= 16'b0000_0000_0000_0000;
array[52048] <= 16'b0000_0000_0000_0000;
array[52049] <= 16'b0000_0000_0000_0000;
array[52050] <= 16'b0000_0000_0000_0000;
array[52051] <= 16'b0000_0000_0000_0000;
array[52052] <= 16'b0000_0000_0000_0000;
array[52053] <= 16'b0000_0000_0000_0000;
array[52054] <= 16'b0000_0000_0000_0000;
array[52055] <= 16'b0000_0000_0000_0000;
array[52056] <= 16'b0000_0000_0000_0000;
array[52057] <= 16'b0000_0000_0000_0000;
array[52058] <= 16'b0000_0000_0000_0000;
array[52059] <= 16'b0000_0000_0000_0000;
array[52060] <= 16'b0000_0000_0000_0000;
array[52061] <= 16'b0000_0000_0000_0000;
array[52062] <= 16'b0000_0000_0000_0000;
array[52063] <= 16'b0000_0000_0000_0000;
array[52064] <= 16'b0000_0000_0000_0000;
array[52065] <= 16'b0000_0000_0000_0000;
array[52066] <= 16'b0000_0000_0000_0000;
array[52067] <= 16'b0000_0000_0000_0000;
array[52068] <= 16'b0000_0000_0000_0000;
array[52069] <= 16'b0000_0000_0000_0000;
array[52070] <= 16'b0000_0000_0000_0000;
array[52071] <= 16'b0000_0000_0000_0000;
array[52072] <= 16'b0000_0000_0000_0000;
array[52073] <= 16'b0000_0000_0000_0000;
array[52074] <= 16'b0000_0000_0000_0000;
array[52075] <= 16'b0000_0000_0000_0000;
array[52076] <= 16'b0000_0000_0000_0000;
array[52077] <= 16'b0000_0000_0000_0000;
array[52078] <= 16'b0000_0000_0000_0000;
array[52079] <= 16'b0000_0000_0000_0000;
array[52080] <= 16'b0000_0000_0000_0000;
array[52081] <= 16'b0000_0000_0000_0000;
array[52082] <= 16'b0000_0000_0000_0000;
array[52083] <= 16'b0000_0000_0000_0000;
array[52084] <= 16'b0000_0000_0000_0000;
array[52085] <= 16'b0000_0000_0000_0000;
array[52086] <= 16'b0000_0000_0000_0000;
array[52087] <= 16'b0000_0000_0000_0000;
array[52088] <= 16'b0000_0000_0000_0000;
array[52089] <= 16'b0000_0000_0000_0000;
array[52090] <= 16'b0000_0000_0000_0000;
array[52091] <= 16'b0000_0000_0000_0000;
array[52092] <= 16'b0000_0000_0000_0000;
array[52093] <= 16'b0000_0000_0000_0000;
array[52094] <= 16'b0000_0000_0000_0000;
array[52095] <= 16'b0000_0000_0000_0000;
array[52096] <= 16'b0000_0000_0000_0000;
array[52097] <= 16'b0000_0000_0000_0000;
array[52098] <= 16'b0000_0000_0000_0000;
array[52099] <= 16'b0000_0000_0000_0000;
array[52100] <= 16'b0000_0000_0000_0000;
array[52101] <= 16'b0000_0000_0000_0000;
array[52102] <= 16'b0000_0000_0000_0000;
array[52103] <= 16'b0000_0000_0000_0000;
array[52104] <= 16'b0000_0000_0000_0000;
array[52105] <= 16'b0000_0000_0000_0000;
array[52106] <= 16'b0000_0000_0000_0000;
array[52107] <= 16'b0000_0000_0000_0000;
array[52108] <= 16'b0000_0000_0000_0000;
array[52109] <= 16'b0000_0000_0000_0000;
array[52110] <= 16'b0000_0000_0000_0000;
array[52111] <= 16'b0000_0000_0000_0000;
array[52112] <= 16'b0000_0000_0000_0000;
array[52113] <= 16'b0000_0000_0000_0000;
array[52114] <= 16'b0000_0000_0000_0000;
array[52115] <= 16'b0000_0000_0000_0000;
array[52116] <= 16'b0000_0000_0000_0000;
array[52117] <= 16'b0000_0000_0000_0000;
array[52118] <= 16'b0000_0000_0000_0000;
array[52119] <= 16'b0000_0000_0000_0000;
array[52120] <= 16'b0000_0000_0000_0000;
array[52121] <= 16'b0000_0000_0000_0000;
array[52122] <= 16'b0000_0000_0000_0000;
array[52123] <= 16'b0000_0000_0000_0000;
array[52124] <= 16'b0000_0000_0000_0000;
array[52125] <= 16'b0000_0000_0000_0000;
array[52126] <= 16'b0000_0000_0000_0000;
array[52127] <= 16'b0000_0000_0000_0000;
array[52128] <= 16'b0000_0000_0000_0000;
array[52129] <= 16'b0000_0000_0000_0000;
array[52130] <= 16'b0000_0000_0000_0000;
array[52131] <= 16'b0000_0000_0000_0000;
array[52132] <= 16'b0000_0000_0000_0000;
array[52133] <= 16'b0000_0000_0000_0000;
array[52134] <= 16'b0000_0000_0000_0000;
array[52135] <= 16'b0000_0000_0000_0000;
array[52136] <= 16'b0000_0000_0000_0000;
array[52137] <= 16'b0000_0000_0000_0000;
array[52138] <= 16'b0000_0000_0000_0000;
array[52139] <= 16'b0000_0000_0000_0000;
array[52140] <= 16'b0000_0000_0000_0000;
array[52141] <= 16'b0000_0000_0000_0000;
array[52142] <= 16'b0000_0000_0000_0000;
array[52143] <= 16'b0000_0000_0000_0000;
array[52144] <= 16'b0000_0000_0000_0000;
array[52145] <= 16'b0000_0000_0000_0000;
array[52146] <= 16'b0000_0000_0000_0000;
array[52147] <= 16'b0000_0000_0000_0000;
array[52148] <= 16'b0000_0000_0000_0000;
array[52149] <= 16'b0000_0000_0000_0000;
array[52150] <= 16'b0000_0000_0000_0000;
array[52151] <= 16'b0000_0000_0000_0000;
array[52152] <= 16'b0000_0000_0000_0000;
array[52153] <= 16'b0000_0000_0000_0000;
array[52154] <= 16'b0000_0000_0000_0000;
array[52155] <= 16'b0000_0000_0000_0000;
array[52156] <= 16'b0000_0000_0000_0000;
array[52157] <= 16'b0000_0000_0000_0000;
array[52158] <= 16'b0000_0000_0000_0000;
array[52159] <= 16'b0000_0000_0000_0000;
array[52160] <= 16'b0000_0000_0000_0000;
array[52161] <= 16'b0000_0000_0000_0000;
array[52162] <= 16'b0000_0000_0000_0000;
array[52163] <= 16'b0000_0000_0000_0000;
array[52164] <= 16'b0000_0000_0000_0000;
array[52165] <= 16'b0000_0000_0000_0000;
array[52166] <= 16'b0000_0000_0000_0000;
array[52167] <= 16'b0000_0000_0000_0000;
array[52168] <= 16'b0000_0000_0000_0000;
array[52169] <= 16'b0000_0000_0000_0000;
array[52170] <= 16'b0000_0000_0000_0000;
array[52171] <= 16'b0000_0000_0000_0000;
array[52172] <= 16'b0000_0000_0000_0000;
array[52173] <= 16'b0000_0000_0000_0000;
array[52174] <= 16'b0000_0000_0000_0000;
array[52175] <= 16'b0000_0000_0000_0000;
array[52176] <= 16'b0000_0000_0000_0000;
array[52177] <= 16'b0000_0000_0000_0000;
array[52178] <= 16'b0000_0000_0000_0000;
array[52179] <= 16'b0000_0000_0000_0000;
array[52180] <= 16'b0000_0000_0000_0000;
array[52181] <= 16'b0000_0000_0000_0000;
array[52182] <= 16'b0000_0000_0000_0000;
array[52183] <= 16'b0000_0000_0000_0000;
array[52184] <= 16'b0000_0000_0000_0000;
array[52185] <= 16'b0000_0000_0000_0000;
array[52186] <= 16'b0000_0000_0000_0000;
array[52187] <= 16'b0000_0000_0000_0000;
array[52188] <= 16'b0000_0000_0000_0000;
array[52189] <= 16'b0000_0000_0000_0000;
array[52190] <= 16'b0000_0000_0000_0000;
array[52191] <= 16'b0000_0000_0000_0000;
array[52192] <= 16'b0000_0000_0000_0000;
array[52193] <= 16'b0000_0000_0000_0000;
array[52194] <= 16'b0000_0000_0000_0000;
array[52195] <= 16'b0000_0000_0000_0000;
array[52196] <= 16'b0000_0000_0000_0000;
array[52197] <= 16'b0000_0000_0000_0000;
array[52198] <= 16'b0000_0000_0000_0000;
array[52199] <= 16'b0000_0000_0000_0000;
array[52200] <= 16'b0000_0000_0000_0000;
array[52201] <= 16'b0000_0000_0000_0000;
array[52202] <= 16'b0000_0000_0000_0000;
array[52203] <= 16'b0000_0000_0000_0000;
array[52204] <= 16'b0000_0000_0000_0000;
array[52205] <= 16'b0000_0000_0000_0000;
array[52206] <= 16'b0000_0000_0000_0000;
array[52207] <= 16'b0000_0000_0000_0000;
array[52208] <= 16'b0000_0000_0000_0000;
array[52209] <= 16'b0000_0000_0000_0000;
array[52210] <= 16'b0000_0000_0000_0000;
array[52211] <= 16'b0000_0000_0000_0000;
array[52212] <= 16'b0000_0000_0000_0000;
array[52213] <= 16'b0000_0000_0000_0000;
array[52214] <= 16'b0000_0000_0000_0000;
array[52215] <= 16'b0000_0000_0000_0000;
array[52216] <= 16'b0000_0000_0000_0000;
array[52217] <= 16'b0000_0000_0000_0000;
array[52218] <= 16'b0000_0000_0000_0000;
array[52219] <= 16'b0000_0000_0000_0000;
array[52220] <= 16'b0000_0000_0000_0000;
array[52221] <= 16'b0000_0000_0000_0000;
array[52222] <= 16'b0000_0000_0000_0000;
array[52223] <= 16'b0000_0000_0000_0000;
array[52224] <= 16'b0000_0000_0000_0000;
array[52225] <= 16'b0000_0000_0000_0000;
array[52226] <= 16'b0000_0000_0000_0000;
array[52227] <= 16'b0000_0000_0000_0000;
array[52228] <= 16'b0000_0000_0000_0000;
array[52229] <= 16'b0000_0000_0000_0000;
array[52230] <= 16'b0000_0000_0000_0000;
array[52231] <= 16'b0000_0000_0000_0000;
array[52232] <= 16'b0000_0000_0000_0000;
array[52233] <= 16'b0000_0000_0000_0000;
array[52234] <= 16'b0000_0000_0000_0000;
array[52235] <= 16'b0000_0000_0000_0000;
array[52236] <= 16'b0000_0000_0000_0000;
array[52237] <= 16'b0000_0000_0000_0000;
array[52238] <= 16'b0000_0000_0000_0000;
array[52239] <= 16'b0000_0000_0000_0000;
array[52240] <= 16'b0000_0000_0000_0000;
array[52241] <= 16'b0000_0000_0000_0000;
array[52242] <= 16'b0000_0000_0000_0000;
array[52243] <= 16'b0000_0000_0000_0000;
array[52244] <= 16'b0000_0000_0000_0000;
array[52245] <= 16'b0000_0000_0000_0000;
array[52246] <= 16'b0000_0000_0000_0000;
array[52247] <= 16'b0000_0000_0000_0000;
array[52248] <= 16'b0000_0000_0000_0000;
array[52249] <= 16'b0000_0000_0000_0000;
array[52250] <= 16'b0000_0000_0000_0000;
array[52251] <= 16'b0000_0000_0000_0000;
array[52252] <= 16'b0000_0000_0000_0000;
array[52253] <= 16'b0000_0000_0000_0000;
array[52254] <= 16'b0000_0000_0000_0000;
array[52255] <= 16'b0000_0000_0000_0000;
array[52256] <= 16'b0000_0000_0000_0000;
array[52257] <= 16'b0000_0000_0000_0000;
array[52258] <= 16'b0000_0000_0000_0000;
array[52259] <= 16'b0000_0000_0000_0000;
array[52260] <= 16'b0000_0000_0000_0000;
array[52261] <= 16'b0000_0000_0000_0000;
array[52262] <= 16'b0000_0000_0000_0000;
array[52263] <= 16'b0000_0000_0000_0000;
array[52264] <= 16'b0000_0000_0000_0000;
array[52265] <= 16'b0000_0000_0000_0000;
array[52266] <= 16'b0000_0000_0000_0000;
array[52267] <= 16'b0000_0000_0000_0000;
array[52268] <= 16'b0000_0000_0000_0000;
array[52269] <= 16'b0000_0000_0000_0000;
array[52270] <= 16'b0000_0000_0000_0000;
array[52271] <= 16'b0000_0000_0000_0000;
array[52272] <= 16'b0000_0000_0000_0000;
array[52273] <= 16'b0000_0000_0000_0000;
array[52274] <= 16'b0000_0000_0000_0000;
array[52275] <= 16'b0000_0000_0000_0000;
array[52276] <= 16'b0000_0000_0000_0000;
array[52277] <= 16'b0000_0000_0000_0000;
array[52278] <= 16'b0000_0000_0000_0000;
array[52279] <= 16'b0000_0000_0000_0000;
array[52280] <= 16'b0000_0000_0000_0000;
array[52281] <= 16'b0000_0000_0000_0000;
array[52282] <= 16'b0000_0000_0000_0000;
array[52283] <= 16'b0000_0000_0000_0000;
array[52284] <= 16'b0000_0000_0000_0000;
array[52285] <= 16'b0000_0000_0000_0000;
array[52286] <= 16'b0000_0000_0000_0000;
array[52287] <= 16'b0000_0000_0000_0000;
array[52288] <= 16'b0000_0000_0000_0000;
array[52289] <= 16'b0000_0000_0000_0000;
array[52290] <= 16'b0000_0000_0000_0000;
array[52291] <= 16'b0000_0000_0000_0000;
array[52292] <= 16'b0000_0000_0000_0000;
array[52293] <= 16'b0000_0000_0000_0000;
array[52294] <= 16'b0000_0000_0000_0000;
array[52295] <= 16'b0000_0000_0000_0000;
array[52296] <= 16'b0000_0000_0000_0000;
array[52297] <= 16'b0000_0000_0000_0000;
array[52298] <= 16'b0000_0000_0000_0000;
array[52299] <= 16'b0000_0000_0000_0000;
array[52300] <= 16'b0000_0000_0000_0000;
array[52301] <= 16'b0000_0000_0000_0000;
array[52302] <= 16'b0000_0000_0000_0000;
array[52303] <= 16'b0000_0000_0000_0000;
array[52304] <= 16'b0000_0000_0000_0000;
array[52305] <= 16'b0000_0000_0000_0000;
array[52306] <= 16'b0000_0000_0000_0000;
array[52307] <= 16'b0000_0000_0000_0000;
array[52308] <= 16'b0000_0000_0000_0000;
array[52309] <= 16'b0000_0000_0000_0000;
array[52310] <= 16'b0000_0000_0000_0000;
array[52311] <= 16'b0000_0000_0000_0000;
array[52312] <= 16'b0000_0000_0000_0000;
array[52313] <= 16'b0000_0000_0000_0000;
array[52314] <= 16'b0000_0000_0000_0000;
array[52315] <= 16'b0000_0000_0000_0000;
array[52316] <= 16'b0000_0000_0000_0000;
array[52317] <= 16'b0000_0000_0000_0000;
array[52318] <= 16'b0000_0000_0000_0000;
array[52319] <= 16'b0000_0000_0000_0000;
array[52320] <= 16'b0000_0000_0000_0000;
array[52321] <= 16'b0000_0000_0000_0000;
array[52322] <= 16'b0000_0000_0000_0000;
array[52323] <= 16'b0000_0000_0000_0000;
array[52324] <= 16'b0000_0000_0000_0000;
array[52325] <= 16'b0000_0000_0000_0000;
array[52326] <= 16'b0000_0000_0000_0000;
array[52327] <= 16'b0000_0000_0000_0000;
array[52328] <= 16'b0000_0000_0000_0000;
array[52329] <= 16'b0000_0000_0000_0000;
array[52330] <= 16'b0000_0000_0000_0000;
array[52331] <= 16'b0000_0000_0000_0000;
array[52332] <= 16'b0000_0000_0000_0000;
array[52333] <= 16'b0000_0000_0000_0000;
array[52334] <= 16'b0000_0000_0000_0000;
array[52335] <= 16'b0000_0000_0000_0000;
array[52336] <= 16'b0000_0000_0000_0000;
array[52337] <= 16'b0000_0000_0000_0000;
array[52338] <= 16'b0000_0000_0000_0000;
array[52339] <= 16'b0000_0000_0000_0000;
array[52340] <= 16'b0000_0000_0000_0000;
array[52341] <= 16'b0000_0000_0000_0000;
array[52342] <= 16'b0000_0000_0000_0000;
array[52343] <= 16'b0000_0000_0000_0000;
array[52344] <= 16'b0000_0000_0000_0000;
array[52345] <= 16'b0000_0000_0000_0000;
array[52346] <= 16'b0000_0000_0000_0000;
array[52347] <= 16'b0000_0000_0000_0000;
array[52348] <= 16'b0000_0000_0000_0000;
array[52349] <= 16'b0000_0000_0000_0000;
array[52350] <= 16'b0000_0000_0000_0000;
array[52351] <= 16'b0000_0000_0000_0000;
array[52352] <= 16'b0000_0000_0000_0000;
array[52353] <= 16'b0000_0000_0000_0000;
array[52354] <= 16'b0000_0000_0000_0000;
array[52355] <= 16'b0000_0000_0000_0000;
array[52356] <= 16'b0000_0000_0000_0000;
array[52357] <= 16'b0000_0000_0000_0000;
array[52358] <= 16'b0000_0000_0000_0000;
array[52359] <= 16'b0000_0000_0000_0000;
array[52360] <= 16'b0000_0000_0000_0000;
array[52361] <= 16'b0000_0000_0000_0000;
array[52362] <= 16'b0000_0000_0000_0000;
array[52363] <= 16'b0000_0000_0000_0000;
array[52364] <= 16'b0000_0000_0000_0000;
array[52365] <= 16'b0000_0000_0000_0000;
array[52366] <= 16'b0000_0000_0000_0000;
array[52367] <= 16'b0000_0000_0000_0000;
array[52368] <= 16'b0000_0000_0000_0000;
array[52369] <= 16'b0000_0000_0000_0000;
array[52370] <= 16'b0000_0000_0000_0000;
array[52371] <= 16'b0000_0000_0000_0000;
array[52372] <= 16'b0000_0000_0000_0000;
array[52373] <= 16'b0000_0000_0000_0000;
array[52374] <= 16'b0000_0000_0000_0000;
array[52375] <= 16'b0000_0000_0000_0000;
array[52376] <= 16'b0000_0000_0000_0000;
array[52377] <= 16'b0000_0000_0000_0000;
array[52378] <= 16'b0000_0000_0000_0000;
array[52379] <= 16'b0000_0000_0000_0000;
array[52380] <= 16'b0000_0000_0000_0000;
array[52381] <= 16'b0000_0000_0000_0000;
array[52382] <= 16'b0000_0000_0000_0000;
array[52383] <= 16'b0000_0000_0000_0000;
array[52384] <= 16'b0000_0000_0000_0000;
array[52385] <= 16'b0000_0000_0000_0000;
array[52386] <= 16'b0000_0000_0000_0000;
array[52387] <= 16'b0000_0000_0000_0000;
array[52388] <= 16'b0000_0000_0000_0000;
array[52389] <= 16'b0000_0000_0000_0000;
array[52390] <= 16'b0000_0000_0000_0000;
array[52391] <= 16'b0000_0000_0000_0000;
array[52392] <= 16'b0000_0000_0000_0000;
array[52393] <= 16'b0000_0000_0000_0000;
array[52394] <= 16'b0000_0000_0000_0000;
array[52395] <= 16'b0000_0000_0000_0000;
array[52396] <= 16'b0000_0000_0000_0000;
array[52397] <= 16'b0000_0000_0000_0000;
array[52398] <= 16'b0000_0000_0000_0000;
array[52399] <= 16'b0000_0000_0000_0000;
array[52400] <= 16'b0000_0000_0000_0000;
array[52401] <= 16'b0000_0000_0000_0000;
array[52402] <= 16'b0000_0000_0000_0000;
array[52403] <= 16'b0000_0000_0000_0000;
array[52404] <= 16'b0000_0000_0000_0000;
array[52405] <= 16'b0000_0000_0000_0000;
array[52406] <= 16'b0000_0000_0000_0000;
array[52407] <= 16'b0000_0000_0000_0000;
array[52408] <= 16'b0000_0000_0000_0000;
array[52409] <= 16'b0000_0000_0000_0000;
array[52410] <= 16'b0000_0000_0000_0000;
array[52411] <= 16'b0000_0000_0000_0000;
array[52412] <= 16'b0000_0000_0000_0000;
array[52413] <= 16'b0000_0000_0000_0000;
array[52414] <= 16'b0000_0000_0000_0000;
array[52415] <= 16'b0000_0000_0000_0000;
array[52416] <= 16'b0000_0000_0000_0000;
array[52417] <= 16'b0000_0000_0000_0000;
array[52418] <= 16'b0000_0000_0000_0000;
array[52419] <= 16'b0000_0000_0000_0000;
array[52420] <= 16'b0000_0000_0000_0000;
array[52421] <= 16'b0000_0000_0000_0000;
array[52422] <= 16'b0000_0000_0000_0000;
array[52423] <= 16'b0000_0000_0000_0000;
array[52424] <= 16'b0000_0000_0000_0000;
array[52425] <= 16'b0000_0000_0000_0000;
array[52426] <= 16'b0000_0000_0000_0000;
array[52427] <= 16'b0000_0000_0000_0000;
array[52428] <= 16'b0000_0000_0000_0000;
array[52429] <= 16'b0000_0000_0000_0000;
array[52430] <= 16'b0000_0000_0000_0000;
array[52431] <= 16'b0000_0000_0000_0000;
array[52432] <= 16'b0000_0000_0000_0000;
array[52433] <= 16'b0000_0000_0000_0000;
array[52434] <= 16'b0000_0000_0000_0000;
array[52435] <= 16'b0000_0000_0000_0000;
array[52436] <= 16'b0000_0000_0000_0000;
array[52437] <= 16'b0000_0000_0000_0000;
array[52438] <= 16'b0000_0000_0000_0000;
array[52439] <= 16'b0000_0000_0000_0000;
array[52440] <= 16'b0000_0000_0000_0000;
array[52441] <= 16'b0000_0000_0000_0000;
array[52442] <= 16'b0000_0000_0000_0000;
array[52443] <= 16'b0000_0000_0000_0000;
array[52444] <= 16'b0000_0000_0000_0000;
array[52445] <= 16'b0000_0000_0000_0000;
array[52446] <= 16'b0000_0000_0000_0000;
array[52447] <= 16'b0000_0000_0000_0000;
array[52448] <= 16'b0000_0000_0000_0000;
array[52449] <= 16'b0000_0000_0000_0000;
array[52450] <= 16'b0000_0000_0000_0000;
array[52451] <= 16'b0000_0000_0000_0000;
array[52452] <= 16'b0000_0000_0000_0000;
array[52453] <= 16'b0000_0000_0000_0000;
array[52454] <= 16'b0000_0000_0000_0000;
array[52455] <= 16'b0000_0000_0000_0000;
array[52456] <= 16'b0000_0000_0000_0000;
array[52457] <= 16'b0000_0000_0000_0000;
array[52458] <= 16'b0000_0000_0000_0000;
array[52459] <= 16'b0000_0000_0000_0000;
array[52460] <= 16'b0000_0000_0000_0000;
array[52461] <= 16'b0000_0000_0000_0000;
array[52462] <= 16'b0000_0000_0000_0000;
array[52463] <= 16'b0000_0000_0000_0000;
array[52464] <= 16'b0000_0000_0000_0000;
array[52465] <= 16'b0000_0000_0000_0000;
array[52466] <= 16'b0000_0000_0000_0000;
array[52467] <= 16'b0000_0000_0000_0000;
array[52468] <= 16'b0000_0000_0000_0000;
array[52469] <= 16'b0000_0000_0000_0000;
array[52470] <= 16'b0000_0000_0000_0000;
array[52471] <= 16'b0000_0000_0000_0000;
array[52472] <= 16'b0000_0000_0000_0000;
array[52473] <= 16'b0000_0000_0000_0000;
array[52474] <= 16'b0000_0000_0000_0000;
array[52475] <= 16'b0000_0000_0000_0000;
array[52476] <= 16'b0000_0000_0000_0000;
array[52477] <= 16'b0000_0000_0000_0000;
array[52478] <= 16'b0000_0000_0000_0000;
array[52479] <= 16'b0000_0000_0000_0000;
array[52480] <= 16'b0000_0000_0000_0000;
array[52481] <= 16'b0000_0000_0000_0000;
array[52482] <= 16'b0000_0000_0000_0000;
array[52483] <= 16'b0000_0000_0000_0000;
array[52484] <= 16'b0000_0000_0000_0000;
array[52485] <= 16'b0000_0000_0000_0000;
array[52486] <= 16'b0000_0000_0000_0000;
array[52487] <= 16'b0000_0000_0000_0000;
array[52488] <= 16'b0000_0000_0000_0000;
array[52489] <= 16'b0000_0000_0000_0000;
array[52490] <= 16'b0000_0000_0000_0000;
array[52491] <= 16'b0000_0000_0000_0000;
array[52492] <= 16'b0000_0000_0000_0000;
array[52493] <= 16'b0000_0000_0000_0000;
array[52494] <= 16'b0000_0000_0000_0000;
array[52495] <= 16'b0000_0000_0000_0000;
array[52496] <= 16'b0000_0000_0000_0000;
array[52497] <= 16'b0000_0000_0000_0000;
array[52498] <= 16'b0000_0000_0000_0000;
array[52499] <= 16'b0000_0000_0000_0000;
array[52500] <= 16'b0000_0000_0000_0000;
array[52501] <= 16'b0000_0000_0000_0000;
array[52502] <= 16'b0000_0000_0000_0000;
array[52503] <= 16'b0000_0000_0000_0000;
array[52504] <= 16'b0000_0000_0000_0000;
array[52505] <= 16'b0000_0000_0000_0000;
array[52506] <= 16'b0000_0000_0000_0000;
array[52507] <= 16'b0000_0000_0000_0000;
array[52508] <= 16'b0000_0000_0000_0000;
array[52509] <= 16'b0000_0000_0000_0000;
array[52510] <= 16'b0000_0000_0000_0000;
array[52511] <= 16'b0000_0000_0000_0000;
array[52512] <= 16'b0000_0000_0000_0000;
array[52513] <= 16'b0000_0000_0000_0000;
array[52514] <= 16'b0000_0000_0000_0000;
array[52515] <= 16'b0000_0000_0000_0000;
array[52516] <= 16'b0000_0000_0000_0000;
array[52517] <= 16'b0000_0000_0000_0000;
array[52518] <= 16'b0000_0000_0000_0000;
array[52519] <= 16'b0000_0000_0000_0000;
array[52520] <= 16'b0000_0000_0000_0000;
array[52521] <= 16'b0000_0000_0000_0000;
array[52522] <= 16'b0000_0000_0000_0000;
array[52523] <= 16'b0000_0000_0000_0000;
array[52524] <= 16'b0000_0000_0000_0000;
array[52525] <= 16'b0000_0000_0000_0000;
array[52526] <= 16'b0000_0000_0000_0000;
array[52527] <= 16'b0000_0000_0000_0000;
array[52528] <= 16'b0000_0000_0000_0000;
array[52529] <= 16'b0000_0000_0000_0000;
array[52530] <= 16'b0000_0000_0000_0000;
array[52531] <= 16'b0000_0000_0000_0000;
array[52532] <= 16'b0000_0000_0000_0000;
array[52533] <= 16'b0000_0000_0000_0000;
array[52534] <= 16'b0000_0000_0000_0000;
array[52535] <= 16'b0000_0000_0000_0000;
array[52536] <= 16'b0000_0000_0000_0000;
array[52537] <= 16'b0000_0000_0000_0000;
array[52538] <= 16'b0000_0000_0000_0000;
array[52539] <= 16'b0000_0000_0000_0000;
array[52540] <= 16'b0000_0000_0000_0000;
array[52541] <= 16'b0000_0000_0000_0000;
array[52542] <= 16'b0000_0000_0000_0000;
array[52543] <= 16'b0000_0000_0000_0000;
array[52544] <= 16'b0000_0000_0000_0000;
array[52545] <= 16'b0000_0000_0000_0000;
array[52546] <= 16'b0000_0000_0000_0000;
array[52547] <= 16'b0000_0000_0000_0000;
array[52548] <= 16'b0000_0000_0000_0000;
array[52549] <= 16'b0000_0000_0000_0000;
array[52550] <= 16'b0000_0000_0000_0000;
array[52551] <= 16'b0000_0000_0000_0000;
array[52552] <= 16'b0000_0000_0000_0000;
array[52553] <= 16'b0000_0000_0000_0000;
array[52554] <= 16'b0000_0000_0000_0000;
array[52555] <= 16'b0000_0000_0000_0000;
array[52556] <= 16'b0000_0000_0000_0000;
array[52557] <= 16'b0000_0000_0000_0000;
array[52558] <= 16'b0000_0000_0000_0000;
array[52559] <= 16'b0000_0000_0000_0000;
array[52560] <= 16'b0000_0000_0000_0000;
array[52561] <= 16'b0000_0000_0000_0000;
array[52562] <= 16'b0000_0000_0000_0000;
array[52563] <= 16'b0000_0000_0000_0000;
array[52564] <= 16'b0000_0000_0000_0000;
array[52565] <= 16'b0000_0000_0000_0000;
array[52566] <= 16'b0000_0000_0000_0000;
array[52567] <= 16'b0000_0000_0000_0000;
array[52568] <= 16'b0000_0000_0000_0000;
array[52569] <= 16'b0000_0000_0000_0000;
array[52570] <= 16'b0000_0000_0000_0000;
array[52571] <= 16'b0000_0000_0000_0000;
array[52572] <= 16'b0000_0000_0000_0000;
array[52573] <= 16'b0000_0000_0000_0000;
array[52574] <= 16'b0000_0000_0000_0000;
array[52575] <= 16'b0000_0000_0000_0000;
array[52576] <= 16'b0000_0000_0000_0000;
array[52577] <= 16'b0000_0000_0000_0000;
array[52578] <= 16'b0000_0000_0000_0000;
array[52579] <= 16'b0000_0000_0000_0000;
array[52580] <= 16'b0000_0000_0000_0000;
array[52581] <= 16'b0000_0000_0000_0000;
array[52582] <= 16'b0000_0000_0000_0000;
array[52583] <= 16'b0000_0000_0000_0000;
array[52584] <= 16'b0000_0000_0000_0000;
array[52585] <= 16'b0000_0000_0000_0000;
array[52586] <= 16'b0000_0000_0000_0000;
array[52587] <= 16'b0000_0000_0000_0000;
array[52588] <= 16'b0000_0000_0000_0000;
array[52589] <= 16'b0000_0000_0000_0000;
array[52590] <= 16'b0000_0000_0000_0000;
array[52591] <= 16'b0000_0000_0000_0000;
array[52592] <= 16'b0000_0000_0000_0000;
array[52593] <= 16'b0000_0000_0000_0000;
array[52594] <= 16'b0000_0000_0000_0000;
array[52595] <= 16'b0000_0000_0000_0000;
array[52596] <= 16'b0000_0000_0000_0000;
array[52597] <= 16'b0000_0000_0000_0000;
array[52598] <= 16'b0000_0000_0000_0000;
array[52599] <= 16'b0000_0000_0000_0000;
array[52600] <= 16'b0000_0000_0000_0000;
array[52601] <= 16'b0000_0000_0000_0000;
array[52602] <= 16'b0000_0000_0000_0000;
array[52603] <= 16'b0000_0000_0000_0000;
array[52604] <= 16'b0000_0000_0000_0000;
array[52605] <= 16'b0000_0000_0000_0000;
array[52606] <= 16'b0000_0000_0000_0000;
array[52607] <= 16'b0000_0000_0000_0000;
array[52608] <= 16'b0000_0000_0000_0000;
array[52609] <= 16'b0000_0000_0000_0000;
array[52610] <= 16'b0000_0000_0000_0000;
array[52611] <= 16'b0000_0000_0000_0000;
array[52612] <= 16'b0000_0000_0000_0000;
array[52613] <= 16'b0000_0000_0000_0000;
array[52614] <= 16'b0000_0000_0000_0000;
array[52615] <= 16'b0000_0000_0000_0000;
array[52616] <= 16'b0000_0000_0000_0000;
array[52617] <= 16'b0000_0000_0000_0000;
array[52618] <= 16'b0000_0000_0000_0000;
array[52619] <= 16'b0000_0000_0000_0000;
array[52620] <= 16'b0000_0000_0000_0000;
array[52621] <= 16'b0000_0000_0000_0000;
array[52622] <= 16'b0000_0000_0000_0000;
array[52623] <= 16'b0000_0000_0000_0000;
array[52624] <= 16'b0000_0000_0000_0000;
array[52625] <= 16'b0000_0000_0000_0000;
array[52626] <= 16'b0000_0000_0000_0000;
array[52627] <= 16'b0000_0000_0000_0000;
array[52628] <= 16'b0000_0000_0000_0000;
array[52629] <= 16'b0000_0000_0000_0000;
array[52630] <= 16'b0000_0000_0000_0000;
array[52631] <= 16'b0000_0000_0000_0000;
array[52632] <= 16'b0000_0000_0000_0000;
array[52633] <= 16'b0000_0000_0000_0000;
array[52634] <= 16'b0000_0000_0000_0000;
array[52635] <= 16'b0000_0000_0000_0000;
array[52636] <= 16'b0000_0000_0000_0000;
array[52637] <= 16'b0000_0000_0000_0000;
array[52638] <= 16'b0000_0000_0000_0000;
array[52639] <= 16'b0000_0000_0000_0000;
array[52640] <= 16'b0000_0000_0000_0000;
array[52641] <= 16'b0000_0000_0000_0000;
array[52642] <= 16'b0000_0000_0000_0000;
array[52643] <= 16'b0000_0000_0000_0000;
array[52644] <= 16'b0000_0000_0000_0000;
array[52645] <= 16'b0000_0000_0000_0000;
array[52646] <= 16'b0000_0000_0000_0000;
array[52647] <= 16'b0000_0000_0000_0000;
array[52648] <= 16'b0000_0000_0000_0000;
array[52649] <= 16'b0000_0000_0000_0000;
array[52650] <= 16'b0000_0000_0000_0000;
array[52651] <= 16'b0000_0000_0000_0000;
array[52652] <= 16'b0000_0000_0000_0000;
array[52653] <= 16'b0000_0000_0000_0000;
array[52654] <= 16'b0000_0000_0000_0000;
array[52655] <= 16'b0000_0000_0000_0000;
array[52656] <= 16'b0000_0000_0000_0000;
array[52657] <= 16'b0000_0000_0000_0000;
array[52658] <= 16'b0000_0000_0000_0000;
array[52659] <= 16'b0000_0000_0000_0000;
array[52660] <= 16'b0000_0000_0000_0000;
array[52661] <= 16'b0000_0000_0000_0000;
array[52662] <= 16'b0000_0000_0000_0000;
array[52663] <= 16'b0000_0000_0000_0000;
array[52664] <= 16'b0000_0000_0000_0000;
array[52665] <= 16'b0000_0000_0000_0000;
array[52666] <= 16'b0000_0000_0000_0000;
array[52667] <= 16'b0000_0000_0000_0000;
array[52668] <= 16'b0000_0000_0000_0000;
array[52669] <= 16'b0000_0000_0000_0000;
array[52670] <= 16'b0000_0000_0000_0000;
array[52671] <= 16'b0000_0000_0000_0000;
array[52672] <= 16'b0000_0000_0000_0000;
array[52673] <= 16'b0000_0000_0000_0000;
array[52674] <= 16'b0000_0000_0000_0000;
array[52675] <= 16'b0000_0000_0000_0000;
array[52676] <= 16'b0000_0000_0000_0000;
array[52677] <= 16'b0000_0000_0000_0000;
array[52678] <= 16'b0000_0000_0000_0000;
array[52679] <= 16'b0000_0000_0000_0000;
array[52680] <= 16'b0000_0000_0000_0000;
array[52681] <= 16'b0000_0000_0000_0000;
array[52682] <= 16'b0000_0000_0000_0000;
array[52683] <= 16'b0000_0000_0000_0000;
array[52684] <= 16'b0000_0000_0000_0000;
array[52685] <= 16'b0000_0000_0000_0000;
array[52686] <= 16'b0000_0000_0000_0000;
array[52687] <= 16'b0000_0000_0000_0000;
array[52688] <= 16'b0000_0000_0000_0000;
array[52689] <= 16'b0000_0000_0000_0000;
array[52690] <= 16'b0000_0000_0000_0000;
array[52691] <= 16'b0000_0000_0000_0000;
array[52692] <= 16'b0000_0000_0000_0000;
array[52693] <= 16'b0000_0000_0000_0000;
array[52694] <= 16'b0000_0000_0000_0000;
array[52695] <= 16'b0000_0000_0000_0000;
array[52696] <= 16'b0000_0000_0000_0000;
array[52697] <= 16'b0000_0000_0000_0000;
array[52698] <= 16'b0000_0000_0000_0000;
array[52699] <= 16'b0000_0000_0000_0000;
array[52700] <= 16'b0000_0000_0000_0000;
array[52701] <= 16'b0000_0000_0000_0000;
array[52702] <= 16'b0000_0000_0000_0000;
array[52703] <= 16'b0000_0000_0000_0000;
array[52704] <= 16'b0000_0000_0000_0000;
array[52705] <= 16'b0000_0000_0000_0000;
array[52706] <= 16'b0000_0000_0000_0000;
array[52707] <= 16'b0000_0000_0000_0000;
array[52708] <= 16'b0000_0000_0000_0000;
array[52709] <= 16'b0000_0000_0000_0000;
array[52710] <= 16'b0000_0000_0000_0000;
array[52711] <= 16'b0000_0000_0000_0000;
array[52712] <= 16'b0000_0000_0000_0000;
array[52713] <= 16'b0000_0000_0000_0000;
array[52714] <= 16'b0000_0000_0000_0000;
array[52715] <= 16'b0000_0000_0000_0000;
array[52716] <= 16'b0000_0000_0000_0000;
array[52717] <= 16'b0000_0000_0000_0000;
array[52718] <= 16'b0000_0000_0000_0000;
array[52719] <= 16'b0000_0000_0000_0000;
array[52720] <= 16'b0000_0000_0000_0000;
array[52721] <= 16'b0000_0000_0000_0000;
array[52722] <= 16'b0000_0000_0000_0000;
array[52723] <= 16'b0000_0000_0000_0000;
array[52724] <= 16'b0000_0000_0000_0000;
array[52725] <= 16'b0000_0000_0000_0000;
array[52726] <= 16'b0000_0000_0000_0000;
array[52727] <= 16'b0000_0000_0000_0000;
array[52728] <= 16'b0000_0000_0000_0000;
array[52729] <= 16'b0000_0000_0000_0000;
array[52730] <= 16'b0000_0000_0000_0000;
array[52731] <= 16'b0000_0000_0000_0000;
array[52732] <= 16'b0000_0000_0000_0000;
array[52733] <= 16'b0000_0000_0000_0000;
array[52734] <= 16'b0000_0000_0000_0000;
array[52735] <= 16'b0000_0000_0000_0000;
array[52736] <= 16'b0000_0000_0000_0000;
array[52737] <= 16'b0000_0000_0000_0000;
array[52738] <= 16'b0000_0000_0000_0000;
array[52739] <= 16'b0000_0000_0000_0000;
array[52740] <= 16'b0000_0000_0000_0000;
array[52741] <= 16'b0000_0000_0000_0000;
array[52742] <= 16'b0000_0000_0000_0000;
array[52743] <= 16'b0000_0000_0000_0000;
array[52744] <= 16'b0000_0000_0000_0000;
array[52745] <= 16'b0000_0000_0000_0000;
array[52746] <= 16'b0000_0000_0000_0000;
array[52747] <= 16'b0000_0000_0000_0000;
array[52748] <= 16'b0000_0000_0000_0000;
array[52749] <= 16'b0000_0000_0000_0000;
array[52750] <= 16'b0000_0000_0000_0000;
array[52751] <= 16'b0000_0000_0000_0000;
array[52752] <= 16'b0000_0000_0000_0000;
array[52753] <= 16'b0000_0000_0000_0000;
array[52754] <= 16'b0000_0000_0000_0000;
array[52755] <= 16'b0000_0000_0000_0000;
array[52756] <= 16'b0000_0000_0000_0000;
array[52757] <= 16'b0000_0000_0000_0000;
array[52758] <= 16'b0000_0000_0000_0000;
array[52759] <= 16'b0000_0000_0000_0000;
array[52760] <= 16'b0000_0000_0000_0000;
array[52761] <= 16'b0000_0000_0000_0000;
array[52762] <= 16'b0000_0000_0000_0000;
array[52763] <= 16'b0000_0000_0000_0000;
array[52764] <= 16'b0000_0000_0000_0000;
array[52765] <= 16'b0000_0000_0000_0000;
array[52766] <= 16'b0000_0000_0000_0000;
array[52767] <= 16'b0000_0000_0000_0000;
array[52768] <= 16'b0000_0000_0000_0000;
array[52769] <= 16'b0000_0000_0000_0000;
array[52770] <= 16'b0000_0000_0000_0000;
array[52771] <= 16'b0000_0000_0000_0000;
array[52772] <= 16'b0000_0000_0000_0000;
array[52773] <= 16'b0000_0000_0000_0000;
array[52774] <= 16'b0000_0000_0000_0000;
array[52775] <= 16'b0000_0000_0000_0000;
array[52776] <= 16'b0000_0000_0000_0000;
array[52777] <= 16'b0000_0000_0000_0000;
array[52778] <= 16'b0000_0000_0000_0000;
array[52779] <= 16'b0000_0000_0000_0000;
array[52780] <= 16'b0000_0000_0000_0000;
array[52781] <= 16'b0000_0000_0000_0000;
array[52782] <= 16'b0000_0000_0000_0000;
array[52783] <= 16'b0000_0000_0000_0000;
array[52784] <= 16'b0000_0000_0000_0000;
array[52785] <= 16'b0000_0000_0000_0000;
array[52786] <= 16'b0000_0000_0000_0000;
array[52787] <= 16'b0000_0000_0000_0000;
array[52788] <= 16'b0000_0000_0000_0000;
array[52789] <= 16'b0000_0000_0000_0000;
array[52790] <= 16'b0000_0000_0000_0000;
array[52791] <= 16'b0000_0000_0000_0000;
array[52792] <= 16'b0000_0000_0000_0000;
array[52793] <= 16'b0000_0000_0000_0000;
array[52794] <= 16'b0000_0000_0000_0000;
array[52795] <= 16'b0000_0000_0000_0000;
array[52796] <= 16'b0000_0000_0000_0000;
array[52797] <= 16'b0000_0000_0000_0000;
array[52798] <= 16'b0000_0000_0000_0000;
array[52799] <= 16'b0000_0000_0000_0000;
array[52800] <= 16'b0000_0000_0000_0000;
array[52801] <= 16'b0000_0000_0000_0000;
array[52802] <= 16'b0000_0000_0000_0000;
array[52803] <= 16'b0000_0000_0000_0000;
array[52804] <= 16'b0000_0000_0000_0000;
array[52805] <= 16'b0000_0000_0000_0000;
array[52806] <= 16'b0000_0000_0000_0000;
array[52807] <= 16'b0000_0000_0000_0000;
array[52808] <= 16'b0000_0000_0000_0000;
array[52809] <= 16'b0000_0000_0000_0000;
array[52810] <= 16'b0000_0000_0000_0000;
array[52811] <= 16'b0000_0000_0000_0000;
array[52812] <= 16'b0000_0000_0000_0000;
array[52813] <= 16'b0000_0000_0000_0000;
array[52814] <= 16'b0000_0000_0000_0000;
array[52815] <= 16'b0000_0000_0000_0000;
array[52816] <= 16'b0000_0000_0000_0000;
array[52817] <= 16'b0000_0000_0000_0000;
array[52818] <= 16'b0000_0000_0000_0000;
array[52819] <= 16'b0000_0000_0000_0000;
array[52820] <= 16'b0000_0000_0000_0000;
array[52821] <= 16'b0000_0000_0000_0000;
array[52822] <= 16'b0000_0000_0000_0000;
array[52823] <= 16'b0000_0000_0000_0000;
array[52824] <= 16'b0000_0000_0000_0000;
array[52825] <= 16'b0000_0000_0000_0000;
array[52826] <= 16'b0000_0000_0000_0000;
array[52827] <= 16'b0000_0000_0000_0000;
array[52828] <= 16'b0000_0000_0000_0000;
array[52829] <= 16'b0000_0000_0000_0000;
array[52830] <= 16'b0000_0000_0000_0000;
array[52831] <= 16'b0000_0000_0000_0000;
array[52832] <= 16'b0000_0000_0000_0000;
array[52833] <= 16'b0000_0000_0000_0000;
array[52834] <= 16'b0000_0000_0000_0000;
array[52835] <= 16'b0000_0000_0000_0000;
array[52836] <= 16'b0000_0000_0000_0000;
array[52837] <= 16'b0000_0000_0000_0000;
array[52838] <= 16'b0000_0000_0000_0000;
array[52839] <= 16'b0000_0000_0000_0000;
array[52840] <= 16'b0000_0000_0000_0000;
array[52841] <= 16'b0000_0000_0000_0000;
array[52842] <= 16'b0000_0000_0000_0000;
array[52843] <= 16'b0000_0000_0000_0000;
array[52844] <= 16'b0000_0000_0000_0000;
array[52845] <= 16'b0000_0000_0000_0000;
array[52846] <= 16'b0000_0000_0000_0000;
array[52847] <= 16'b0000_0000_0000_0000;
array[52848] <= 16'b0000_0000_0000_0000;
array[52849] <= 16'b0000_0000_0000_0000;
array[52850] <= 16'b0000_0000_0000_0000;
array[52851] <= 16'b0000_0000_0000_0000;
array[52852] <= 16'b0000_0000_0000_0000;
array[52853] <= 16'b0000_0000_0000_0000;
array[52854] <= 16'b0000_0000_0000_0000;
array[52855] <= 16'b0000_0000_0000_0000;
array[52856] <= 16'b0000_0000_0000_0000;
array[52857] <= 16'b0000_0000_0000_0000;
array[52858] <= 16'b0000_0000_0000_0000;
array[52859] <= 16'b0000_0000_0000_0000;
array[52860] <= 16'b0000_0000_0000_0000;
array[52861] <= 16'b0000_0000_0000_0000;
array[52862] <= 16'b0000_0000_0000_0000;
array[52863] <= 16'b0000_0000_0000_0000;
array[52864] <= 16'b0000_0000_0000_0000;
array[52865] <= 16'b0000_0000_0000_0000;
array[52866] <= 16'b0000_0000_0000_0000;
array[52867] <= 16'b0000_0000_0000_0000;
array[52868] <= 16'b0000_0000_0000_0000;
array[52869] <= 16'b0000_0000_0000_0000;
array[52870] <= 16'b0000_0000_0000_0000;
array[52871] <= 16'b0000_0000_0000_0000;
array[52872] <= 16'b0000_0000_0000_0000;
array[52873] <= 16'b0000_0000_0000_0000;
array[52874] <= 16'b0000_0000_0000_0000;
array[52875] <= 16'b0000_0000_0000_0000;
array[52876] <= 16'b0000_0000_0000_0000;
array[52877] <= 16'b0000_0000_0000_0000;
array[52878] <= 16'b0000_0000_0000_0000;
array[52879] <= 16'b0000_0000_0000_0000;
array[52880] <= 16'b0000_0000_0000_0000;
array[52881] <= 16'b0000_0000_0000_0000;
array[52882] <= 16'b0000_0000_0000_0000;
array[52883] <= 16'b0000_0000_0000_0000;
array[52884] <= 16'b0000_0000_0000_0000;
array[52885] <= 16'b0000_0000_0000_0000;
array[52886] <= 16'b0000_0000_0000_0000;
array[52887] <= 16'b0000_0000_0000_0000;
array[52888] <= 16'b0000_0000_0000_0000;
array[52889] <= 16'b0000_0000_0000_0000;
array[52890] <= 16'b0000_0000_0000_0000;
array[52891] <= 16'b0000_0000_0000_0000;
array[52892] <= 16'b0000_0000_0000_0000;
array[52893] <= 16'b0000_0000_0000_0000;
array[52894] <= 16'b0000_0000_0000_0000;
array[52895] <= 16'b0000_0000_0000_0000;
array[52896] <= 16'b0000_0000_0000_0000;
array[52897] <= 16'b0000_0000_0000_0000;
array[52898] <= 16'b0000_0000_0000_0000;
array[52899] <= 16'b0000_0000_0000_0000;
array[52900] <= 16'b0000_0000_0000_0000;
array[52901] <= 16'b0000_0000_0000_0000;
array[52902] <= 16'b0000_0000_0000_0000;
array[52903] <= 16'b0000_0000_0000_0000;
array[52904] <= 16'b0000_0000_0000_0000;
array[52905] <= 16'b0000_0000_0000_0000;
array[52906] <= 16'b0000_0000_0000_0000;
array[52907] <= 16'b0000_0000_0000_0000;
array[52908] <= 16'b0000_0000_0000_0000;
array[52909] <= 16'b0000_0000_0000_0000;
array[52910] <= 16'b0000_0000_0000_0000;
array[52911] <= 16'b0000_0000_0000_0000;
array[52912] <= 16'b0000_0000_0000_0000;
array[52913] <= 16'b0000_0000_0000_0000;
array[52914] <= 16'b0000_0000_0000_0000;
array[52915] <= 16'b0000_0000_0000_0000;
array[52916] <= 16'b0000_0000_0000_0000;
array[52917] <= 16'b0000_0000_0000_0000;
array[52918] <= 16'b0000_0000_0000_0000;
array[52919] <= 16'b0000_0000_0000_0000;
array[52920] <= 16'b0000_0000_0000_0000;
array[52921] <= 16'b0000_0000_0000_0000;
array[52922] <= 16'b0000_0000_0000_0000;
array[52923] <= 16'b0000_0000_0000_0000;
array[52924] <= 16'b0000_0000_0000_0000;
array[52925] <= 16'b0000_0000_0000_0000;
array[52926] <= 16'b0000_0000_0000_0000;
array[52927] <= 16'b0000_0000_0000_0000;
array[52928] <= 16'b0000_0000_0000_0000;
array[52929] <= 16'b0000_0000_0000_0000;
array[52930] <= 16'b0000_0000_0000_0000;
array[52931] <= 16'b0000_0000_0000_0000;
array[52932] <= 16'b0000_0000_0000_0000;
array[52933] <= 16'b0000_0000_0000_0000;
array[52934] <= 16'b0000_0000_0000_0000;
array[52935] <= 16'b0000_0000_0000_0000;
array[52936] <= 16'b0000_0000_0000_0000;
array[52937] <= 16'b0000_0000_0000_0000;
array[52938] <= 16'b0000_0000_0000_0000;
array[52939] <= 16'b0000_0000_0000_0000;
array[52940] <= 16'b0000_0000_0000_0000;
array[52941] <= 16'b0000_0000_0000_0000;
array[52942] <= 16'b0000_0000_0000_0000;
array[52943] <= 16'b0000_0000_0000_0000;
array[52944] <= 16'b0000_0000_0000_0000;
array[52945] <= 16'b0000_0000_0000_0000;
array[52946] <= 16'b0000_0000_0000_0000;
array[52947] <= 16'b0000_0000_0000_0000;
array[52948] <= 16'b0000_0000_0000_0000;
array[52949] <= 16'b0000_0000_0000_0000;
array[52950] <= 16'b0000_0000_0000_0000;
array[52951] <= 16'b0000_0000_0000_0000;
array[52952] <= 16'b0000_0000_0000_0000;
array[52953] <= 16'b0000_0000_0000_0000;
array[52954] <= 16'b0000_0000_0000_0000;
array[52955] <= 16'b0000_0000_0000_0000;
array[52956] <= 16'b0000_0000_0000_0000;
array[52957] <= 16'b0000_0000_0000_0000;
array[52958] <= 16'b0000_0000_0000_0000;
array[52959] <= 16'b0000_0000_0000_0000;
array[52960] <= 16'b0000_0000_0000_0000;
array[52961] <= 16'b0000_0000_0000_0000;
array[52962] <= 16'b0000_0000_0000_0000;
array[52963] <= 16'b0000_0000_0000_0000;
array[52964] <= 16'b0000_0000_0000_0000;
array[52965] <= 16'b0000_0000_0000_0000;
array[52966] <= 16'b0000_0000_0000_0000;
array[52967] <= 16'b0000_0000_0000_0000;
array[52968] <= 16'b0000_0000_0000_0000;
array[52969] <= 16'b0000_0000_0000_0000;
array[52970] <= 16'b0000_0000_0000_0000;
array[52971] <= 16'b0000_0000_0000_0000;
array[52972] <= 16'b0000_0000_0000_0000;
array[52973] <= 16'b0000_0000_0000_0000;
array[52974] <= 16'b0000_0000_0000_0000;
array[52975] <= 16'b0000_0000_0000_0000;
array[52976] <= 16'b0000_0000_0000_0000;
array[52977] <= 16'b0000_0000_0000_0000;
array[52978] <= 16'b0000_0000_0000_0000;
array[52979] <= 16'b0000_0000_0000_0000;
array[52980] <= 16'b0000_0000_0000_0000;
array[52981] <= 16'b0000_0000_0000_0000;
array[52982] <= 16'b0000_0000_0000_0000;
array[52983] <= 16'b0000_0000_0000_0000;
array[52984] <= 16'b0000_0000_0000_0000;
array[52985] <= 16'b0000_0000_0000_0000;
array[52986] <= 16'b0000_0000_0000_0000;
array[52987] <= 16'b0000_0000_0000_0000;
array[52988] <= 16'b0000_0000_0000_0000;
array[52989] <= 16'b0000_0000_0000_0000;
array[52990] <= 16'b0000_0000_0000_0000;
array[52991] <= 16'b0000_0000_0000_0000;
array[52992] <= 16'b0000_0000_0000_0000;
array[52993] <= 16'b0000_0000_0000_0000;
array[52994] <= 16'b0000_0000_0000_0000;
array[52995] <= 16'b0000_0000_0000_0000;
array[52996] <= 16'b0000_0000_0000_0000;
array[52997] <= 16'b0000_0000_0000_0000;
array[52998] <= 16'b0000_0000_0000_0000;
array[52999] <= 16'b0000_0000_0000_0000;
array[53000] <= 16'b0000_0000_0000_0000;
array[53001] <= 16'b0000_0000_0000_0000;
array[53002] <= 16'b0000_0000_0000_0000;
array[53003] <= 16'b0000_0000_0000_0000;
array[53004] <= 16'b0000_0000_0000_0000;
array[53005] <= 16'b0000_0000_0000_0000;
array[53006] <= 16'b0000_0000_0000_0000;
array[53007] <= 16'b0000_0000_0000_0000;
array[53008] <= 16'b0000_0000_0000_0000;
array[53009] <= 16'b0000_0000_0000_0000;
array[53010] <= 16'b0000_0000_0000_0000;
array[53011] <= 16'b0000_0000_0000_0000;
array[53012] <= 16'b0000_0000_0000_0000;
array[53013] <= 16'b0000_0000_0000_0000;
array[53014] <= 16'b0000_0000_0000_0000;
array[53015] <= 16'b0000_0000_0000_0000;
array[53016] <= 16'b0000_0000_0000_0000;
array[53017] <= 16'b0000_0000_0000_0000;
array[53018] <= 16'b0000_0000_0000_0000;
array[53019] <= 16'b0000_0000_0000_0000;
array[53020] <= 16'b0000_0000_0000_0000;
array[53021] <= 16'b0000_0000_0000_0000;
array[53022] <= 16'b0000_0000_0000_0000;
array[53023] <= 16'b0000_0000_0000_0000;
array[53024] <= 16'b0000_0000_0000_0000;
array[53025] <= 16'b0000_0000_0000_0000;
array[53026] <= 16'b0000_0000_0000_0000;
array[53027] <= 16'b0000_0000_0000_0000;
array[53028] <= 16'b0000_0000_0000_0000;
array[53029] <= 16'b0000_0000_0000_0000;
array[53030] <= 16'b0000_0000_0000_0000;
array[53031] <= 16'b0000_0000_0000_0000;
array[53032] <= 16'b0000_0000_0000_0000;
array[53033] <= 16'b0000_0000_0000_0000;
array[53034] <= 16'b0000_0000_0000_0000;
array[53035] <= 16'b0000_0000_0000_0000;
array[53036] <= 16'b0000_0000_0000_0000;
array[53037] <= 16'b0000_0000_0000_0000;
array[53038] <= 16'b0000_0000_0000_0000;
array[53039] <= 16'b0000_0000_0000_0000;
array[53040] <= 16'b0000_0000_0000_0000;
array[53041] <= 16'b0000_0000_0000_0000;
array[53042] <= 16'b0000_0000_0000_0000;
array[53043] <= 16'b0000_0000_0000_0000;
array[53044] <= 16'b0000_0000_0000_0000;
array[53045] <= 16'b0000_0000_0000_0000;
array[53046] <= 16'b0000_0000_0000_0000;
array[53047] <= 16'b0000_0000_0000_0000;
array[53048] <= 16'b0000_0000_0000_0000;
array[53049] <= 16'b0000_0000_0000_0000;
array[53050] <= 16'b0000_0000_0000_0000;
array[53051] <= 16'b0000_0000_0000_0000;
array[53052] <= 16'b0000_0000_0000_0000;
array[53053] <= 16'b0000_0000_0000_0000;
array[53054] <= 16'b0000_0000_0000_0000;
array[53055] <= 16'b0000_0000_0000_0000;
array[53056] <= 16'b0000_0000_0000_0000;
array[53057] <= 16'b0000_0000_0000_0000;
array[53058] <= 16'b0000_0000_0000_0000;
array[53059] <= 16'b0000_0000_0000_0000;
array[53060] <= 16'b0000_0000_0000_0000;
array[53061] <= 16'b0000_0000_0000_0000;
array[53062] <= 16'b0000_0000_0000_0000;
array[53063] <= 16'b0000_0000_0000_0000;
array[53064] <= 16'b0000_0000_0000_0000;
array[53065] <= 16'b0000_0000_0000_0000;
array[53066] <= 16'b0000_0000_0000_0000;
array[53067] <= 16'b0000_0000_0000_0000;
array[53068] <= 16'b0000_0000_0000_0000;
array[53069] <= 16'b0000_0000_0000_0000;
array[53070] <= 16'b0000_0000_0000_0000;
array[53071] <= 16'b0000_0000_0000_0000;
array[53072] <= 16'b0000_0000_0000_0000;
array[53073] <= 16'b0000_0000_0000_0000;
array[53074] <= 16'b0000_0000_0000_0000;
array[53075] <= 16'b0000_0000_0000_0000;
array[53076] <= 16'b0000_0000_0000_0000;
array[53077] <= 16'b0000_0000_0000_0000;
array[53078] <= 16'b0000_0000_0000_0000;
array[53079] <= 16'b0000_0000_0000_0000;
array[53080] <= 16'b0000_0000_0000_0000;
array[53081] <= 16'b0000_0000_0000_0000;
array[53082] <= 16'b0000_0000_0000_0000;
array[53083] <= 16'b0000_0000_0000_0000;
array[53084] <= 16'b0000_0000_0000_0000;
array[53085] <= 16'b0000_0000_0000_0000;
array[53086] <= 16'b0000_0000_0000_0000;
array[53087] <= 16'b0000_0000_0000_0000;
array[53088] <= 16'b0000_0000_0000_0000;
array[53089] <= 16'b0000_0000_0000_0000;
array[53090] <= 16'b0000_0000_0000_0000;
array[53091] <= 16'b0000_0000_0000_0000;
array[53092] <= 16'b0000_0000_0000_0000;
array[53093] <= 16'b0000_0000_0000_0000;
array[53094] <= 16'b0000_0000_0000_0000;
array[53095] <= 16'b0000_0000_0000_0000;
array[53096] <= 16'b0000_0000_0000_0000;
array[53097] <= 16'b0000_0000_0000_0000;
array[53098] <= 16'b0000_0000_0000_0000;
array[53099] <= 16'b0000_0000_0000_0000;
array[53100] <= 16'b0000_0000_0000_0000;
array[53101] <= 16'b0000_0000_0000_0000;
array[53102] <= 16'b0000_0000_0000_0000;
array[53103] <= 16'b0000_0000_0000_0000;
array[53104] <= 16'b0000_0000_0000_0000;
array[53105] <= 16'b0000_0000_0000_0000;
array[53106] <= 16'b0000_0000_0000_0000;
array[53107] <= 16'b0000_0000_0000_0000;
array[53108] <= 16'b0000_0000_0000_0000;
array[53109] <= 16'b0000_0000_0000_0000;
array[53110] <= 16'b0000_0000_0000_0000;
array[53111] <= 16'b0000_0000_0000_0000;
array[53112] <= 16'b0000_0000_0000_0000;
array[53113] <= 16'b0000_0000_0000_0000;
array[53114] <= 16'b0000_0000_0000_0000;
array[53115] <= 16'b0000_0000_0000_0000;
array[53116] <= 16'b0000_0000_0000_0000;
array[53117] <= 16'b0000_0000_0000_0000;
array[53118] <= 16'b0000_0000_0000_0000;
array[53119] <= 16'b0000_0000_0000_0000;
array[53120] <= 16'b0000_0000_0000_0000;
array[53121] <= 16'b0000_0000_0000_0000;
array[53122] <= 16'b0000_0000_0000_0000;
array[53123] <= 16'b0000_0000_0000_0000;
array[53124] <= 16'b0000_0000_0000_0000;
array[53125] <= 16'b0000_0000_0000_0000;
array[53126] <= 16'b0000_0000_0000_0000;
array[53127] <= 16'b0000_0000_0000_0000;
array[53128] <= 16'b0000_0000_0000_0000;
array[53129] <= 16'b0000_0000_0000_0000;
array[53130] <= 16'b0000_0000_0000_0000;
array[53131] <= 16'b0000_0000_0000_0000;
array[53132] <= 16'b0000_0000_0000_0000;
array[53133] <= 16'b0000_0000_0000_0000;
array[53134] <= 16'b0000_0000_0000_0000;
array[53135] <= 16'b0000_0000_0000_0000;
array[53136] <= 16'b0000_0000_0000_0000;
array[53137] <= 16'b0000_0000_0000_0000;
array[53138] <= 16'b0000_0000_0000_0000;
array[53139] <= 16'b0000_0000_0000_0000;
array[53140] <= 16'b0000_0000_0000_0000;
array[53141] <= 16'b0000_0000_0000_0000;
array[53142] <= 16'b0000_0000_0000_0000;
array[53143] <= 16'b0000_0000_0000_0000;
array[53144] <= 16'b0000_0000_0000_0000;
array[53145] <= 16'b0000_0000_0000_0000;
array[53146] <= 16'b0000_0000_0000_0000;
array[53147] <= 16'b0000_0000_0000_0000;
array[53148] <= 16'b0000_0000_0000_0000;
array[53149] <= 16'b0000_0000_0000_0000;
array[53150] <= 16'b0000_0000_0000_0000;
array[53151] <= 16'b0000_0000_0000_0000;
array[53152] <= 16'b0000_0000_0000_0000;
array[53153] <= 16'b0000_0000_0000_0000;
array[53154] <= 16'b0000_0000_0000_0000;
array[53155] <= 16'b0000_0000_0000_0000;
array[53156] <= 16'b0000_0000_0000_0000;
array[53157] <= 16'b0000_0000_0000_0000;
array[53158] <= 16'b0000_0000_0000_0000;
array[53159] <= 16'b0000_0000_0000_0000;
array[53160] <= 16'b0000_0000_0000_0000;
array[53161] <= 16'b0000_0000_0000_0000;
array[53162] <= 16'b0000_0000_0000_0000;
array[53163] <= 16'b0000_0000_0000_0000;
array[53164] <= 16'b0000_0000_0000_0000;
array[53165] <= 16'b0000_0000_0000_0000;
array[53166] <= 16'b0000_0000_0000_0000;
array[53167] <= 16'b0000_0000_0000_0000;
array[53168] <= 16'b0000_0000_0000_0000;
array[53169] <= 16'b0000_0000_0000_0000;
array[53170] <= 16'b0000_0000_0000_0000;
array[53171] <= 16'b0000_0000_0000_0000;
array[53172] <= 16'b0000_0000_0000_0000;
array[53173] <= 16'b0000_0000_0000_0000;
array[53174] <= 16'b0000_0000_0000_0000;
array[53175] <= 16'b0000_0000_0000_0000;
array[53176] <= 16'b0000_0000_0000_0000;
array[53177] <= 16'b0000_0000_0000_0000;
array[53178] <= 16'b0000_0000_0000_0000;
array[53179] <= 16'b0000_0000_0000_0000;
array[53180] <= 16'b0000_0000_0000_0000;
array[53181] <= 16'b0000_0000_0000_0000;
array[53182] <= 16'b0000_0000_0000_0000;
array[53183] <= 16'b0000_0000_0000_0000;
array[53184] <= 16'b0000_0000_0000_0000;
array[53185] <= 16'b0000_0000_0000_0000;
array[53186] <= 16'b0000_0000_0000_0000;
array[53187] <= 16'b0000_0000_0000_0000;
array[53188] <= 16'b0000_0000_0000_0000;
array[53189] <= 16'b0000_0000_0000_0000;
array[53190] <= 16'b0000_0000_0000_0000;
array[53191] <= 16'b0000_0000_0000_0000;
array[53192] <= 16'b0000_0000_0000_0000;
array[53193] <= 16'b0000_0000_0000_0000;
array[53194] <= 16'b0000_0000_0000_0000;
array[53195] <= 16'b0000_0000_0000_0000;
array[53196] <= 16'b0000_0000_0000_0000;
array[53197] <= 16'b0000_0000_0000_0000;
array[53198] <= 16'b0000_0000_0000_0000;
array[53199] <= 16'b0000_0000_0000_0000;
array[53200] <= 16'b0000_0000_0000_0000;
array[53201] <= 16'b0000_0000_0000_0000;
array[53202] <= 16'b0000_0000_0000_0000;
array[53203] <= 16'b0000_0000_0000_0000;
array[53204] <= 16'b0000_0000_0000_0000;
array[53205] <= 16'b0000_0000_0000_0000;
array[53206] <= 16'b0000_0000_0000_0000;
array[53207] <= 16'b0000_0000_0000_0000;
array[53208] <= 16'b0000_0000_0000_0000;
array[53209] <= 16'b0000_0000_0000_0000;
array[53210] <= 16'b0000_0000_0000_0000;
array[53211] <= 16'b0000_0000_0000_0000;
array[53212] <= 16'b0000_0000_0000_0000;
array[53213] <= 16'b0000_0000_0000_0000;
array[53214] <= 16'b0000_0000_0000_0000;
array[53215] <= 16'b0000_0000_0000_0000;
array[53216] <= 16'b0000_0000_0000_0000;
array[53217] <= 16'b0000_0000_0000_0000;
array[53218] <= 16'b0000_0000_0000_0000;
array[53219] <= 16'b0000_0000_0000_0000;
array[53220] <= 16'b0000_0000_0000_0000;
array[53221] <= 16'b0000_0000_0000_0000;
array[53222] <= 16'b0000_0000_0000_0000;
array[53223] <= 16'b0000_0000_0000_0000;
array[53224] <= 16'b0000_0000_0000_0000;
array[53225] <= 16'b0000_0000_0000_0000;
array[53226] <= 16'b0000_0000_0000_0000;
array[53227] <= 16'b0000_0000_0000_0000;
array[53228] <= 16'b0000_0000_0000_0000;
array[53229] <= 16'b0000_0000_0000_0000;
array[53230] <= 16'b0000_0000_0000_0000;
array[53231] <= 16'b0000_0000_0000_0000;
array[53232] <= 16'b0000_0000_0000_0000;
array[53233] <= 16'b0000_0000_0000_0000;
array[53234] <= 16'b0000_0000_0000_0000;
array[53235] <= 16'b0000_0000_0000_0000;
array[53236] <= 16'b0000_0000_0000_0000;
array[53237] <= 16'b0000_0000_0000_0000;
array[53238] <= 16'b0000_0000_0000_0000;
array[53239] <= 16'b0000_0000_0000_0000;
array[53240] <= 16'b0000_0000_0000_0000;
array[53241] <= 16'b0000_0000_0000_0000;
array[53242] <= 16'b0000_0000_0000_0000;
array[53243] <= 16'b0000_0000_0000_0000;
array[53244] <= 16'b0000_0000_0000_0000;
array[53245] <= 16'b0000_0000_0000_0000;
array[53246] <= 16'b0000_0000_0000_0000;
array[53247] <= 16'b0000_0000_0000_0000;
array[53248] <= 16'b0000_0000_0000_0000;
array[53249] <= 16'b0000_0000_0000_0000;
array[53250] <= 16'b0000_0000_0000_0000;
array[53251] <= 16'b0000_0000_0000_0000;
array[53252] <= 16'b0000_0000_0000_0000;
array[53253] <= 16'b0000_0000_0000_0000;
array[53254] <= 16'b0000_0000_0000_0000;
array[53255] <= 16'b0000_0000_0000_0000;
array[53256] <= 16'b0000_0000_0000_0000;
array[53257] <= 16'b0000_0000_0000_0000;
array[53258] <= 16'b0000_0000_0000_0000;
array[53259] <= 16'b0000_0000_0000_0000;
array[53260] <= 16'b0000_0000_0000_0000;
array[53261] <= 16'b0000_0000_0000_0000;
array[53262] <= 16'b0000_0000_0000_0000;
array[53263] <= 16'b0000_0000_0000_0000;
array[53264] <= 16'b0000_0000_0000_0000;
array[53265] <= 16'b0000_0000_0000_0000;
array[53266] <= 16'b0000_0000_0000_0000;
array[53267] <= 16'b0000_0000_0000_0000;
array[53268] <= 16'b0000_0000_0000_0000;
array[53269] <= 16'b0000_0000_0000_0000;
array[53270] <= 16'b0000_0000_0000_0000;
array[53271] <= 16'b0000_0000_0000_0000;
array[53272] <= 16'b0000_0000_0000_0000;
array[53273] <= 16'b0000_0000_0000_0000;
array[53274] <= 16'b0000_0000_0000_0000;
array[53275] <= 16'b0000_0000_0000_0000;
array[53276] <= 16'b0000_0000_0000_0000;
array[53277] <= 16'b0000_0000_0000_0000;
array[53278] <= 16'b0000_0000_0000_0000;
array[53279] <= 16'b0000_0000_0000_0000;
array[53280] <= 16'b0000_0000_0000_0000;
array[53281] <= 16'b0000_0000_0000_0000;
array[53282] <= 16'b0000_0000_0000_0000;
array[53283] <= 16'b0000_0000_0000_0000;
array[53284] <= 16'b0000_0000_0000_0000;
array[53285] <= 16'b0000_0000_0000_0000;
array[53286] <= 16'b0000_0000_0000_0000;
array[53287] <= 16'b0000_0000_0000_0000;
array[53288] <= 16'b0000_0000_0000_0000;
array[53289] <= 16'b0000_0000_0000_0000;
array[53290] <= 16'b0000_0000_0000_0000;
array[53291] <= 16'b0000_0000_0000_0000;
array[53292] <= 16'b0000_0000_0000_0000;
array[53293] <= 16'b0000_0000_0000_0000;
array[53294] <= 16'b0000_0000_0000_0000;
array[53295] <= 16'b0000_0000_0000_0000;
array[53296] <= 16'b0000_0000_0000_0000;
array[53297] <= 16'b0000_0000_0000_0000;
array[53298] <= 16'b0000_0000_0000_0000;
array[53299] <= 16'b0000_0000_0000_0000;
array[53300] <= 16'b0000_0000_0000_0000;
array[53301] <= 16'b0000_0000_0000_0000;
array[53302] <= 16'b0000_0000_0000_0000;
array[53303] <= 16'b0000_0000_0000_0000;
array[53304] <= 16'b0000_0000_0000_0000;
array[53305] <= 16'b0000_0000_0000_0000;
array[53306] <= 16'b0000_0000_0000_0000;
array[53307] <= 16'b0000_0000_0000_0000;
array[53308] <= 16'b0000_0000_0000_0000;
array[53309] <= 16'b0000_0000_0000_0000;
array[53310] <= 16'b0000_0000_0000_0000;
array[53311] <= 16'b0000_0000_0000_0000;
array[53312] <= 16'b0000_0000_0000_0000;
array[53313] <= 16'b0000_0000_0000_0000;
array[53314] <= 16'b0000_0000_0000_0000;
array[53315] <= 16'b0000_0000_0000_0000;
array[53316] <= 16'b0000_0000_0000_0000;
array[53317] <= 16'b0000_0000_0000_0000;
array[53318] <= 16'b0000_0000_0000_0000;
array[53319] <= 16'b0000_0000_0000_0000;
array[53320] <= 16'b0000_0000_0000_0000;
array[53321] <= 16'b0000_0000_0000_0000;
array[53322] <= 16'b0000_0000_0000_0000;
array[53323] <= 16'b0000_0000_0000_0000;
array[53324] <= 16'b0000_0000_0000_0000;
array[53325] <= 16'b0000_0000_0000_0000;
array[53326] <= 16'b0000_0000_0000_0000;
array[53327] <= 16'b0000_0000_0000_0000;
array[53328] <= 16'b0000_0000_0000_0000;
array[53329] <= 16'b0000_0000_0000_0000;
array[53330] <= 16'b0000_0000_0000_0000;
array[53331] <= 16'b0000_0000_0000_0000;
array[53332] <= 16'b0000_0000_0000_0000;
array[53333] <= 16'b0000_0000_0000_0000;
array[53334] <= 16'b0000_0000_0000_0000;
array[53335] <= 16'b0000_0000_0000_0000;
array[53336] <= 16'b0000_0000_0000_0000;
array[53337] <= 16'b0000_0000_0000_0000;
array[53338] <= 16'b0000_0000_0000_0000;
array[53339] <= 16'b0000_0000_0000_0000;
array[53340] <= 16'b0000_0000_0000_0000;
array[53341] <= 16'b0000_0000_0000_0000;
array[53342] <= 16'b0000_0000_0000_0000;
array[53343] <= 16'b0000_0000_0000_0000;
array[53344] <= 16'b0000_0000_0000_0000;
array[53345] <= 16'b0000_0000_0000_0000;
array[53346] <= 16'b0000_0000_0000_0000;
array[53347] <= 16'b0000_0000_0000_0000;
array[53348] <= 16'b0000_0000_0000_0000;
array[53349] <= 16'b0000_0000_0000_0000;
array[53350] <= 16'b0000_0000_0000_0000;
array[53351] <= 16'b0000_0000_0000_0000;
array[53352] <= 16'b0000_0000_0000_0000;
array[53353] <= 16'b0000_0000_0000_0000;
array[53354] <= 16'b0000_0000_0000_0000;
array[53355] <= 16'b0000_0000_0000_0000;
array[53356] <= 16'b0000_0000_0000_0000;
array[53357] <= 16'b0000_0000_0000_0000;
array[53358] <= 16'b0000_0000_0000_0000;
array[53359] <= 16'b0000_0000_0000_0000;
array[53360] <= 16'b0000_0000_0000_0000;
array[53361] <= 16'b0000_0000_0000_0000;
array[53362] <= 16'b0000_0000_0000_0000;
array[53363] <= 16'b0000_0000_0000_0000;
array[53364] <= 16'b0000_0000_0000_0000;
array[53365] <= 16'b0000_0000_0000_0000;
array[53366] <= 16'b0000_0000_0000_0000;
array[53367] <= 16'b0000_0000_0000_0000;
array[53368] <= 16'b0000_0000_0000_0000;
array[53369] <= 16'b0000_0000_0000_0000;
array[53370] <= 16'b0000_0000_0000_0000;
array[53371] <= 16'b0000_0000_0000_0000;
array[53372] <= 16'b0000_0000_0000_0000;
array[53373] <= 16'b0000_0000_0000_0000;
array[53374] <= 16'b0000_0000_0000_0000;
array[53375] <= 16'b0000_0000_0000_0000;
array[53376] <= 16'b0000_0000_0000_0000;
array[53377] <= 16'b0000_0000_0000_0000;
array[53378] <= 16'b0000_0000_0000_0000;
array[53379] <= 16'b0000_0000_0000_0000;
array[53380] <= 16'b0000_0000_0000_0000;
array[53381] <= 16'b0000_0000_0000_0000;
array[53382] <= 16'b0000_0000_0000_0000;
array[53383] <= 16'b0000_0000_0000_0000;
array[53384] <= 16'b0000_0000_0000_0000;
array[53385] <= 16'b0000_0000_0000_0000;
array[53386] <= 16'b0000_0000_0000_0000;
array[53387] <= 16'b0000_0000_0000_0000;
array[53388] <= 16'b0000_0000_0000_0000;
array[53389] <= 16'b0000_0000_0000_0000;
array[53390] <= 16'b0000_0000_0000_0000;
array[53391] <= 16'b0000_0000_0000_0000;
array[53392] <= 16'b0000_0000_0000_0000;
array[53393] <= 16'b0000_0000_0000_0000;
array[53394] <= 16'b0000_0000_0000_0000;
array[53395] <= 16'b0000_0000_0000_0000;
array[53396] <= 16'b0000_0000_0000_0000;
array[53397] <= 16'b0000_0000_0000_0000;
array[53398] <= 16'b0000_0000_0000_0000;
array[53399] <= 16'b0000_0000_0000_0000;
array[53400] <= 16'b0000_0000_0000_0000;
array[53401] <= 16'b0000_0000_0000_0000;
array[53402] <= 16'b0000_0000_0000_0000;
array[53403] <= 16'b0000_0000_0000_0000;
array[53404] <= 16'b0000_0000_0000_0000;
array[53405] <= 16'b0000_0000_0000_0000;
array[53406] <= 16'b0000_0000_0000_0000;
array[53407] <= 16'b0000_0000_0000_0000;
array[53408] <= 16'b0000_0000_0000_0000;
array[53409] <= 16'b0000_0000_0000_0000;
array[53410] <= 16'b0000_0000_0000_0000;
array[53411] <= 16'b0000_0000_0000_0000;
array[53412] <= 16'b0000_0000_0000_0000;
array[53413] <= 16'b0000_0000_0000_0000;
array[53414] <= 16'b0000_0000_0000_0000;
array[53415] <= 16'b0000_0000_0000_0000;
array[53416] <= 16'b0000_0000_0000_0000;
array[53417] <= 16'b0000_0000_0000_0000;
array[53418] <= 16'b0000_0000_0000_0000;
array[53419] <= 16'b0000_0000_0000_0000;
array[53420] <= 16'b0000_0000_0000_0000;
array[53421] <= 16'b0000_0000_0000_0000;
array[53422] <= 16'b0000_0000_0000_0000;
array[53423] <= 16'b0000_0000_0000_0000;
array[53424] <= 16'b0000_0000_0000_0000;
array[53425] <= 16'b0000_0000_0000_0000;
array[53426] <= 16'b0000_0000_0000_0000;
array[53427] <= 16'b0000_0000_0000_0000;
array[53428] <= 16'b0000_0000_0000_0000;
array[53429] <= 16'b0000_0000_0000_0000;
array[53430] <= 16'b0000_0000_0000_0000;
array[53431] <= 16'b0000_0000_0000_0000;
array[53432] <= 16'b0000_0000_0000_0000;
array[53433] <= 16'b0000_0000_0000_0000;
array[53434] <= 16'b0000_0000_0000_0000;
array[53435] <= 16'b0000_0000_0000_0000;
array[53436] <= 16'b0000_0000_0000_0000;
array[53437] <= 16'b0000_0000_0000_0000;
array[53438] <= 16'b0000_0000_0000_0000;
array[53439] <= 16'b0000_0000_0000_0000;
array[53440] <= 16'b0000_0000_0000_0000;
array[53441] <= 16'b0000_0000_0000_0000;
array[53442] <= 16'b0000_0000_0000_0000;
array[53443] <= 16'b0000_0000_0000_0000;
array[53444] <= 16'b0000_0000_0000_0000;
array[53445] <= 16'b0000_0000_0000_0000;
array[53446] <= 16'b0000_0000_0000_0000;
array[53447] <= 16'b0000_0000_0000_0000;
array[53448] <= 16'b0000_0000_0000_0000;
array[53449] <= 16'b0000_0000_0000_0000;
array[53450] <= 16'b0000_0000_0000_0000;
array[53451] <= 16'b0000_0000_0000_0000;
array[53452] <= 16'b0000_0000_0000_0000;
array[53453] <= 16'b0000_0000_0000_0000;
array[53454] <= 16'b0000_0000_0000_0000;
array[53455] <= 16'b0000_0000_0000_0000;
array[53456] <= 16'b0000_0000_0000_0000;
array[53457] <= 16'b0000_0000_0000_0000;
array[53458] <= 16'b0000_0000_0000_0000;
array[53459] <= 16'b0000_0000_0000_0000;
array[53460] <= 16'b0000_0000_0000_0000;
array[53461] <= 16'b0000_0000_0000_0000;
array[53462] <= 16'b0000_0000_0000_0000;
array[53463] <= 16'b0000_0000_0000_0000;
array[53464] <= 16'b0000_0000_0000_0000;
array[53465] <= 16'b0000_0000_0000_0000;
array[53466] <= 16'b0000_0000_0000_0000;
array[53467] <= 16'b0000_0000_0000_0000;
array[53468] <= 16'b0000_0000_0000_0000;
array[53469] <= 16'b0000_0000_0000_0000;
array[53470] <= 16'b0000_0000_0000_0000;
array[53471] <= 16'b0000_0000_0000_0000;
array[53472] <= 16'b0000_0000_0000_0000;
array[53473] <= 16'b0000_0000_0000_0000;
array[53474] <= 16'b0000_0000_0000_0000;
array[53475] <= 16'b0000_0000_0000_0000;
array[53476] <= 16'b0000_0000_0000_0000;
array[53477] <= 16'b0000_0000_0000_0000;
array[53478] <= 16'b0000_0000_0000_0000;
array[53479] <= 16'b0000_0000_0000_0000;
array[53480] <= 16'b0000_0000_0000_0000;
array[53481] <= 16'b0000_0000_0000_0000;
array[53482] <= 16'b0000_0000_0000_0000;
array[53483] <= 16'b0000_0000_0000_0000;
array[53484] <= 16'b0000_0000_0000_0000;
array[53485] <= 16'b0000_0000_0000_0000;
array[53486] <= 16'b0000_0000_0000_0000;
array[53487] <= 16'b0000_0000_0000_0000;
array[53488] <= 16'b0000_0000_0000_0000;
array[53489] <= 16'b0000_0000_0000_0000;
array[53490] <= 16'b0000_0000_0000_0000;
array[53491] <= 16'b0000_0000_0000_0000;
array[53492] <= 16'b0000_0000_0000_0000;
array[53493] <= 16'b0000_0000_0000_0000;
array[53494] <= 16'b0000_0000_0000_0000;
array[53495] <= 16'b0000_0000_0000_0000;
array[53496] <= 16'b0000_0000_0000_0000;
array[53497] <= 16'b0000_0000_0000_0000;
array[53498] <= 16'b0000_0000_0000_0000;
array[53499] <= 16'b0000_0000_0000_0000;
array[53500] <= 16'b0000_0000_0000_0000;
array[53501] <= 16'b0000_0000_0000_0000;
array[53502] <= 16'b0000_0000_0000_0000;
array[53503] <= 16'b0000_0000_0000_0000;
array[53504] <= 16'b0000_0000_0000_0000;
array[53505] <= 16'b0000_0000_0000_0000;
array[53506] <= 16'b0000_0000_0000_0000;
array[53507] <= 16'b0000_0000_0000_0000;
array[53508] <= 16'b0000_0000_0000_0000;
array[53509] <= 16'b0000_0000_0000_0000;
array[53510] <= 16'b0000_0000_0000_0000;
array[53511] <= 16'b0000_0000_0000_0000;
array[53512] <= 16'b0000_0000_0000_0000;
array[53513] <= 16'b0000_0000_0000_0000;
array[53514] <= 16'b0000_0000_0000_0000;
array[53515] <= 16'b0000_0000_0000_0000;
array[53516] <= 16'b0000_0000_0000_0000;
array[53517] <= 16'b0000_0000_0000_0000;
array[53518] <= 16'b0000_0000_0000_0000;
array[53519] <= 16'b0000_0000_0000_0000;
array[53520] <= 16'b0000_0000_0000_0000;
array[53521] <= 16'b0000_0000_0000_0000;
array[53522] <= 16'b0000_0000_0000_0000;
array[53523] <= 16'b0000_0000_0000_0000;
array[53524] <= 16'b0000_0000_0000_0000;
array[53525] <= 16'b0000_0000_0000_0000;
array[53526] <= 16'b0000_0000_0000_0000;
array[53527] <= 16'b0000_0000_0000_0000;
array[53528] <= 16'b0000_0000_0000_0000;
array[53529] <= 16'b0000_0000_0000_0000;
array[53530] <= 16'b0000_0000_0000_0000;
array[53531] <= 16'b0000_0000_0000_0000;
array[53532] <= 16'b0000_0000_0000_0000;
array[53533] <= 16'b0000_0000_0000_0000;
array[53534] <= 16'b0000_0000_0000_0000;
array[53535] <= 16'b0000_0000_0000_0000;
array[53536] <= 16'b0000_0000_0000_0000;
array[53537] <= 16'b0000_0000_0000_0000;
array[53538] <= 16'b0000_0000_0000_0000;
array[53539] <= 16'b0000_0000_0000_0000;
array[53540] <= 16'b0000_0000_0000_0000;
array[53541] <= 16'b0000_0000_0000_0000;
array[53542] <= 16'b0000_0000_0000_0000;
array[53543] <= 16'b0000_0000_0000_0000;
array[53544] <= 16'b0000_0000_0000_0000;
array[53545] <= 16'b0000_0000_0000_0000;
array[53546] <= 16'b0000_0000_0000_0000;
array[53547] <= 16'b0000_0000_0000_0000;
array[53548] <= 16'b0000_0000_0000_0000;
array[53549] <= 16'b0000_0000_0000_0000;
array[53550] <= 16'b0000_0000_0000_0000;
array[53551] <= 16'b0000_0000_0000_0000;
array[53552] <= 16'b0000_0000_0000_0000;
array[53553] <= 16'b0000_0000_0000_0000;
array[53554] <= 16'b0000_0000_0000_0000;
array[53555] <= 16'b0000_0000_0000_0000;
array[53556] <= 16'b0000_0000_0000_0000;
array[53557] <= 16'b0000_0000_0000_0000;
array[53558] <= 16'b0000_0000_0000_0000;
array[53559] <= 16'b0000_0000_0000_0000;
array[53560] <= 16'b0000_0000_0000_0000;
array[53561] <= 16'b0000_0000_0000_0000;
array[53562] <= 16'b0000_0000_0000_0000;
array[53563] <= 16'b0000_0000_0000_0000;
array[53564] <= 16'b0000_0000_0000_0000;
array[53565] <= 16'b0000_0000_0000_0000;
array[53566] <= 16'b0000_0000_0000_0000;
array[53567] <= 16'b0000_0000_0000_0000;
array[53568] <= 16'b0000_0000_0000_0000;
array[53569] <= 16'b0000_0000_0000_0000;
array[53570] <= 16'b0000_0000_0000_0000;
array[53571] <= 16'b0000_0000_0000_0000;
array[53572] <= 16'b0000_0000_0000_0000;
array[53573] <= 16'b0000_0000_0000_0000;
array[53574] <= 16'b0000_0000_0000_0000;
array[53575] <= 16'b0000_0000_0000_0000;
array[53576] <= 16'b0000_0000_0000_0000;
array[53577] <= 16'b0000_0000_0000_0000;
array[53578] <= 16'b0000_0000_0000_0000;
array[53579] <= 16'b0000_0000_0000_0000;
array[53580] <= 16'b0000_0000_0000_0000;
array[53581] <= 16'b0000_0000_0000_0000;
array[53582] <= 16'b0000_0000_0000_0000;
array[53583] <= 16'b0000_0000_0000_0000;
array[53584] <= 16'b0000_0000_0000_0000;
array[53585] <= 16'b0000_0000_0000_0000;
array[53586] <= 16'b0000_0000_0000_0000;
array[53587] <= 16'b0000_0000_0000_0000;
array[53588] <= 16'b0000_0000_0000_0000;
array[53589] <= 16'b0000_0000_0000_0000;
array[53590] <= 16'b0000_0000_0000_0000;
array[53591] <= 16'b0000_0000_0000_0000;
array[53592] <= 16'b0000_0000_0000_0000;
array[53593] <= 16'b0000_0000_0000_0000;
array[53594] <= 16'b0000_0000_0000_0000;
array[53595] <= 16'b0000_0000_0000_0000;
array[53596] <= 16'b0000_0000_0000_0000;
array[53597] <= 16'b0000_0000_0000_0000;
array[53598] <= 16'b0000_0000_0000_0000;
array[53599] <= 16'b0000_0000_0000_0000;
array[53600] <= 16'b0000_0000_0000_0000;
array[53601] <= 16'b0000_0000_0000_0000;
array[53602] <= 16'b0000_0000_0000_0000;
array[53603] <= 16'b0000_0000_0000_0000;
array[53604] <= 16'b0000_0000_0000_0000;
array[53605] <= 16'b0000_0000_0000_0000;
array[53606] <= 16'b0000_0000_0000_0000;
array[53607] <= 16'b0000_0000_0000_0000;
array[53608] <= 16'b0000_0000_0000_0000;
array[53609] <= 16'b0000_0000_0000_0000;
array[53610] <= 16'b0000_0000_0000_0000;
array[53611] <= 16'b0000_0000_0000_0000;
array[53612] <= 16'b0000_0000_0000_0000;
array[53613] <= 16'b0000_0000_0000_0000;
array[53614] <= 16'b0000_0000_0000_0000;
array[53615] <= 16'b0000_0000_0000_0000;
array[53616] <= 16'b0000_0000_0000_0000;
array[53617] <= 16'b0000_0000_0000_0000;
array[53618] <= 16'b0000_0000_0000_0000;
array[53619] <= 16'b0000_0000_0000_0000;
array[53620] <= 16'b0000_0000_0000_0000;
array[53621] <= 16'b0000_0000_0000_0000;
array[53622] <= 16'b0000_0000_0000_0000;
array[53623] <= 16'b0000_0000_0000_0000;
array[53624] <= 16'b0000_0000_0000_0000;
array[53625] <= 16'b0000_0000_0000_0000;
array[53626] <= 16'b0000_0000_0000_0000;
array[53627] <= 16'b0000_0000_0000_0000;
array[53628] <= 16'b0000_0000_0000_0000;
array[53629] <= 16'b0000_0000_0000_0000;
array[53630] <= 16'b0000_0000_0000_0000;
array[53631] <= 16'b0000_0000_0000_0000;
array[53632] <= 16'b0000_0000_0000_0000;
array[53633] <= 16'b0000_0000_0000_0000;
array[53634] <= 16'b0000_0000_0000_0000;
array[53635] <= 16'b0000_0000_0000_0000;
array[53636] <= 16'b0000_0000_0000_0000;
array[53637] <= 16'b0000_0000_0000_0000;
array[53638] <= 16'b0000_0000_0000_0000;
array[53639] <= 16'b0000_0000_0000_0000;
array[53640] <= 16'b0000_0000_0000_0000;
array[53641] <= 16'b0000_0000_0000_0000;
array[53642] <= 16'b0000_0000_0000_0000;
array[53643] <= 16'b0000_0000_0000_0000;
array[53644] <= 16'b0000_0000_0000_0000;
array[53645] <= 16'b0000_0000_0000_0000;
array[53646] <= 16'b0000_0000_0000_0000;
array[53647] <= 16'b0000_0000_0000_0000;
array[53648] <= 16'b0000_0000_0000_0000;
array[53649] <= 16'b0000_0000_0000_0000;
array[53650] <= 16'b0000_0000_0000_0000;
array[53651] <= 16'b0000_0000_0000_0000;
array[53652] <= 16'b0000_0000_0000_0000;
array[53653] <= 16'b0000_0000_0000_0000;
array[53654] <= 16'b0000_0000_0000_0000;
array[53655] <= 16'b0000_0000_0000_0000;
array[53656] <= 16'b0000_0000_0000_0000;
array[53657] <= 16'b0000_0000_0000_0000;
array[53658] <= 16'b0000_0000_0000_0000;
array[53659] <= 16'b0000_0000_0000_0000;
array[53660] <= 16'b0000_0000_0000_0000;
array[53661] <= 16'b0000_0000_0000_0000;
array[53662] <= 16'b0000_0000_0000_0000;
array[53663] <= 16'b0000_0000_0000_0000;
array[53664] <= 16'b0000_0000_0000_0000;
array[53665] <= 16'b0000_0000_0000_0000;
array[53666] <= 16'b0000_0000_0000_0000;
array[53667] <= 16'b0000_0000_0000_0000;
array[53668] <= 16'b0000_0000_0000_0000;
array[53669] <= 16'b0000_0000_0000_0000;
array[53670] <= 16'b0000_0000_0000_0000;
array[53671] <= 16'b0000_0000_0000_0000;
array[53672] <= 16'b0000_0000_0000_0000;
array[53673] <= 16'b0000_0000_0000_0000;
array[53674] <= 16'b0000_0000_0000_0000;
array[53675] <= 16'b0000_0000_0000_0000;
array[53676] <= 16'b0000_0000_0000_0000;
array[53677] <= 16'b0000_0000_0000_0000;
array[53678] <= 16'b0000_0000_0000_0000;
array[53679] <= 16'b0000_0000_0000_0000;
array[53680] <= 16'b0000_0000_0000_0000;
array[53681] <= 16'b0000_0000_0000_0000;
array[53682] <= 16'b0000_0000_0000_0000;
array[53683] <= 16'b0000_0000_0000_0000;
array[53684] <= 16'b0000_0000_0000_0000;
array[53685] <= 16'b0000_0000_0000_0000;
array[53686] <= 16'b0000_0000_0000_0000;
array[53687] <= 16'b0000_0000_0000_0000;
array[53688] <= 16'b0000_0000_0000_0000;
array[53689] <= 16'b0000_0000_0000_0000;
array[53690] <= 16'b0000_0000_0000_0000;
array[53691] <= 16'b0000_0000_0000_0000;
array[53692] <= 16'b0000_0000_0000_0000;
array[53693] <= 16'b0000_0000_0000_0000;
array[53694] <= 16'b0000_0000_0000_0000;
array[53695] <= 16'b0000_0000_0000_0000;
array[53696] <= 16'b0000_0000_0000_0000;
array[53697] <= 16'b0000_0000_0000_0000;
array[53698] <= 16'b0000_0000_0000_0000;
array[53699] <= 16'b0000_0000_0000_0000;
array[53700] <= 16'b0000_0000_0000_0000;
array[53701] <= 16'b0000_0000_0000_0000;
array[53702] <= 16'b0000_0000_0000_0000;
array[53703] <= 16'b0000_0000_0000_0000;
array[53704] <= 16'b0000_0000_0000_0000;
array[53705] <= 16'b0000_0000_0000_0000;
array[53706] <= 16'b0000_0000_0000_0000;
array[53707] <= 16'b0000_0000_0000_0000;
array[53708] <= 16'b0000_0000_0000_0000;
array[53709] <= 16'b0000_0000_0000_0000;
array[53710] <= 16'b0000_0000_0000_0000;
array[53711] <= 16'b0000_0000_0000_0000;
array[53712] <= 16'b0000_0000_0000_0000;
array[53713] <= 16'b0000_0000_0000_0000;
array[53714] <= 16'b0000_0000_0000_0000;
array[53715] <= 16'b0000_0000_0000_0000;
array[53716] <= 16'b0000_0000_0000_0000;
array[53717] <= 16'b0000_0000_0000_0000;
array[53718] <= 16'b0000_0000_0000_0000;
array[53719] <= 16'b0000_0000_0000_0000;
array[53720] <= 16'b0000_0000_0000_0000;
array[53721] <= 16'b0000_0000_0000_0000;
array[53722] <= 16'b0000_0000_0000_0000;
array[53723] <= 16'b0000_0000_0000_0000;
array[53724] <= 16'b0000_0000_0000_0000;
array[53725] <= 16'b0000_0000_0000_0000;
array[53726] <= 16'b0000_0000_0000_0000;
array[53727] <= 16'b0000_0000_0000_0000;
array[53728] <= 16'b0000_0000_0000_0000;
array[53729] <= 16'b0000_0000_0000_0000;
array[53730] <= 16'b0000_0000_0000_0000;
array[53731] <= 16'b0000_0000_0000_0000;
array[53732] <= 16'b0000_0000_0000_0000;
array[53733] <= 16'b0000_0000_0000_0000;
array[53734] <= 16'b0000_0000_0000_0000;
array[53735] <= 16'b0000_0000_0000_0000;
array[53736] <= 16'b0000_0000_0000_0000;
array[53737] <= 16'b0000_0000_0000_0000;
array[53738] <= 16'b0000_0000_0000_0000;
array[53739] <= 16'b0000_0000_0000_0000;
array[53740] <= 16'b0000_0000_0000_0000;
array[53741] <= 16'b0000_0000_0000_0000;
array[53742] <= 16'b0000_0000_0000_0000;
array[53743] <= 16'b0000_0000_0000_0000;
array[53744] <= 16'b0000_0000_0000_0000;
array[53745] <= 16'b0000_0000_0000_0000;
array[53746] <= 16'b0000_0000_0000_0000;
array[53747] <= 16'b0000_0000_0000_0000;
array[53748] <= 16'b0000_0000_0000_0000;
array[53749] <= 16'b0000_0000_0000_0000;
array[53750] <= 16'b0000_0000_0000_0000;
array[53751] <= 16'b0000_0000_0000_0000;
array[53752] <= 16'b0000_0000_0000_0000;
array[53753] <= 16'b0000_0000_0000_0000;
array[53754] <= 16'b0000_0000_0000_0000;
array[53755] <= 16'b0000_0000_0000_0000;
array[53756] <= 16'b0000_0000_0000_0000;
array[53757] <= 16'b0000_0000_0000_0000;
array[53758] <= 16'b0000_0000_0000_0000;
array[53759] <= 16'b0000_0000_0000_0000;
array[53760] <= 16'b0000_0000_0000_0000;
array[53761] <= 16'b0000_0000_0000_0000;
array[53762] <= 16'b0000_0000_0000_0000;
array[53763] <= 16'b0000_0000_0000_0000;
array[53764] <= 16'b0000_0000_0000_0000;
array[53765] <= 16'b0000_0000_0000_0000;
array[53766] <= 16'b0000_0000_0000_0000;
array[53767] <= 16'b0000_0000_0000_0000;
array[53768] <= 16'b0000_0000_0000_0000;
array[53769] <= 16'b0000_0000_0000_0000;
array[53770] <= 16'b0000_0000_0000_0000;
array[53771] <= 16'b0000_0000_0000_0000;
array[53772] <= 16'b0000_0000_0000_0000;
array[53773] <= 16'b0000_0000_0000_0000;
array[53774] <= 16'b0000_0000_0000_0000;
array[53775] <= 16'b0000_0000_0000_0000;
array[53776] <= 16'b0000_0000_0000_0000;
array[53777] <= 16'b0000_0000_0000_0000;
array[53778] <= 16'b0000_0000_0000_0000;
array[53779] <= 16'b0000_0000_0000_0000;
array[53780] <= 16'b0000_0000_0000_0000;
array[53781] <= 16'b0000_0000_0000_0000;
array[53782] <= 16'b0000_0000_0000_0000;
array[53783] <= 16'b0000_0000_0000_0000;
array[53784] <= 16'b0000_0000_0000_0000;
array[53785] <= 16'b0000_0000_0000_0000;
array[53786] <= 16'b0000_0000_0000_0000;
array[53787] <= 16'b0000_0000_0000_0000;
array[53788] <= 16'b0000_0000_0000_0000;
array[53789] <= 16'b0000_0000_0000_0000;
array[53790] <= 16'b0000_0000_0000_0000;
array[53791] <= 16'b0000_0000_0000_0000;
array[53792] <= 16'b0000_0000_0000_0000;
array[53793] <= 16'b0000_0000_0000_0000;
array[53794] <= 16'b0000_0000_0000_0000;
array[53795] <= 16'b0000_0000_0000_0000;
array[53796] <= 16'b0000_0000_0000_0000;
array[53797] <= 16'b0000_0000_0000_0000;
array[53798] <= 16'b0000_0000_0000_0000;
array[53799] <= 16'b0000_0000_0000_0000;
array[53800] <= 16'b0000_0000_0000_0000;
array[53801] <= 16'b0000_0000_0000_0000;
array[53802] <= 16'b0000_0000_0000_0000;
array[53803] <= 16'b0000_0000_0000_0000;
array[53804] <= 16'b0000_0000_0000_0000;
array[53805] <= 16'b0000_0000_0000_0000;
array[53806] <= 16'b0000_0000_0000_0000;
array[53807] <= 16'b0000_0000_0000_0000;
array[53808] <= 16'b0000_0000_0000_0000;
array[53809] <= 16'b0000_0000_0000_0000;
array[53810] <= 16'b0000_0000_0000_0000;
array[53811] <= 16'b0000_0000_0000_0000;
array[53812] <= 16'b0000_0000_0000_0000;
array[53813] <= 16'b0000_0000_0000_0000;
array[53814] <= 16'b0000_0000_0000_0000;
array[53815] <= 16'b0000_0000_0000_0000;
array[53816] <= 16'b0000_0000_0000_0000;
array[53817] <= 16'b0000_0000_0000_0000;
array[53818] <= 16'b0000_0000_0000_0000;
array[53819] <= 16'b0000_0000_0000_0000;
array[53820] <= 16'b0000_0000_0000_0000;
array[53821] <= 16'b0000_0000_0000_0000;
array[53822] <= 16'b0000_0000_0000_0000;
array[53823] <= 16'b0000_0000_0000_0000;
array[53824] <= 16'b0000_0000_0000_0000;
array[53825] <= 16'b0000_0000_0000_0000;
array[53826] <= 16'b0000_0000_0000_0000;
array[53827] <= 16'b0000_0000_0000_0000;
array[53828] <= 16'b0000_0000_0000_0000;
array[53829] <= 16'b0000_0000_0000_0000;
array[53830] <= 16'b0000_0000_0000_0000;
array[53831] <= 16'b0000_0000_0000_0000;
array[53832] <= 16'b0000_0000_0000_0000;
array[53833] <= 16'b0000_0000_0000_0000;
array[53834] <= 16'b0000_0000_0000_0000;
array[53835] <= 16'b0000_0000_0000_0000;
array[53836] <= 16'b0000_0000_0000_0000;
array[53837] <= 16'b0000_0000_0000_0000;
array[53838] <= 16'b0000_0000_0000_0000;
array[53839] <= 16'b0000_0000_0000_0000;
array[53840] <= 16'b0000_0000_0000_0000;
array[53841] <= 16'b0000_0000_0000_0000;
array[53842] <= 16'b0000_0000_0000_0000;
array[53843] <= 16'b0000_0000_0000_0000;
array[53844] <= 16'b0000_0000_0000_0000;
array[53845] <= 16'b0000_0000_0000_0000;
array[53846] <= 16'b0000_0000_0000_0000;
array[53847] <= 16'b0000_0000_0000_0000;
array[53848] <= 16'b0000_0000_0000_0000;
array[53849] <= 16'b0000_0000_0000_0000;
array[53850] <= 16'b0000_0000_0000_0000;
array[53851] <= 16'b0000_0000_0000_0000;
array[53852] <= 16'b0000_0000_0000_0000;
array[53853] <= 16'b0000_0000_0000_0000;
array[53854] <= 16'b0000_0000_0000_0000;
array[53855] <= 16'b0000_0000_0000_0000;
array[53856] <= 16'b0000_0000_0000_0000;
array[53857] <= 16'b0000_0000_0000_0000;
array[53858] <= 16'b0000_0000_0000_0000;
array[53859] <= 16'b0000_0000_0000_0000;
array[53860] <= 16'b0000_0000_0000_0000;
array[53861] <= 16'b0000_0000_0000_0000;
array[53862] <= 16'b0000_0000_0000_0000;
array[53863] <= 16'b0000_0000_0000_0000;
array[53864] <= 16'b0000_0000_0000_0000;
array[53865] <= 16'b0000_0000_0000_0000;
array[53866] <= 16'b0000_0000_0000_0000;
array[53867] <= 16'b0000_0000_0000_0000;
array[53868] <= 16'b0000_0000_0000_0000;
array[53869] <= 16'b0000_0000_0000_0000;
array[53870] <= 16'b0000_0000_0000_0000;
array[53871] <= 16'b0000_0000_0000_0000;
array[53872] <= 16'b0000_0000_0000_0000;
array[53873] <= 16'b0000_0000_0000_0000;
array[53874] <= 16'b0000_0000_0000_0000;
array[53875] <= 16'b0000_0000_0000_0000;
array[53876] <= 16'b0000_0000_0000_0000;
array[53877] <= 16'b0000_0000_0000_0000;
array[53878] <= 16'b0000_0000_0000_0000;
array[53879] <= 16'b0000_0000_0000_0000;
array[53880] <= 16'b0000_0000_0000_0000;
array[53881] <= 16'b0000_0000_0000_0000;
array[53882] <= 16'b0000_0000_0000_0000;
array[53883] <= 16'b0000_0000_0000_0000;
array[53884] <= 16'b0000_0000_0000_0000;
array[53885] <= 16'b0000_0000_0000_0000;
array[53886] <= 16'b0000_0000_0000_0000;
array[53887] <= 16'b0000_0000_0000_0000;
array[53888] <= 16'b0000_0000_0000_0000;
array[53889] <= 16'b0000_0000_0000_0000;
array[53890] <= 16'b0000_0000_0000_0000;
array[53891] <= 16'b0000_0000_0000_0000;
array[53892] <= 16'b0000_0000_0000_0000;
array[53893] <= 16'b0000_0000_0000_0000;
array[53894] <= 16'b0000_0000_0000_0000;
array[53895] <= 16'b0000_0000_0000_0000;
array[53896] <= 16'b0000_0000_0000_0000;
array[53897] <= 16'b0000_0000_0000_0000;
array[53898] <= 16'b0000_0000_0000_0000;
array[53899] <= 16'b0000_0000_0000_0000;
array[53900] <= 16'b0000_0000_0000_0000;
array[53901] <= 16'b0000_0000_0000_0000;
array[53902] <= 16'b0000_0000_0000_0000;
array[53903] <= 16'b0000_0000_0000_0000;
array[53904] <= 16'b0000_0000_0000_0000;
array[53905] <= 16'b0000_0000_0000_0000;
array[53906] <= 16'b0000_0000_0000_0000;
array[53907] <= 16'b0000_0000_0000_0000;
array[53908] <= 16'b0000_0000_0000_0000;
array[53909] <= 16'b0000_0000_0000_0000;
array[53910] <= 16'b0000_0000_0000_0000;
array[53911] <= 16'b0000_0000_0000_0000;
array[53912] <= 16'b0000_0000_0000_0000;
array[53913] <= 16'b0000_0000_0000_0000;
array[53914] <= 16'b0000_0000_0000_0000;
array[53915] <= 16'b0000_0000_0000_0000;
array[53916] <= 16'b0000_0000_0000_0000;
array[53917] <= 16'b0000_0000_0000_0000;
array[53918] <= 16'b0000_0000_0000_0000;
array[53919] <= 16'b0000_0000_0000_0000;
array[53920] <= 16'b0000_0000_0000_0000;
array[53921] <= 16'b0000_0000_0000_0000;
array[53922] <= 16'b0000_0000_0000_0000;
array[53923] <= 16'b0000_0000_0000_0000;
array[53924] <= 16'b0000_0000_0000_0000;
array[53925] <= 16'b0000_0000_0000_0000;
array[53926] <= 16'b0000_0000_0000_0000;
array[53927] <= 16'b0000_0000_0000_0000;
array[53928] <= 16'b0000_0000_0000_0000;
array[53929] <= 16'b0000_0000_0000_0000;
array[53930] <= 16'b0000_0000_0000_0000;
array[53931] <= 16'b0000_0000_0000_0000;
array[53932] <= 16'b0000_0000_0000_0000;
array[53933] <= 16'b0000_0000_0000_0000;
array[53934] <= 16'b0000_0000_0000_0000;
array[53935] <= 16'b0000_0000_0000_0000;
array[53936] <= 16'b0000_0000_0000_0000;
array[53937] <= 16'b0000_0000_0000_0000;
array[53938] <= 16'b0000_0000_0000_0000;
array[53939] <= 16'b0000_0000_0000_0000;
array[53940] <= 16'b0000_0000_0000_0000;
array[53941] <= 16'b0000_0000_0000_0000;
array[53942] <= 16'b0000_0000_0000_0000;
array[53943] <= 16'b0000_0000_0000_0000;
array[53944] <= 16'b0000_0000_0000_0000;
array[53945] <= 16'b0000_0000_0000_0000;
array[53946] <= 16'b0000_0000_0000_0000;
array[53947] <= 16'b0000_0000_0000_0000;
array[53948] <= 16'b0000_0000_0000_0000;
array[53949] <= 16'b0000_0000_0000_0000;
array[53950] <= 16'b0000_0000_0000_0000;
array[53951] <= 16'b0000_0000_0000_0000;
array[53952] <= 16'b0000_0000_0000_0000;
array[53953] <= 16'b0000_0000_0000_0000;
array[53954] <= 16'b0000_0000_0000_0000;
array[53955] <= 16'b0000_0000_0000_0000;
array[53956] <= 16'b0000_0000_0000_0000;
array[53957] <= 16'b0000_0000_0000_0000;
array[53958] <= 16'b0000_0000_0000_0000;
array[53959] <= 16'b0000_0000_0000_0000;
array[53960] <= 16'b0000_0000_0000_0000;
array[53961] <= 16'b0000_0000_0000_0000;
array[53962] <= 16'b0000_0000_0000_0000;
array[53963] <= 16'b0000_0000_0000_0000;
array[53964] <= 16'b0000_0000_0000_0000;
array[53965] <= 16'b0000_0000_0000_0000;
array[53966] <= 16'b0000_0000_0000_0000;
array[53967] <= 16'b0000_0000_0000_0000;
array[53968] <= 16'b0000_0000_0000_0000;
array[53969] <= 16'b0000_0000_0000_0000;
array[53970] <= 16'b0000_0000_0000_0000;
array[53971] <= 16'b0000_0000_0000_0000;
array[53972] <= 16'b0000_0000_0000_0000;
array[53973] <= 16'b0000_0000_0000_0000;
array[53974] <= 16'b0000_0000_0000_0000;
array[53975] <= 16'b0000_0000_0000_0000;
array[53976] <= 16'b0000_0000_0000_0000;
array[53977] <= 16'b0000_0000_0000_0000;
array[53978] <= 16'b0000_0000_0000_0000;
array[53979] <= 16'b0000_0000_0000_0000;
array[53980] <= 16'b0000_0000_0000_0000;
array[53981] <= 16'b0000_0000_0000_0000;
array[53982] <= 16'b0000_0000_0000_0000;
array[53983] <= 16'b0000_0000_0000_0000;
array[53984] <= 16'b0000_0000_0000_0000;
array[53985] <= 16'b0000_0000_0000_0000;
array[53986] <= 16'b0000_0000_0000_0000;
array[53987] <= 16'b0000_0000_0000_0000;
array[53988] <= 16'b0000_0000_0000_0000;
array[53989] <= 16'b0000_0000_0000_0000;
array[53990] <= 16'b0000_0000_0000_0000;
array[53991] <= 16'b0000_0000_0000_0000;
array[53992] <= 16'b0000_0000_0000_0000;
array[53993] <= 16'b0000_0000_0000_0000;
array[53994] <= 16'b0000_0000_0000_0000;
array[53995] <= 16'b0000_0000_0000_0000;
array[53996] <= 16'b0000_0000_0000_0000;
array[53997] <= 16'b0000_0000_0000_0000;
array[53998] <= 16'b0000_0000_0000_0000;
array[53999] <= 16'b0000_0000_0000_0000;
array[54000] <= 16'b0000_0000_0000_0000;
array[54001] <= 16'b0000_0000_0000_0000;
array[54002] <= 16'b0000_0000_0000_0000;
array[54003] <= 16'b0000_0000_0000_0000;
array[54004] <= 16'b0000_0000_0000_0000;
array[54005] <= 16'b0000_0000_0000_0000;
array[54006] <= 16'b0000_0000_0000_0000;
array[54007] <= 16'b0000_0000_0000_0000;
array[54008] <= 16'b0000_0000_0000_0000;
array[54009] <= 16'b0000_0000_0000_0000;
array[54010] <= 16'b0000_0000_0000_0000;
array[54011] <= 16'b0000_0000_0000_0000;
array[54012] <= 16'b0000_0000_0000_0000;
array[54013] <= 16'b0000_0000_0000_0000;
array[54014] <= 16'b0000_0000_0000_0000;
array[54015] <= 16'b0000_0000_0000_0000;
array[54016] <= 16'b0000_0000_0000_0000;
array[54017] <= 16'b0000_0000_0000_0000;
array[54018] <= 16'b0000_0000_0000_0000;
array[54019] <= 16'b0000_0000_0000_0000;
array[54020] <= 16'b0000_0000_0000_0000;
array[54021] <= 16'b0000_0000_0000_0000;
array[54022] <= 16'b0000_0000_0000_0000;
array[54023] <= 16'b0000_0000_0000_0000;
array[54024] <= 16'b0000_0000_0000_0000;
array[54025] <= 16'b0000_0000_0000_0000;
array[54026] <= 16'b0000_0000_0000_0000;
array[54027] <= 16'b0000_0000_0000_0000;
array[54028] <= 16'b0000_0000_0000_0000;
array[54029] <= 16'b0000_0000_0000_0000;
array[54030] <= 16'b0000_0000_0000_0000;
array[54031] <= 16'b0000_0000_0000_0000;
array[54032] <= 16'b0000_0000_0000_0000;
array[54033] <= 16'b0000_0000_0000_0000;
array[54034] <= 16'b0000_0000_0000_0000;
array[54035] <= 16'b0000_0000_0000_0000;
array[54036] <= 16'b0000_0000_0000_0000;
array[54037] <= 16'b0000_0000_0000_0000;
array[54038] <= 16'b0000_0000_0000_0000;
array[54039] <= 16'b0000_0000_0000_0000;
array[54040] <= 16'b0000_0000_0000_0000;
array[54041] <= 16'b0000_0000_0000_0000;
array[54042] <= 16'b0000_0000_0000_0000;
array[54043] <= 16'b0000_0000_0000_0000;
array[54044] <= 16'b0000_0000_0000_0000;
array[54045] <= 16'b0000_0000_0000_0000;
array[54046] <= 16'b0000_0000_0000_0000;
array[54047] <= 16'b0000_0000_0000_0000;
array[54048] <= 16'b0000_0000_0000_0000;
array[54049] <= 16'b0000_0000_0000_0000;
array[54050] <= 16'b0000_0000_0000_0000;
array[54051] <= 16'b0000_0000_0000_0000;
array[54052] <= 16'b0000_0000_0000_0000;
array[54053] <= 16'b0000_0000_0000_0000;
array[54054] <= 16'b0000_0000_0000_0000;
array[54055] <= 16'b0000_0000_0000_0000;
array[54056] <= 16'b0000_0000_0000_0000;
array[54057] <= 16'b0000_0000_0000_0000;
array[54058] <= 16'b0000_0000_0000_0000;
array[54059] <= 16'b0000_0000_0000_0000;
array[54060] <= 16'b0000_0000_0000_0000;
array[54061] <= 16'b0000_0000_0000_0000;
array[54062] <= 16'b0000_0000_0000_0000;
array[54063] <= 16'b0000_0000_0000_0000;
array[54064] <= 16'b0000_0000_0000_0000;
array[54065] <= 16'b0000_0000_0000_0000;
array[54066] <= 16'b0000_0000_0000_0000;
array[54067] <= 16'b0000_0000_0000_0000;
array[54068] <= 16'b0000_0000_0000_0000;
array[54069] <= 16'b0000_0000_0000_0000;
array[54070] <= 16'b0000_0000_0000_0000;
array[54071] <= 16'b0000_0000_0000_0000;
array[54072] <= 16'b0000_0000_0000_0000;
array[54073] <= 16'b0000_0000_0000_0000;
array[54074] <= 16'b0000_0000_0000_0000;
array[54075] <= 16'b0000_0000_0000_0000;
array[54076] <= 16'b0000_0000_0000_0000;
array[54077] <= 16'b0000_0000_0000_0000;
array[54078] <= 16'b0000_0000_0000_0000;
array[54079] <= 16'b0000_0000_0000_0000;
array[54080] <= 16'b0000_0000_0000_0000;
array[54081] <= 16'b0000_0000_0000_0000;
array[54082] <= 16'b0000_0000_0000_0000;
array[54083] <= 16'b0000_0000_0000_0000;
array[54084] <= 16'b0000_0000_0000_0000;
array[54085] <= 16'b0000_0000_0000_0000;
array[54086] <= 16'b0000_0000_0000_0000;
array[54087] <= 16'b0000_0000_0000_0000;
array[54088] <= 16'b0000_0000_0000_0000;
array[54089] <= 16'b0000_0000_0000_0000;
array[54090] <= 16'b0000_0000_0000_0000;
array[54091] <= 16'b0000_0000_0000_0000;
array[54092] <= 16'b0000_0000_0000_0000;
array[54093] <= 16'b0000_0000_0000_0000;
array[54094] <= 16'b0000_0000_0000_0000;
array[54095] <= 16'b0000_0000_0000_0000;
array[54096] <= 16'b0000_0000_0000_0000;
array[54097] <= 16'b0000_0000_0000_0000;
array[54098] <= 16'b0000_0000_0000_0000;
array[54099] <= 16'b0000_0000_0000_0000;
array[54100] <= 16'b0000_0000_0000_0000;
array[54101] <= 16'b0000_0000_0000_0000;
array[54102] <= 16'b0000_0000_0000_0000;
array[54103] <= 16'b0000_0000_0000_0000;
array[54104] <= 16'b0000_0000_0000_0000;
array[54105] <= 16'b0000_0000_0000_0000;
array[54106] <= 16'b0000_0000_0000_0000;
array[54107] <= 16'b0000_0000_0000_0000;
array[54108] <= 16'b0000_0000_0000_0000;
array[54109] <= 16'b0000_0000_0000_0000;
array[54110] <= 16'b0000_0000_0000_0000;
array[54111] <= 16'b0000_0000_0000_0000;
array[54112] <= 16'b0000_0000_0000_0000;
array[54113] <= 16'b0000_0000_0000_0000;
array[54114] <= 16'b0000_0000_0000_0000;
array[54115] <= 16'b0000_0000_0000_0000;
array[54116] <= 16'b0000_0000_0000_0000;
array[54117] <= 16'b0000_0000_0000_0000;
array[54118] <= 16'b0000_0000_0000_0000;
array[54119] <= 16'b0000_0000_0000_0000;
array[54120] <= 16'b0000_0000_0000_0000;
array[54121] <= 16'b0000_0000_0000_0000;
array[54122] <= 16'b0000_0000_0000_0000;
array[54123] <= 16'b0000_0000_0000_0000;
array[54124] <= 16'b0000_0000_0000_0000;
array[54125] <= 16'b0000_0000_0000_0000;
array[54126] <= 16'b0000_0000_0000_0000;
array[54127] <= 16'b0000_0000_0000_0000;
array[54128] <= 16'b0000_0000_0000_0000;
array[54129] <= 16'b0000_0000_0000_0000;
array[54130] <= 16'b0000_0000_0000_0000;
array[54131] <= 16'b0000_0000_0000_0000;
array[54132] <= 16'b0000_0000_0000_0000;
array[54133] <= 16'b0000_0000_0000_0000;
array[54134] <= 16'b0000_0000_0000_0000;
array[54135] <= 16'b0000_0000_0000_0000;
array[54136] <= 16'b0000_0000_0000_0000;
array[54137] <= 16'b0000_0000_0000_0000;
array[54138] <= 16'b0000_0000_0000_0000;
array[54139] <= 16'b0000_0000_0000_0000;
array[54140] <= 16'b0000_0000_0000_0000;
array[54141] <= 16'b0000_0000_0000_0000;
array[54142] <= 16'b0000_0000_0000_0000;
array[54143] <= 16'b0000_0000_0000_0000;
array[54144] <= 16'b0000_0000_0000_0000;
array[54145] <= 16'b0000_0000_0000_0000;
array[54146] <= 16'b0000_0000_0000_0000;
array[54147] <= 16'b0000_0000_0000_0000;
array[54148] <= 16'b0000_0000_0000_0000;
array[54149] <= 16'b0000_0000_0000_0000;
array[54150] <= 16'b0000_0000_0000_0000;
array[54151] <= 16'b0000_0000_0000_0000;
array[54152] <= 16'b0000_0000_0000_0000;
array[54153] <= 16'b0000_0000_0000_0000;
array[54154] <= 16'b0000_0000_0000_0000;
array[54155] <= 16'b0000_0000_0000_0000;
array[54156] <= 16'b0000_0000_0000_0000;
array[54157] <= 16'b0000_0000_0000_0000;
array[54158] <= 16'b0000_0000_0000_0000;
array[54159] <= 16'b0000_0000_0000_0000;
array[54160] <= 16'b0000_0000_0000_0000;
array[54161] <= 16'b0000_0000_0000_0000;
array[54162] <= 16'b0000_0000_0000_0000;
array[54163] <= 16'b0000_0000_0000_0000;
array[54164] <= 16'b0000_0000_0000_0000;
array[54165] <= 16'b0000_0000_0000_0000;
array[54166] <= 16'b0000_0000_0000_0000;
array[54167] <= 16'b0000_0000_0000_0000;
array[54168] <= 16'b0000_0000_0000_0000;
array[54169] <= 16'b0000_0000_0000_0000;
array[54170] <= 16'b0000_0000_0000_0000;
array[54171] <= 16'b0000_0000_0000_0000;
array[54172] <= 16'b0000_0000_0000_0000;
array[54173] <= 16'b0000_0000_0000_0000;
array[54174] <= 16'b0000_0000_0000_0000;
array[54175] <= 16'b0000_0000_0000_0000;
array[54176] <= 16'b0000_0000_0000_0000;
array[54177] <= 16'b0000_0000_0000_0000;
array[54178] <= 16'b0000_0000_0000_0000;
array[54179] <= 16'b0000_0000_0000_0000;
array[54180] <= 16'b0000_0000_0000_0000;
array[54181] <= 16'b0000_0000_0000_0000;
array[54182] <= 16'b0000_0000_0000_0000;
array[54183] <= 16'b0000_0000_0000_0000;
array[54184] <= 16'b0000_0000_0000_0000;
array[54185] <= 16'b0000_0000_0000_0000;
array[54186] <= 16'b0000_0000_0000_0000;
array[54187] <= 16'b0000_0000_0000_0000;
array[54188] <= 16'b0000_0000_0000_0000;
array[54189] <= 16'b0000_0000_0000_0000;
array[54190] <= 16'b0000_0000_0000_0000;
array[54191] <= 16'b0000_0000_0000_0000;
array[54192] <= 16'b0000_0000_0000_0000;
array[54193] <= 16'b0000_0000_0000_0000;
array[54194] <= 16'b0000_0000_0000_0000;
array[54195] <= 16'b0000_0000_0000_0000;
array[54196] <= 16'b0000_0000_0000_0000;
array[54197] <= 16'b0000_0000_0000_0000;
array[54198] <= 16'b0000_0000_0000_0000;
array[54199] <= 16'b0000_0000_0000_0000;
array[54200] <= 16'b0000_0000_0000_0000;
array[54201] <= 16'b0000_0000_0000_0000;
array[54202] <= 16'b0000_0000_0000_0000;
array[54203] <= 16'b0000_0000_0000_0000;
array[54204] <= 16'b0000_0000_0000_0000;
array[54205] <= 16'b0000_0000_0000_0000;
array[54206] <= 16'b0000_0000_0000_0000;
array[54207] <= 16'b0000_0000_0000_0000;
array[54208] <= 16'b0000_0000_0000_0000;
array[54209] <= 16'b0000_0000_0000_0000;
array[54210] <= 16'b0000_0000_0000_0000;
array[54211] <= 16'b0000_0000_0000_0000;
array[54212] <= 16'b0000_0000_0000_0000;
array[54213] <= 16'b0000_0000_0000_0000;
array[54214] <= 16'b0000_0000_0000_0000;
array[54215] <= 16'b0000_0000_0000_0000;
array[54216] <= 16'b0000_0000_0000_0000;
array[54217] <= 16'b0000_0000_0000_0000;
array[54218] <= 16'b0000_0000_0000_0000;
array[54219] <= 16'b0000_0000_0000_0000;
array[54220] <= 16'b0000_0000_0000_0000;
array[54221] <= 16'b0000_0000_0000_0000;
array[54222] <= 16'b0000_0000_0000_0000;
array[54223] <= 16'b0000_0000_0000_0000;
array[54224] <= 16'b0000_0000_0000_0000;
array[54225] <= 16'b0000_0000_0000_0000;
array[54226] <= 16'b0000_0000_0000_0000;
array[54227] <= 16'b0000_0000_0000_0000;
array[54228] <= 16'b0000_0000_0000_0000;
array[54229] <= 16'b0000_0000_0000_0000;
array[54230] <= 16'b0000_0000_0000_0000;
array[54231] <= 16'b0000_0000_0000_0000;
array[54232] <= 16'b0000_0000_0000_0000;
array[54233] <= 16'b0000_0000_0000_0000;
array[54234] <= 16'b0000_0000_0000_0000;
array[54235] <= 16'b0000_0000_0000_0000;
array[54236] <= 16'b0000_0000_0000_0000;
array[54237] <= 16'b0000_0000_0000_0000;
array[54238] <= 16'b0000_0000_0000_0000;
array[54239] <= 16'b0000_0000_0000_0000;
array[54240] <= 16'b0000_0000_0000_0000;
array[54241] <= 16'b0000_0000_0000_0000;
array[54242] <= 16'b0000_0000_0000_0000;
array[54243] <= 16'b0000_0000_0000_0000;
array[54244] <= 16'b0000_0000_0000_0000;
array[54245] <= 16'b0000_0000_0000_0000;
array[54246] <= 16'b0000_0000_0000_0000;
array[54247] <= 16'b0000_0000_0000_0000;
array[54248] <= 16'b0000_0000_0000_0000;
array[54249] <= 16'b0000_0000_0000_0000;
array[54250] <= 16'b0000_0000_0000_0000;
array[54251] <= 16'b0000_0000_0000_0000;
array[54252] <= 16'b0000_0000_0000_0000;
array[54253] <= 16'b0000_0000_0000_0000;
array[54254] <= 16'b0000_0000_0000_0000;
array[54255] <= 16'b0000_0000_0000_0000;
array[54256] <= 16'b0000_0000_0000_0000;
array[54257] <= 16'b0000_0000_0000_0000;
array[54258] <= 16'b0000_0000_0000_0000;
array[54259] <= 16'b0000_0000_0000_0000;
array[54260] <= 16'b0000_0000_0000_0000;
array[54261] <= 16'b0000_0000_0000_0000;
array[54262] <= 16'b0000_0000_0000_0000;
array[54263] <= 16'b0000_0000_0000_0000;
array[54264] <= 16'b0000_0000_0000_0000;
array[54265] <= 16'b0000_0000_0000_0000;
array[54266] <= 16'b0000_0000_0000_0000;
array[54267] <= 16'b0000_0000_0000_0000;
array[54268] <= 16'b0000_0000_0000_0000;
array[54269] <= 16'b0000_0000_0000_0000;
array[54270] <= 16'b0000_0000_0000_0000;
array[54271] <= 16'b0000_0000_0000_0000;
array[54272] <= 16'b0000_0000_0000_0000;
array[54273] <= 16'b0000_0000_0000_0000;
array[54274] <= 16'b0000_0000_0000_0000;
array[54275] <= 16'b0000_0000_0000_0000;
array[54276] <= 16'b0000_0000_0000_0000;
array[54277] <= 16'b0000_0000_0000_0000;
array[54278] <= 16'b0000_0000_0000_0000;
array[54279] <= 16'b0000_0000_0000_0000;
array[54280] <= 16'b0000_0000_0000_0000;
array[54281] <= 16'b0000_0000_0000_0000;
array[54282] <= 16'b0000_0000_0000_0000;
array[54283] <= 16'b0000_0000_0000_0000;
array[54284] <= 16'b0000_0000_0000_0000;
array[54285] <= 16'b0000_0000_0000_0000;
array[54286] <= 16'b0000_0000_0000_0000;
array[54287] <= 16'b0000_0000_0000_0000;
array[54288] <= 16'b0000_0000_0000_0000;
array[54289] <= 16'b0000_0000_0000_0000;
array[54290] <= 16'b0000_0000_0000_0000;
array[54291] <= 16'b0000_0000_0000_0000;
array[54292] <= 16'b0000_0000_0000_0000;
array[54293] <= 16'b0000_0000_0000_0000;
array[54294] <= 16'b0000_0000_0000_0000;
array[54295] <= 16'b0000_0000_0000_0000;
array[54296] <= 16'b0000_0000_0000_0000;
array[54297] <= 16'b0000_0000_0000_0000;
array[54298] <= 16'b0000_0000_0000_0000;
array[54299] <= 16'b0000_0000_0000_0000;
array[54300] <= 16'b0000_0000_0000_0000;
array[54301] <= 16'b0000_0000_0000_0000;
array[54302] <= 16'b0000_0000_0000_0000;
array[54303] <= 16'b0000_0000_0000_0000;
array[54304] <= 16'b0000_0000_0000_0000;
array[54305] <= 16'b0000_0000_0000_0000;
array[54306] <= 16'b0000_0000_0000_0000;
array[54307] <= 16'b0000_0000_0000_0000;
array[54308] <= 16'b0000_0000_0000_0000;
array[54309] <= 16'b0000_0000_0000_0000;
array[54310] <= 16'b0000_0000_0000_0000;
array[54311] <= 16'b0000_0000_0000_0000;
array[54312] <= 16'b0000_0000_0000_0000;
array[54313] <= 16'b0000_0000_0000_0000;
array[54314] <= 16'b0000_0000_0000_0000;
array[54315] <= 16'b0000_0000_0000_0000;
array[54316] <= 16'b0000_0000_0000_0000;
array[54317] <= 16'b0000_0000_0000_0000;
array[54318] <= 16'b0000_0000_0000_0000;
array[54319] <= 16'b0000_0000_0000_0000;
array[54320] <= 16'b0000_0000_0000_0000;
array[54321] <= 16'b0000_0000_0000_0000;
array[54322] <= 16'b0000_0000_0000_0000;
array[54323] <= 16'b0000_0000_0000_0000;
array[54324] <= 16'b0000_0000_0000_0000;
array[54325] <= 16'b0000_0000_0000_0000;
array[54326] <= 16'b0000_0000_0000_0000;
array[54327] <= 16'b0000_0000_0000_0000;
array[54328] <= 16'b0000_0000_0000_0000;
array[54329] <= 16'b0000_0000_0000_0000;
array[54330] <= 16'b0000_0000_0000_0000;
array[54331] <= 16'b0000_0000_0000_0000;
array[54332] <= 16'b0000_0000_0000_0000;
array[54333] <= 16'b0000_0000_0000_0000;
array[54334] <= 16'b0000_0000_0000_0000;
array[54335] <= 16'b0000_0000_0000_0000;
array[54336] <= 16'b0000_0000_0000_0000;
array[54337] <= 16'b0000_0000_0000_0000;
array[54338] <= 16'b0000_0000_0000_0000;
array[54339] <= 16'b0000_0000_0000_0000;
array[54340] <= 16'b0000_0000_0000_0000;
array[54341] <= 16'b0000_0000_0000_0000;
array[54342] <= 16'b0000_0000_0000_0000;
array[54343] <= 16'b0000_0000_0000_0000;
array[54344] <= 16'b0000_0000_0000_0000;
array[54345] <= 16'b0000_0000_0000_0000;
array[54346] <= 16'b0000_0000_0000_0000;
array[54347] <= 16'b0000_0000_0000_0000;
array[54348] <= 16'b0000_0000_0000_0000;
array[54349] <= 16'b0000_0000_0000_0000;
array[54350] <= 16'b0000_0000_0000_0000;
array[54351] <= 16'b0000_0000_0000_0000;
array[54352] <= 16'b0000_0000_0000_0000;
array[54353] <= 16'b0000_0000_0000_0000;
array[54354] <= 16'b0000_0000_0000_0000;
array[54355] <= 16'b0000_0000_0000_0000;
array[54356] <= 16'b0000_0000_0000_0000;
array[54357] <= 16'b0000_0000_0000_0000;
array[54358] <= 16'b0000_0000_0000_0000;
array[54359] <= 16'b0000_0000_0000_0000;
array[54360] <= 16'b0000_0000_0000_0000;
array[54361] <= 16'b0000_0000_0000_0000;
array[54362] <= 16'b0000_0000_0000_0000;
array[54363] <= 16'b0000_0000_0000_0000;
array[54364] <= 16'b0000_0000_0000_0000;
array[54365] <= 16'b0000_0000_0000_0000;
array[54366] <= 16'b0000_0000_0000_0000;
array[54367] <= 16'b0000_0000_0000_0000;
array[54368] <= 16'b0000_0000_0000_0000;
array[54369] <= 16'b0000_0000_0000_0000;
array[54370] <= 16'b0000_0000_0000_0000;
array[54371] <= 16'b0000_0000_0000_0000;
array[54372] <= 16'b0000_0000_0000_0000;
array[54373] <= 16'b0000_0000_0000_0000;
array[54374] <= 16'b0000_0000_0000_0000;
array[54375] <= 16'b0000_0000_0000_0000;
array[54376] <= 16'b0000_0000_0000_0000;
array[54377] <= 16'b0000_0000_0000_0000;
array[54378] <= 16'b0000_0000_0000_0000;
array[54379] <= 16'b0000_0000_0000_0000;
array[54380] <= 16'b0000_0000_0000_0000;
array[54381] <= 16'b0000_0000_0000_0000;
array[54382] <= 16'b0000_0000_0000_0000;
array[54383] <= 16'b0000_0000_0000_0000;
array[54384] <= 16'b0000_0000_0000_0000;
array[54385] <= 16'b0000_0000_0000_0000;
array[54386] <= 16'b0000_0000_0000_0000;
array[54387] <= 16'b0000_0000_0000_0000;
array[54388] <= 16'b0000_0000_0000_0000;
array[54389] <= 16'b0000_0000_0000_0000;
array[54390] <= 16'b0000_0000_0000_0000;
array[54391] <= 16'b0000_0000_0000_0000;
array[54392] <= 16'b0000_0000_0000_0000;
array[54393] <= 16'b0000_0000_0000_0000;
array[54394] <= 16'b0000_0000_0000_0000;
array[54395] <= 16'b0000_0000_0000_0000;
array[54396] <= 16'b0000_0000_0000_0000;
array[54397] <= 16'b0000_0000_0000_0000;
array[54398] <= 16'b0000_0000_0000_0000;
array[54399] <= 16'b0000_0000_0000_0000;
array[54400] <= 16'b0000_0000_0000_0000;
array[54401] <= 16'b0000_0000_0000_0000;
array[54402] <= 16'b0000_0000_0000_0000;
array[54403] <= 16'b0000_0000_0000_0000;
array[54404] <= 16'b0000_0000_0000_0000;
array[54405] <= 16'b0000_0000_0000_0000;
array[54406] <= 16'b0000_0000_0000_0000;
array[54407] <= 16'b0000_0000_0000_0000;
array[54408] <= 16'b0000_0000_0000_0000;
array[54409] <= 16'b0000_0000_0000_0000;
array[54410] <= 16'b0000_0000_0000_0000;
array[54411] <= 16'b0000_0000_0000_0000;
array[54412] <= 16'b0000_0000_0000_0000;
array[54413] <= 16'b0000_0000_0000_0000;
array[54414] <= 16'b0000_0000_0000_0000;
array[54415] <= 16'b0000_0000_0000_0000;
array[54416] <= 16'b0000_0000_0000_0000;
array[54417] <= 16'b0000_0000_0000_0000;
array[54418] <= 16'b0000_0000_0000_0000;
array[54419] <= 16'b0000_0000_0000_0000;
array[54420] <= 16'b0000_0000_0000_0000;
array[54421] <= 16'b0000_0000_0000_0000;
array[54422] <= 16'b0000_0000_0000_0000;
array[54423] <= 16'b0000_0000_0000_0000;
array[54424] <= 16'b0000_0000_0000_0000;
array[54425] <= 16'b0000_0000_0000_0000;
array[54426] <= 16'b0000_0000_0000_0000;
array[54427] <= 16'b0000_0000_0000_0000;
array[54428] <= 16'b0000_0000_0000_0000;
array[54429] <= 16'b0000_0000_0000_0000;
array[54430] <= 16'b0000_0000_0000_0000;
array[54431] <= 16'b0000_0000_0000_0000;
array[54432] <= 16'b0000_0000_0000_0000;
array[54433] <= 16'b0000_0000_0000_0000;
array[54434] <= 16'b0000_0000_0000_0000;
array[54435] <= 16'b0000_0000_0000_0000;
array[54436] <= 16'b0000_0000_0000_0000;
array[54437] <= 16'b0000_0000_0000_0000;
array[54438] <= 16'b0000_0000_0000_0000;
array[54439] <= 16'b0000_0000_0000_0000;
array[54440] <= 16'b0000_0000_0000_0000;
array[54441] <= 16'b0000_0000_0000_0000;
array[54442] <= 16'b0000_0000_0000_0000;
array[54443] <= 16'b0000_0000_0000_0000;
array[54444] <= 16'b0000_0000_0000_0000;
array[54445] <= 16'b0000_0000_0000_0000;
array[54446] <= 16'b0000_0000_0000_0000;
array[54447] <= 16'b0000_0000_0000_0000;
array[54448] <= 16'b0000_0000_0000_0000;
array[54449] <= 16'b0000_0000_0000_0000;
array[54450] <= 16'b0000_0000_0000_0000;
array[54451] <= 16'b0000_0000_0000_0000;
array[54452] <= 16'b0000_0000_0000_0000;
array[54453] <= 16'b0000_0000_0000_0000;
array[54454] <= 16'b0000_0000_0000_0000;
array[54455] <= 16'b0000_0000_0000_0000;
array[54456] <= 16'b0000_0000_0000_0000;
array[54457] <= 16'b0000_0000_0000_0000;
array[54458] <= 16'b0000_0000_0000_0000;
array[54459] <= 16'b0000_0000_0000_0000;
array[54460] <= 16'b0000_0000_0000_0000;
array[54461] <= 16'b0000_0000_0000_0000;
array[54462] <= 16'b0000_0000_0000_0000;
array[54463] <= 16'b0000_0000_0000_0000;
array[54464] <= 16'b0000_0000_0000_0000;
array[54465] <= 16'b0000_0000_0000_0000;
array[54466] <= 16'b0000_0000_0000_0000;
array[54467] <= 16'b0000_0000_0000_0000;
array[54468] <= 16'b0000_0000_0000_0000;
array[54469] <= 16'b0000_0000_0000_0000;
array[54470] <= 16'b0000_0000_0000_0000;
array[54471] <= 16'b0000_0000_0000_0000;
array[54472] <= 16'b0000_0000_0000_0000;
array[54473] <= 16'b0000_0000_0000_0000;
array[54474] <= 16'b0000_0000_0000_0000;
array[54475] <= 16'b0000_0000_0000_0000;
array[54476] <= 16'b0000_0000_0000_0000;
array[54477] <= 16'b0000_0000_0000_0000;
array[54478] <= 16'b0000_0000_0000_0000;
array[54479] <= 16'b0000_0000_0000_0000;
array[54480] <= 16'b0000_0000_0000_0000;
array[54481] <= 16'b0000_0000_0000_0000;
array[54482] <= 16'b0000_0000_0000_0000;
array[54483] <= 16'b0000_0000_0000_0000;
array[54484] <= 16'b0000_0000_0000_0000;
array[54485] <= 16'b0000_0000_0000_0000;
array[54486] <= 16'b0000_0000_0000_0000;
array[54487] <= 16'b0000_0000_0000_0000;
array[54488] <= 16'b0000_0000_0000_0000;
array[54489] <= 16'b0000_0000_0000_0000;
array[54490] <= 16'b0000_0000_0000_0000;
array[54491] <= 16'b0000_0000_0000_0000;
array[54492] <= 16'b0000_0000_0000_0000;
array[54493] <= 16'b0000_0000_0000_0000;
array[54494] <= 16'b0000_0000_0000_0000;
array[54495] <= 16'b0000_0000_0000_0000;
array[54496] <= 16'b0000_0000_0000_0000;
array[54497] <= 16'b0000_0000_0000_0000;
array[54498] <= 16'b0000_0000_0000_0000;
array[54499] <= 16'b0000_0000_0000_0000;
array[54500] <= 16'b0000_0000_0000_0000;
array[54501] <= 16'b0000_0000_0000_0000;
array[54502] <= 16'b0000_0000_0000_0000;
array[54503] <= 16'b0000_0000_0000_0000;
array[54504] <= 16'b0000_0000_0000_0000;
array[54505] <= 16'b0000_0000_0000_0000;
array[54506] <= 16'b0000_0000_0000_0000;
array[54507] <= 16'b0000_0000_0000_0000;
array[54508] <= 16'b0000_0000_0000_0000;
array[54509] <= 16'b0000_0000_0000_0000;
array[54510] <= 16'b0000_0000_0000_0000;
array[54511] <= 16'b0000_0000_0000_0000;
array[54512] <= 16'b0000_0000_0000_0000;
array[54513] <= 16'b0000_0000_0000_0000;
array[54514] <= 16'b0000_0000_0000_0000;
array[54515] <= 16'b0000_0000_0000_0000;
array[54516] <= 16'b0000_0000_0000_0000;
array[54517] <= 16'b0000_0000_0000_0000;
array[54518] <= 16'b0000_0000_0000_0000;
array[54519] <= 16'b0000_0000_0000_0000;
array[54520] <= 16'b0000_0000_0000_0000;
array[54521] <= 16'b0000_0000_0000_0000;
array[54522] <= 16'b0000_0000_0000_0000;
array[54523] <= 16'b0000_0000_0000_0000;
array[54524] <= 16'b0000_0000_0000_0000;
array[54525] <= 16'b0000_0000_0000_0000;
array[54526] <= 16'b0000_0000_0000_0000;
array[54527] <= 16'b0000_0000_0000_0000;
array[54528] <= 16'b0000_0000_0000_0000;
array[54529] <= 16'b0000_0000_0000_0000;
array[54530] <= 16'b0000_0000_0000_0000;
array[54531] <= 16'b0000_0000_0000_0000;
array[54532] <= 16'b0000_0000_0000_0000;
array[54533] <= 16'b0000_0000_0000_0000;
array[54534] <= 16'b0000_0000_0000_0000;
array[54535] <= 16'b0000_0000_0000_0000;
array[54536] <= 16'b0000_0000_0000_0000;
array[54537] <= 16'b0000_0000_0000_0000;
array[54538] <= 16'b0000_0000_0000_0000;
array[54539] <= 16'b0000_0000_0000_0000;
array[54540] <= 16'b0000_0000_0000_0000;
array[54541] <= 16'b0000_0000_0000_0000;
array[54542] <= 16'b0000_0000_0000_0000;
array[54543] <= 16'b0000_0000_0000_0000;
array[54544] <= 16'b0000_0000_0000_0000;
array[54545] <= 16'b0000_0000_0000_0000;
array[54546] <= 16'b0000_0000_0000_0000;
array[54547] <= 16'b0000_0000_0000_0000;
array[54548] <= 16'b0000_0000_0000_0000;
array[54549] <= 16'b0000_0000_0000_0000;
array[54550] <= 16'b0000_0000_0000_0000;
array[54551] <= 16'b0000_0000_0000_0000;
array[54552] <= 16'b0000_0000_0000_0000;
array[54553] <= 16'b0000_0000_0000_0000;
array[54554] <= 16'b0000_0000_0000_0000;
array[54555] <= 16'b0000_0000_0000_0000;
array[54556] <= 16'b0000_0000_0000_0000;
array[54557] <= 16'b0000_0000_0000_0000;
array[54558] <= 16'b0000_0000_0000_0000;
array[54559] <= 16'b0000_0000_0000_0000;
array[54560] <= 16'b0000_0000_0000_0000;
array[54561] <= 16'b0000_0000_0000_0000;
array[54562] <= 16'b0000_0000_0000_0000;
array[54563] <= 16'b0000_0000_0000_0000;
array[54564] <= 16'b0000_0000_0000_0000;
array[54565] <= 16'b0000_0000_0000_0000;
array[54566] <= 16'b0000_0000_0000_0000;
array[54567] <= 16'b0000_0000_0000_0000;
array[54568] <= 16'b0000_0000_0000_0000;
array[54569] <= 16'b0000_0000_0000_0000;
array[54570] <= 16'b0000_0000_0000_0000;
array[54571] <= 16'b0000_0000_0000_0000;
array[54572] <= 16'b0000_0000_0000_0000;
array[54573] <= 16'b0000_0000_0000_0000;
array[54574] <= 16'b0000_0000_0000_0000;
array[54575] <= 16'b0000_0000_0000_0000;
array[54576] <= 16'b0000_0000_0000_0000;
array[54577] <= 16'b0000_0000_0000_0000;
array[54578] <= 16'b0000_0000_0000_0000;
array[54579] <= 16'b0000_0000_0000_0000;
array[54580] <= 16'b0000_0000_0000_0000;
array[54581] <= 16'b0000_0000_0000_0000;
array[54582] <= 16'b0000_0000_0000_0000;
array[54583] <= 16'b0000_0000_0000_0000;
array[54584] <= 16'b0000_0000_0000_0000;
array[54585] <= 16'b0000_0000_0000_0000;
array[54586] <= 16'b0000_0000_0000_0000;
array[54587] <= 16'b0000_0000_0000_0000;
array[54588] <= 16'b0000_0000_0000_0000;
array[54589] <= 16'b0000_0000_0000_0000;
array[54590] <= 16'b0000_0000_0000_0000;
array[54591] <= 16'b0000_0000_0000_0000;
array[54592] <= 16'b0000_0000_0000_0000;
array[54593] <= 16'b0000_0000_0000_0000;
array[54594] <= 16'b0000_0000_0000_0000;
array[54595] <= 16'b0000_0000_0000_0000;
array[54596] <= 16'b0000_0000_0000_0000;
array[54597] <= 16'b0000_0000_0000_0000;
array[54598] <= 16'b0000_0000_0000_0000;
array[54599] <= 16'b0000_0000_0000_0000;
array[54600] <= 16'b0000_0000_0000_0000;
array[54601] <= 16'b0000_0000_0000_0000;
array[54602] <= 16'b0000_0000_0000_0000;
array[54603] <= 16'b0000_0000_0000_0000;
array[54604] <= 16'b0000_0000_0000_0000;
array[54605] <= 16'b0000_0000_0000_0000;
array[54606] <= 16'b0000_0000_0000_0000;
array[54607] <= 16'b0000_0000_0000_0000;
array[54608] <= 16'b0000_0000_0000_0000;
array[54609] <= 16'b0000_0000_0000_0000;
array[54610] <= 16'b0000_0000_0000_0000;
array[54611] <= 16'b0000_0000_0000_0000;
array[54612] <= 16'b0000_0000_0000_0000;
array[54613] <= 16'b0000_0000_0000_0000;
array[54614] <= 16'b0000_0000_0000_0000;
array[54615] <= 16'b0000_0000_0000_0000;
array[54616] <= 16'b0000_0000_0000_0000;
array[54617] <= 16'b0000_0000_0000_0000;
array[54618] <= 16'b0000_0000_0000_0000;
array[54619] <= 16'b0000_0000_0000_0000;
array[54620] <= 16'b0000_0000_0000_0000;
array[54621] <= 16'b0000_0000_0000_0000;
array[54622] <= 16'b0000_0000_0000_0000;
array[54623] <= 16'b0000_0000_0000_0000;
array[54624] <= 16'b0000_0000_0000_0000;
array[54625] <= 16'b0000_0000_0000_0000;
array[54626] <= 16'b0000_0000_0000_0000;
array[54627] <= 16'b0000_0000_0000_0000;
array[54628] <= 16'b0000_0000_0000_0000;
array[54629] <= 16'b0000_0000_0000_0000;
array[54630] <= 16'b0000_0000_0000_0000;
array[54631] <= 16'b0000_0000_0000_0000;
array[54632] <= 16'b0000_0000_0000_0000;
array[54633] <= 16'b0000_0000_0000_0000;
array[54634] <= 16'b0000_0000_0000_0000;
array[54635] <= 16'b0000_0000_0000_0000;
array[54636] <= 16'b0000_0000_0000_0000;
array[54637] <= 16'b0000_0000_0000_0000;
array[54638] <= 16'b0000_0000_0000_0000;
array[54639] <= 16'b0000_0000_0000_0000;
array[54640] <= 16'b0000_0000_0000_0000;
array[54641] <= 16'b0000_0000_0000_0000;
array[54642] <= 16'b0000_0000_0000_0000;
array[54643] <= 16'b0000_0000_0000_0000;
array[54644] <= 16'b0000_0000_0000_0000;
array[54645] <= 16'b0000_0000_0000_0000;
array[54646] <= 16'b0000_0000_0000_0000;
array[54647] <= 16'b0000_0000_0000_0000;
array[54648] <= 16'b0000_0000_0000_0000;
array[54649] <= 16'b0000_0000_0000_0000;
array[54650] <= 16'b0000_0000_0000_0000;
array[54651] <= 16'b0000_0000_0000_0000;
array[54652] <= 16'b0000_0000_0000_0000;
array[54653] <= 16'b0000_0000_0000_0000;
array[54654] <= 16'b0000_0000_0000_0000;
array[54655] <= 16'b0000_0000_0000_0000;
array[54656] <= 16'b0000_0000_0000_0000;
array[54657] <= 16'b0000_0000_0000_0000;
array[54658] <= 16'b0000_0000_0000_0000;
array[54659] <= 16'b0000_0000_0000_0000;
array[54660] <= 16'b0000_0000_0000_0000;
array[54661] <= 16'b0000_0000_0000_0000;
array[54662] <= 16'b0000_0000_0000_0000;
array[54663] <= 16'b0000_0000_0000_0000;
array[54664] <= 16'b0000_0000_0000_0000;
array[54665] <= 16'b0000_0000_0000_0000;
array[54666] <= 16'b0000_0000_0000_0000;
array[54667] <= 16'b0000_0000_0000_0000;
array[54668] <= 16'b0000_0000_0000_0000;
array[54669] <= 16'b0000_0000_0000_0000;
array[54670] <= 16'b0000_0000_0000_0000;
array[54671] <= 16'b0000_0000_0000_0000;
array[54672] <= 16'b0000_0000_0000_0000;
array[54673] <= 16'b0000_0000_0000_0000;
array[54674] <= 16'b0000_0000_0000_0000;
array[54675] <= 16'b0000_0000_0000_0000;
array[54676] <= 16'b0000_0000_0000_0000;
array[54677] <= 16'b0000_0000_0000_0000;
array[54678] <= 16'b0000_0000_0000_0000;
array[54679] <= 16'b0000_0000_0000_0000;
array[54680] <= 16'b0000_0000_0000_0000;
array[54681] <= 16'b0000_0000_0000_0000;
array[54682] <= 16'b0000_0000_0000_0000;
array[54683] <= 16'b0000_0000_0000_0000;
array[54684] <= 16'b0000_0000_0000_0000;
array[54685] <= 16'b0000_0000_0000_0000;
array[54686] <= 16'b0000_0000_0000_0000;
array[54687] <= 16'b0000_0000_0000_0000;
array[54688] <= 16'b0000_0000_0000_0000;
array[54689] <= 16'b0000_0000_0000_0000;
array[54690] <= 16'b0000_0000_0000_0000;
array[54691] <= 16'b0000_0000_0000_0000;
array[54692] <= 16'b0000_0000_0000_0000;
array[54693] <= 16'b0000_0000_0000_0000;
array[54694] <= 16'b0000_0000_0000_0000;
array[54695] <= 16'b0000_0000_0000_0000;
array[54696] <= 16'b0000_0000_0000_0000;
array[54697] <= 16'b0000_0000_0000_0000;
array[54698] <= 16'b0000_0000_0000_0000;
array[54699] <= 16'b0000_0000_0000_0000;
array[54700] <= 16'b0000_0000_0000_0000;
array[54701] <= 16'b0000_0000_0000_0000;
array[54702] <= 16'b0000_0000_0000_0000;
array[54703] <= 16'b0000_0000_0000_0000;
array[54704] <= 16'b0000_0000_0000_0000;
array[54705] <= 16'b0000_0000_0000_0000;
array[54706] <= 16'b0000_0000_0000_0000;
array[54707] <= 16'b0000_0000_0000_0000;
array[54708] <= 16'b0000_0000_0000_0000;
array[54709] <= 16'b0000_0000_0000_0000;
array[54710] <= 16'b0000_0000_0000_0000;
array[54711] <= 16'b0000_0000_0000_0000;
array[54712] <= 16'b0000_0000_0000_0000;
array[54713] <= 16'b0000_0000_0000_0000;
array[54714] <= 16'b0000_0000_0000_0000;
array[54715] <= 16'b0000_0000_0000_0000;
array[54716] <= 16'b0000_0000_0000_0000;
array[54717] <= 16'b0000_0000_0000_0000;
array[54718] <= 16'b0000_0000_0000_0000;
array[54719] <= 16'b0000_0000_0000_0000;
array[54720] <= 16'b0000_0000_0000_0000;
array[54721] <= 16'b0000_0000_0000_0000;
array[54722] <= 16'b0000_0000_0000_0000;
array[54723] <= 16'b0000_0000_0000_0000;
array[54724] <= 16'b0000_0000_0000_0000;
array[54725] <= 16'b0000_0000_0000_0000;
array[54726] <= 16'b0000_0000_0000_0000;
array[54727] <= 16'b0000_0000_0000_0000;
array[54728] <= 16'b0000_0000_0000_0000;
array[54729] <= 16'b0000_0000_0000_0000;
array[54730] <= 16'b0000_0000_0000_0000;
array[54731] <= 16'b0000_0000_0000_0000;
array[54732] <= 16'b0000_0000_0000_0000;
array[54733] <= 16'b0000_0000_0000_0000;
array[54734] <= 16'b0000_0000_0000_0000;
array[54735] <= 16'b0000_0000_0000_0000;
array[54736] <= 16'b0000_0000_0000_0000;
array[54737] <= 16'b0000_0000_0000_0000;
array[54738] <= 16'b0000_0000_0000_0000;
array[54739] <= 16'b0000_0000_0000_0000;
array[54740] <= 16'b0000_0000_0000_0000;
array[54741] <= 16'b0000_0000_0000_0000;
array[54742] <= 16'b0000_0000_0000_0000;
array[54743] <= 16'b0000_0000_0000_0000;
array[54744] <= 16'b0000_0000_0000_0000;
array[54745] <= 16'b0000_0000_0000_0000;
array[54746] <= 16'b0000_0000_0000_0000;
array[54747] <= 16'b0000_0000_0000_0000;
array[54748] <= 16'b0000_0000_0000_0000;
array[54749] <= 16'b0000_0000_0000_0000;
array[54750] <= 16'b0000_0000_0000_0000;
array[54751] <= 16'b0000_0000_0000_0000;
array[54752] <= 16'b0000_0000_0000_0000;
array[54753] <= 16'b0000_0000_0000_0000;
array[54754] <= 16'b0000_0000_0000_0000;
array[54755] <= 16'b0000_0000_0000_0000;
array[54756] <= 16'b0000_0000_0000_0000;
array[54757] <= 16'b0000_0000_0000_0000;
array[54758] <= 16'b0000_0000_0000_0000;
array[54759] <= 16'b0000_0000_0000_0000;
array[54760] <= 16'b0000_0000_0000_0000;
array[54761] <= 16'b0000_0000_0000_0000;
array[54762] <= 16'b0000_0000_0000_0000;
array[54763] <= 16'b0000_0000_0000_0000;
array[54764] <= 16'b0000_0000_0000_0000;
array[54765] <= 16'b0000_0000_0000_0000;
array[54766] <= 16'b0000_0000_0000_0000;
array[54767] <= 16'b0000_0000_0000_0000;
array[54768] <= 16'b0000_0000_0000_0000;
array[54769] <= 16'b0000_0000_0000_0000;
array[54770] <= 16'b0000_0000_0000_0000;
array[54771] <= 16'b0000_0000_0000_0000;
array[54772] <= 16'b0000_0000_0000_0000;
array[54773] <= 16'b0000_0000_0000_0000;
array[54774] <= 16'b0000_0000_0000_0000;
array[54775] <= 16'b0000_0000_0000_0000;
array[54776] <= 16'b0000_0000_0000_0000;
array[54777] <= 16'b0000_0000_0000_0000;
array[54778] <= 16'b0000_0000_0000_0000;
array[54779] <= 16'b0000_0000_0000_0000;
array[54780] <= 16'b0000_0000_0000_0000;
array[54781] <= 16'b0000_0000_0000_0000;
array[54782] <= 16'b0000_0000_0000_0000;
array[54783] <= 16'b0000_0000_0000_0000;
array[54784] <= 16'b0000_0000_0000_0000;
array[54785] <= 16'b0000_0000_0000_0000;
array[54786] <= 16'b0000_0000_0000_0000;
array[54787] <= 16'b0000_0000_0000_0000;
array[54788] <= 16'b0000_0000_0000_0000;
array[54789] <= 16'b0000_0000_0000_0000;
array[54790] <= 16'b0000_0000_0000_0000;
array[54791] <= 16'b0000_0000_0000_0000;
array[54792] <= 16'b0000_0000_0000_0000;
array[54793] <= 16'b0000_0000_0000_0000;
array[54794] <= 16'b0000_0000_0000_0000;
array[54795] <= 16'b0000_0000_0000_0000;
array[54796] <= 16'b0000_0000_0000_0000;
array[54797] <= 16'b0000_0000_0000_0000;
array[54798] <= 16'b0000_0000_0000_0000;
array[54799] <= 16'b0000_0000_0000_0000;
array[54800] <= 16'b0000_0000_0000_0000;
array[54801] <= 16'b0000_0000_0000_0000;
array[54802] <= 16'b0000_0000_0000_0000;
array[54803] <= 16'b0000_0000_0000_0000;
array[54804] <= 16'b0000_0000_0000_0000;
array[54805] <= 16'b0000_0000_0000_0000;
array[54806] <= 16'b0000_0000_0000_0000;
array[54807] <= 16'b0000_0000_0000_0000;
array[54808] <= 16'b0000_0000_0000_0000;
array[54809] <= 16'b0000_0000_0000_0000;
array[54810] <= 16'b0000_0000_0000_0000;
array[54811] <= 16'b0000_0000_0000_0000;
array[54812] <= 16'b0000_0000_0000_0000;
array[54813] <= 16'b0000_0000_0000_0000;
array[54814] <= 16'b0000_0000_0000_0000;
array[54815] <= 16'b0000_0000_0000_0000;
array[54816] <= 16'b0000_0000_0000_0000;
array[54817] <= 16'b0000_0000_0000_0000;
array[54818] <= 16'b0000_0000_0000_0000;
array[54819] <= 16'b0000_0000_0000_0000;
array[54820] <= 16'b0000_0000_0000_0000;
array[54821] <= 16'b0000_0000_0000_0000;
array[54822] <= 16'b0000_0000_0000_0000;
array[54823] <= 16'b0000_0000_0000_0000;
array[54824] <= 16'b0000_0000_0000_0000;
array[54825] <= 16'b0000_0000_0000_0000;
array[54826] <= 16'b0000_0000_0000_0000;
array[54827] <= 16'b0000_0000_0000_0000;
array[54828] <= 16'b0000_0000_0000_0000;
array[54829] <= 16'b0000_0000_0000_0000;
array[54830] <= 16'b0000_0000_0000_0000;
array[54831] <= 16'b0000_0000_0000_0000;
array[54832] <= 16'b0000_0000_0000_0000;
array[54833] <= 16'b0000_0000_0000_0000;
array[54834] <= 16'b0000_0000_0000_0000;
array[54835] <= 16'b0000_0000_0000_0000;
array[54836] <= 16'b0000_0000_0000_0000;
array[54837] <= 16'b0000_0000_0000_0000;
array[54838] <= 16'b0000_0000_0000_0000;
array[54839] <= 16'b0000_0000_0000_0000;
array[54840] <= 16'b0000_0000_0000_0000;
array[54841] <= 16'b0000_0000_0000_0000;
array[54842] <= 16'b0000_0000_0000_0000;
array[54843] <= 16'b0000_0000_0000_0000;
array[54844] <= 16'b0000_0000_0000_0000;
array[54845] <= 16'b0000_0000_0000_0000;
array[54846] <= 16'b0000_0000_0000_0000;
array[54847] <= 16'b0000_0000_0000_0000;
array[54848] <= 16'b0000_0000_0000_0000;
array[54849] <= 16'b0000_0000_0000_0000;
array[54850] <= 16'b0000_0000_0000_0000;
array[54851] <= 16'b0000_0000_0000_0000;
array[54852] <= 16'b0000_0000_0000_0000;
array[54853] <= 16'b0000_0000_0000_0000;
array[54854] <= 16'b0000_0000_0000_0000;
array[54855] <= 16'b0000_0000_0000_0000;
array[54856] <= 16'b0000_0000_0000_0000;
array[54857] <= 16'b0000_0000_0000_0000;
array[54858] <= 16'b0000_0000_0000_0000;
array[54859] <= 16'b0000_0000_0000_0000;
array[54860] <= 16'b0000_0000_0000_0000;
array[54861] <= 16'b0000_0000_0000_0000;
array[54862] <= 16'b0000_0000_0000_0000;
array[54863] <= 16'b0000_0000_0000_0000;
array[54864] <= 16'b0000_0000_0000_0000;
array[54865] <= 16'b0000_0000_0000_0000;
array[54866] <= 16'b0000_0000_0000_0000;
array[54867] <= 16'b0000_0000_0000_0000;
array[54868] <= 16'b0000_0000_0000_0000;
array[54869] <= 16'b0000_0000_0000_0000;
array[54870] <= 16'b0000_0000_0000_0000;
array[54871] <= 16'b0000_0000_0000_0000;
array[54872] <= 16'b0000_0000_0000_0000;
array[54873] <= 16'b0000_0000_0000_0000;
array[54874] <= 16'b0000_0000_0000_0000;
array[54875] <= 16'b0000_0000_0000_0000;
array[54876] <= 16'b0000_0000_0000_0000;
array[54877] <= 16'b0000_0000_0000_0000;
array[54878] <= 16'b0000_0000_0000_0000;
array[54879] <= 16'b0000_0000_0000_0000;
array[54880] <= 16'b0000_0000_0000_0000;
array[54881] <= 16'b0000_0000_0000_0000;
array[54882] <= 16'b0000_0000_0000_0000;
array[54883] <= 16'b0000_0000_0000_0000;
array[54884] <= 16'b0000_0000_0000_0000;
array[54885] <= 16'b0000_0000_0000_0000;
array[54886] <= 16'b0000_0000_0000_0000;
array[54887] <= 16'b0000_0000_0000_0000;
array[54888] <= 16'b0000_0000_0000_0000;
array[54889] <= 16'b0000_0000_0000_0000;
array[54890] <= 16'b0000_0000_0000_0000;
array[54891] <= 16'b0000_0000_0000_0000;
array[54892] <= 16'b0000_0000_0000_0000;
array[54893] <= 16'b0000_0000_0000_0000;
array[54894] <= 16'b0000_0000_0000_0000;
array[54895] <= 16'b0000_0000_0000_0000;
array[54896] <= 16'b0000_0000_0000_0000;
array[54897] <= 16'b0000_0000_0000_0000;
array[54898] <= 16'b0000_0000_0000_0000;
array[54899] <= 16'b0000_0000_0000_0000;
array[54900] <= 16'b0000_0000_0000_0000;
array[54901] <= 16'b0000_0000_0000_0000;
array[54902] <= 16'b0000_0000_0000_0000;
array[54903] <= 16'b0000_0000_0000_0000;
array[54904] <= 16'b0000_0000_0000_0000;
array[54905] <= 16'b0000_0000_0000_0000;
array[54906] <= 16'b0000_0000_0000_0000;
array[54907] <= 16'b0000_0000_0000_0000;
array[54908] <= 16'b0000_0000_0000_0000;
array[54909] <= 16'b0000_0000_0000_0000;
array[54910] <= 16'b0000_0000_0000_0000;
array[54911] <= 16'b0000_0000_0000_0000;
array[54912] <= 16'b0000_0000_0000_0000;
array[54913] <= 16'b0000_0000_0000_0000;
array[54914] <= 16'b0000_0000_0000_0000;
array[54915] <= 16'b0000_0000_0000_0000;
array[54916] <= 16'b0000_0000_0000_0000;
array[54917] <= 16'b0000_0000_0000_0000;
array[54918] <= 16'b0000_0000_0000_0000;
array[54919] <= 16'b0000_0000_0000_0000;
array[54920] <= 16'b0000_0000_0000_0000;
array[54921] <= 16'b0000_0000_0000_0000;
array[54922] <= 16'b0000_0000_0000_0000;
array[54923] <= 16'b0000_0000_0000_0000;
array[54924] <= 16'b0000_0000_0000_0000;
array[54925] <= 16'b0000_0000_0000_0000;
array[54926] <= 16'b0000_0000_0000_0000;
array[54927] <= 16'b0000_0000_0000_0000;
array[54928] <= 16'b0000_0000_0000_0000;
array[54929] <= 16'b0000_0000_0000_0000;
array[54930] <= 16'b0000_0000_0000_0000;
array[54931] <= 16'b0000_0000_0000_0000;
array[54932] <= 16'b0000_0000_0000_0000;
array[54933] <= 16'b0000_0000_0000_0000;
array[54934] <= 16'b0000_0000_0000_0000;
array[54935] <= 16'b0000_0000_0000_0000;
array[54936] <= 16'b0000_0000_0000_0000;
array[54937] <= 16'b0000_0000_0000_0000;
array[54938] <= 16'b0000_0000_0000_0000;
array[54939] <= 16'b0000_0000_0000_0000;
array[54940] <= 16'b0000_0000_0000_0000;
array[54941] <= 16'b0000_0000_0000_0000;
array[54942] <= 16'b0000_0000_0000_0000;
array[54943] <= 16'b0000_0000_0000_0000;
array[54944] <= 16'b0000_0000_0000_0000;
array[54945] <= 16'b0000_0000_0000_0000;
array[54946] <= 16'b0000_0000_0000_0000;
array[54947] <= 16'b0000_0000_0000_0000;
array[54948] <= 16'b0000_0000_0000_0000;
array[54949] <= 16'b0000_0000_0000_0000;
array[54950] <= 16'b0000_0000_0000_0000;
array[54951] <= 16'b0000_0000_0000_0000;
array[54952] <= 16'b0000_0000_0000_0000;
array[54953] <= 16'b0000_0000_0000_0000;
array[54954] <= 16'b0000_0000_0000_0000;
array[54955] <= 16'b0000_0000_0000_0000;
array[54956] <= 16'b0000_0000_0000_0000;
array[54957] <= 16'b0000_0000_0000_0000;
array[54958] <= 16'b0000_0000_0000_0000;
array[54959] <= 16'b0000_0000_0000_0000;
array[54960] <= 16'b0000_0000_0000_0000;
array[54961] <= 16'b0000_0000_0000_0000;
array[54962] <= 16'b0000_0000_0000_0000;
array[54963] <= 16'b0000_0000_0000_0000;
array[54964] <= 16'b0000_0000_0000_0000;
array[54965] <= 16'b0000_0000_0000_0000;
array[54966] <= 16'b0000_0000_0000_0000;
array[54967] <= 16'b0000_0000_0000_0000;
array[54968] <= 16'b0000_0000_0000_0000;
array[54969] <= 16'b0000_0000_0000_0000;
array[54970] <= 16'b0000_0000_0000_0000;
array[54971] <= 16'b0000_0000_0000_0000;
array[54972] <= 16'b0000_0000_0000_0000;
array[54973] <= 16'b0000_0000_0000_0000;
array[54974] <= 16'b0000_0000_0000_0000;
array[54975] <= 16'b0000_0000_0000_0000;
array[54976] <= 16'b0000_0000_0000_0000;
array[54977] <= 16'b0000_0000_0000_0000;
array[54978] <= 16'b0000_0000_0000_0000;
array[54979] <= 16'b0000_0000_0000_0000;
array[54980] <= 16'b0000_0000_0000_0000;
array[54981] <= 16'b0000_0000_0000_0000;
array[54982] <= 16'b0000_0000_0000_0000;
array[54983] <= 16'b0000_0000_0000_0000;
array[54984] <= 16'b0000_0000_0000_0000;
array[54985] <= 16'b0000_0000_0000_0000;
array[54986] <= 16'b0000_0000_0000_0000;
array[54987] <= 16'b0000_0000_0000_0000;
array[54988] <= 16'b0000_0000_0000_0000;
array[54989] <= 16'b0000_0000_0000_0000;
array[54990] <= 16'b0000_0000_0000_0000;
array[54991] <= 16'b0000_0000_0000_0000;
array[54992] <= 16'b0000_0000_0000_0000;
array[54993] <= 16'b0000_0000_0000_0000;
array[54994] <= 16'b0000_0000_0000_0000;
array[54995] <= 16'b0000_0000_0000_0000;
array[54996] <= 16'b0000_0000_0000_0000;
array[54997] <= 16'b0000_0000_0000_0000;
array[54998] <= 16'b0000_0000_0000_0000;
array[54999] <= 16'b0000_0000_0000_0000;
array[55000] <= 16'b0000_0000_0000_0000;
array[55001] <= 16'b0000_0000_0000_0000;
array[55002] <= 16'b0000_0000_0000_0000;
array[55003] <= 16'b0000_0000_0000_0000;
array[55004] <= 16'b0000_0000_0000_0000;
array[55005] <= 16'b0000_0000_0000_0000;
array[55006] <= 16'b0000_0000_0000_0000;
array[55007] <= 16'b0000_0000_0000_0000;
array[55008] <= 16'b0000_0000_0000_0000;
array[55009] <= 16'b0000_0000_0000_0000;
array[55010] <= 16'b0000_0000_0000_0000;
array[55011] <= 16'b0000_0000_0000_0000;
array[55012] <= 16'b0000_0000_0000_0000;
array[55013] <= 16'b0000_0000_0000_0000;
array[55014] <= 16'b0000_0000_0000_0000;
array[55015] <= 16'b0000_0000_0000_0000;
array[55016] <= 16'b0000_0000_0000_0000;
array[55017] <= 16'b0000_0000_0000_0000;
array[55018] <= 16'b0000_0000_0000_0000;
array[55019] <= 16'b0000_0000_0000_0000;
array[55020] <= 16'b0000_0000_0000_0000;
array[55021] <= 16'b0000_0000_0000_0000;
array[55022] <= 16'b0000_0000_0000_0000;
array[55023] <= 16'b0000_0000_0000_0000;
array[55024] <= 16'b0000_0000_0000_0000;
array[55025] <= 16'b0000_0000_0000_0000;
array[55026] <= 16'b0000_0000_0000_0000;
array[55027] <= 16'b0000_0000_0000_0000;
array[55028] <= 16'b0000_0000_0000_0000;
array[55029] <= 16'b0000_0000_0000_0000;
array[55030] <= 16'b0000_0000_0000_0000;
array[55031] <= 16'b0000_0000_0000_0000;
array[55032] <= 16'b0000_0000_0000_0000;
array[55033] <= 16'b0000_0000_0000_0000;
array[55034] <= 16'b0000_0000_0000_0000;
array[55035] <= 16'b0000_0000_0000_0000;
array[55036] <= 16'b0000_0000_0000_0000;
array[55037] <= 16'b0000_0000_0000_0000;
array[55038] <= 16'b0000_0000_0000_0000;
array[55039] <= 16'b0000_0000_0000_0000;
array[55040] <= 16'b0000_0000_0000_0000;
array[55041] <= 16'b0000_0000_0000_0000;
array[55042] <= 16'b0000_0000_0000_0000;
array[55043] <= 16'b0000_0000_0000_0000;
array[55044] <= 16'b0000_0000_0000_0000;
array[55045] <= 16'b0000_0000_0000_0000;
array[55046] <= 16'b0000_0000_0000_0000;
array[55047] <= 16'b0000_0000_0000_0000;
array[55048] <= 16'b0000_0000_0000_0000;
array[55049] <= 16'b0000_0000_0000_0000;
array[55050] <= 16'b0000_0000_0000_0000;
array[55051] <= 16'b0000_0000_0000_0000;
array[55052] <= 16'b0000_0000_0000_0000;
array[55053] <= 16'b0000_0000_0000_0000;
array[55054] <= 16'b0000_0000_0000_0000;
array[55055] <= 16'b0000_0000_0000_0000;
array[55056] <= 16'b0000_0000_0000_0000;
array[55057] <= 16'b0000_0000_0000_0000;
array[55058] <= 16'b0000_0000_0000_0000;
array[55059] <= 16'b0000_0000_0000_0000;
array[55060] <= 16'b0000_0000_0000_0000;
array[55061] <= 16'b0000_0000_0000_0000;
array[55062] <= 16'b0000_0000_0000_0000;
array[55063] <= 16'b0000_0000_0000_0000;
array[55064] <= 16'b0000_0000_0000_0000;
array[55065] <= 16'b0000_0000_0000_0000;
array[55066] <= 16'b0000_0000_0000_0000;
array[55067] <= 16'b0000_0000_0000_0000;
array[55068] <= 16'b0000_0000_0000_0000;
array[55069] <= 16'b0000_0000_0000_0000;
array[55070] <= 16'b0000_0000_0000_0000;
array[55071] <= 16'b0000_0000_0000_0000;
array[55072] <= 16'b0000_0000_0000_0000;
array[55073] <= 16'b0000_0000_0000_0000;
array[55074] <= 16'b0000_0000_0000_0000;
array[55075] <= 16'b0000_0000_0000_0000;
array[55076] <= 16'b0000_0000_0000_0000;
array[55077] <= 16'b0000_0000_0000_0000;
array[55078] <= 16'b0000_0000_0000_0000;
array[55079] <= 16'b0000_0000_0000_0000;
array[55080] <= 16'b0000_0000_0000_0000;
array[55081] <= 16'b0000_0000_0000_0000;
array[55082] <= 16'b0000_0000_0000_0000;
array[55083] <= 16'b0000_0000_0000_0000;
array[55084] <= 16'b0000_0000_0000_0000;
array[55085] <= 16'b0000_0000_0000_0000;
array[55086] <= 16'b0000_0000_0000_0000;
array[55087] <= 16'b0000_0000_0000_0000;
array[55088] <= 16'b0000_0000_0000_0000;
array[55089] <= 16'b0000_0000_0000_0000;
array[55090] <= 16'b0000_0000_0000_0000;
array[55091] <= 16'b0000_0000_0000_0000;
array[55092] <= 16'b0000_0000_0000_0000;
array[55093] <= 16'b0000_0000_0000_0000;
array[55094] <= 16'b0000_0000_0000_0000;
array[55095] <= 16'b0000_0000_0000_0000;
array[55096] <= 16'b0000_0000_0000_0000;
array[55097] <= 16'b0000_0000_0000_0000;
array[55098] <= 16'b0000_0000_0000_0000;
array[55099] <= 16'b0000_0000_0000_0000;
array[55100] <= 16'b0000_0000_0000_0000;
array[55101] <= 16'b0000_0000_0000_0000;
array[55102] <= 16'b0000_0000_0000_0000;
array[55103] <= 16'b0000_0000_0000_0000;
array[55104] <= 16'b0000_0000_0000_0000;
array[55105] <= 16'b0000_0000_0000_0000;
array[55106] <= 16'b0000_0000_0000_0000;
array[55107] <= 16'b0000_0000_0000_0000;
array[55108] <= 16'b0000_0000_0000_0000;
array[55109] <= 16'b0000_0000_0000_0000;
array[55110] <= 16'b0000_0000_0000_0000;
array[55111] <= 16'b0000_0000_0000_0000;
array[55112] <= 16'b0000_0000_0000_0000;
array[55113] <= 16'b0000_0000_0000_0000;
array[55114] <= 16'b0000_0000_0000_0000;
array[55115] <= 16'b0000_0000_0000_0000;
array[55116] <= 16'b0000_0000_0000_0000;
array[55117] <= 16'b0000_0000_0000_0000;
array[55118] <= 16'b0000_0000_0000_0000;
array[55119] <= 16'b0000_0000_0000_0000;
array[55120] <= 16'b0000_0000_0000_0000;
array[55121] <= 16'b0000_0000_0000_0000;
array[55122] <= 16'b0000_0000_0000_0000;
array[55123] <= 16'b0000_0000_0000_0000;
array[55124] <= 16'b0000_0000_0000_0000;
array[55125] <= 16'b0000_0000_0000_0000;
array[55126] <= 16'b0000_0000_0000_0000;
array[55127] <= 16'b0000_0000_0000_0000;
array[55128] <= 16'b0000_0000_0000_0000;
array[55129] <= 16'b0000_0000_0000_0000;
array[55130] <= 16'b0000_0000_0000_0000;
array[55131] <= 16'b0000_0000_0000_0000;
array[55132] <= 16'b0000_0000_0000_0000;
array[55133] <= 16'b0000_0000_0000_0000;
array[55134] <= 16'b0000_0000_0000_0000;
array[55135] <= 16'b0000_0000_0000_0000;
array[55136] <= 16'b0000_0000_0000_0000;
array[55137] <= 16'b0000_0000_0000_0000;
array[55138] <= 16'b0000_0000_0000_0000;
array[55139] <= 16'b0000_0000_0000_0000;
array[55140] <= 16'b0000_0000_0000_0000;
array[55141] <= 16'b0000_0000_0000_0000;
array[55142] <= 16'b0000_0000_0000_0000;
array[55143] <= 16'b0000_0000_0000_0000;
array[55144] <= 16'b0000_0000_0000_0000;
array[55145] <= 16'b0000_0000_0000_0000;
array[55146] <= 16'b0000_0000_0000_0000;
array[55147] <= 16'b0000_0000_0000_0000;
array[55148] <= 16'b0000_0000_0000_0000;
array[55149] <= 16'b0000_0000_0000_0000;
array[55150] <= 16'b0000_0000_0000_0000;
array[55151] <= 16'b0000_0000_0000_0000;
array[55152] <= 16'b0000_0000_0000_0000;
array[55153] <= 16'b0000_0000_0000_0000;
array[55154] <= 16'b0000_0000_0000_0000;
array[55155] <= 16'b0000_0000_0000_0000;
array[55156] <= 16'b0000_0000_0000_0000;
array[55157] <= 16'b0000_0000_0000_0000;
array[55158] <= 16'b0000_0000_0000_0000;
array[55159] <= 16'b0000_0000_0000_0000;
array[55160] <= 16'b0000_0000_0000_0000;
array[55161] <= 16'b0000_0000_0000_0000;
array[55162] <= 16'b0000_0000_0000_0000;
array[55163] <= 16'b0000_0000_0000_0000;
array[55164] <= 16'b0000_0000_0000_0000;
array[55165] <= 16'b0000_0000_0000_0000;
array[55166] <= 16'b0000_0000_0000_0000;
array[55167] <= 16'b0000_0000_0000_0000;
array[55168] <= 16'b0000_0000_0000_0000;
array[55169] <= 16'b0000_0000_0000_0000;
array[55170] <= 16'b0000_0000_0000_0000;
array[55171] <= 16'b0000_0000_0000_0000;
array[55172] <= 16'b0000_0000_0000_0000;
array[55173] <= 16'b0000_0000_0000_0000;
array[55174] <= 16'b0000_0000_0000_0000;
array[55175] <= 16'b0000_0000_0000_0000;
array[55176] <= 16'b0000_0000_0000_0000;
array[55177] <= 16'b0000_0000_0000_0000;
array[55178] <= 16'b0000_0000_0000_0000;
array[55179] <= 16'b0000_0000_0000_0000;
array[55180] <= 16'b0000_0000_0000_0000;
array[55181] <= 16'b0000_0000_0000_0000;
array[55182] <= 16'b0000_0000_0000_0000;
array[55183] <= 16'b0000_0000_0000_0000;
array[55184] <= 16'b0000_0000_0000_0000;
array[55185] <= 16'b0000_0000_0000_0000;
array[55186] <= 16'b0000_0000_0000_0000;
array[55187] <= 16'b0000_0000_0000_0000;
array[55188] <= 16'b0000_0000_0000_0000;
array[55189] <= 16'b0000_0000_0000_0000;
array[55190] <= 16'b0000_0000_0000_0000;
array[55191] <= 16'b0000_0000_0000_0000;
array[55192] <= 16'b0000_0000_0000_0000;
array[55193] <= 16'b0000_0000_0000_0000;
array[55194] <= 16'b0000_0000_0000_0000;
array[55195] <= 16'b0000_0000_0000_0000;
array[55196] <= 16'b0000_0000_0000_0000;
array[55197] <= 16'b0000_0000_0000_0000;
array[55198] <= 16'b0000_0000_0000_0000;
array[55199] <= 16'b0000_0000_0000_0000;
array[55200] <= 16'b0000_0000_0000_0000;
array[55201] <= 16'b0000_0000_0000_0000;
array[55202] <= 16'b0000_0000_0000_0000;
array[55203] <= 16'b0000_0000_0000_0000;
array[55204] <= 16'b0000_0000_0000_0000;
array[55205] <= 16'b0000_0000_0000_0000;
array[55206] <= 16'b0000_0000_0000_0000;
array[55207] <= 16'b0000_0000_0000_0000;
array[55208] <= 16'b0000_0000_0000_0000;
array[55209] <= 16'b0000_0000_0000_0000;
array[55210] <= 16'b0000_0000_0000_0000;
array[55211] <= 16'b0000_0000_0000_0000;
array[55212] <= 16'b0000_0000_0000_0000;
array[55213] <= 16'b0000_0000_0000_0000;
array[55214] <= 16'b0000_0000_0000_0000;
array[55215] <= 16'b0000_0000_0000_0000;
array[55216] <= 16'b0000_0000_0000_0000;
array[55217] <= 16'b0000_0000_0000_0000;
array[55218] <= 16'b0000_0000_0000_0000;
array[55219] <= 16'b0000_0000_0000_0000;
array[55220] <= 16'b0000_0000_0000_0000;
array[55221] <= 16'b0000_0000_0000_0000;
array[55222] <= 16'b0000_0000_0000_0000;
array[55223] <= 16'b0000_0000_0000_0000;
array[55224] <= 16'b0000_0000_0000_0000;
array[55225] <= 16'b0000_0000_0000_0000;
array[55226] <= 16'b0000_0000_0000_0000;
array[55227] <= 16'b0000_0000_0000_0000;
array[55228] <= 16'b0000_0000_0000_0000;
array[55229] <= 16'b0000_0000_0000_0000;
array[55230] <= 16'b0000_0000_0000_0000;
array[55231] <= 16'b0000_0000_0000_0000;
array[55232] <= 16'b0000_0000_0000_0000;
array[55233] <= 16'b0000_0000_0000_0000;
array[55234] <= 16'b0000_0000_0000_0000;
array[55235] <= 16'b0000_0000_0000_0000;
array[55236] <= 16'b0000_0000_0000_0000;
array[55237] <= 16'b0000_0000_0000_0000;
array[55238] <= 16'b0000_0000_0000_0000;
array[55239] <= 16'b0000_0000_0000_0000;
array[55240] <= 16'b0000_0000_0000_0000;
array[55241] <= 16'b0000_0000_0000_0000;
array[55242] <= 16'b0000_0000_0000_0000;
array[55243] <= 16'b0000_0000_0000_0000;
array[55244] <= 16'b0000_0000_0000_0000;
array[55245] <= 16'b0000_0000_0000_0000;
array[55246] <= 16'b0000_0000_0000_0000;
array[55247] <= 16'b0000_0000_0000_0000;
array[55248] <= 16'b0000_0000_0000_0000;
array[55249] <= 16'b0000_0000_0000_0000;
array[55250] <= 16'b0000_0000_0000_0000;
array[55251] <= 16'b0000_0000_0000_0000;
array[55252] <= 16'b0000_0000_0000_0000;
array[55253] <= 16'b0000_0000_0000_0000;
array[55254] <= 16'b0000_0000_0000_0000;
array[55255] <= 16'b0000_0000_0000_0000;
array[55256] <= 16'b0000_0000_0000_0000;
array[55257] <= 16'b0000_0000_0000_0000;
array[55258] <= 16'b0000_0000_0000_0000;
array[55259] <= 16'b0000_0000_0000_0000;
array[55260] <= 16'b0000_0000_0000_0000;
array[55261] <= 16'b0000_0000_0000_0000;
array[55262] <= 16'b0000_0000_0000_0000;
array[55263] <= 16'b0000_0000_0000_0000;
array[55264] <= 16'b0000_0000_0000_0000;
array[55265] <= 16'b0000_0000_0000_0000;
array[55266] <= 16'b0000_0000_0000_0000;
array[55267] <= 16'b0000_0000_0000_0000;
array[55268] <= 16'b0000_0000_0000_0000;
array[55269] <= 16'b0000_0000_0000_0000;
array[55270] <= 16'b0000_0000_0000_0000;
array[55271] <= 16'b0000_0000_0000_0000;
array[55272] <= 16'b0000_0000_0000_0000;
array[55273] <= 16'b0000_0000_0000_0000;
array[55274] <= 16'b0000_0000_0000_0000;
array[55275] <= 16'b0000_0000_0000_0000;
array[55276] <= 16'b0000_0000_0000_0000;
array[55277] <= 16'b0000_0000_0000_0000;
array[55278] <= 16'b0000_0000_0000_0000;
array[55279] <= 16'b0000_0000_0000_0000;
array[55280] <= 16'b0000_0000_0000_0000;
array[55281] <= 16'b0000_0000_0000_0000;
array[55282] <= 16'b0000_0000_0000_0000;
array[55283] <= 16'b0000_0000_0000_0000;
array[55284] <= 16'b0000_0000_0000_0000;
array[55285] <= 16'b0000_0000_0000_0000;
array[55286] <= 16'b0000_0000_0000_0000;
array[55287] <= 16'b0000_0000_0000_0000;
array[55288] <= 16'b0000_0000_0000_0000;
array[55289] <= 16'b0000_0000_0000_0000;
array[55290] <= 16'b0000_0000_0000_0000;
array[55291] <= 16'b0000_0000_0000_0000;
array[55292] <= 16'b0000_0000_0000_0000;
array[55293] <= 16'b0000_0000_0000_0000;
array[55294] <= 16'b0000_0000_0000_0000;
array[55295] <= 16'b0000_0000_0000_0000;
array[55296] <= 16'b0000_0000_0000_0000;
array[55297] <= 16'b0000_0000_0000_0000;
array[55298] <= 16'b0000_0000_0000_0000;
array[55299] <= 16'b0000_0000_0000_0000;
array[55300] <= 16'b0000_0000_0000_0000;
array[55301] <= 16'b0000_0000_0000_0000;
array[55302] <= 16'b0000_0000_0000_0000;
array[55303] <= 16'b0000_0000_0000_0000;
array[55304] <= 16'b0000_0000_0000_0000;
array[55305] <= 16'b0000_0000_0000_0000;
array[55306] <= 16'b0000_0000_0000_0000;
array[55307] <= 16'b0000_0000_0000_0000;
array[55308] <= 16'b0000_0000_0000_0000;
array[55309] <= 16'b0000_0000_0000_0000;
array[55310] <= 16'b0000_0000_0000_0000;
array[55311] <= 16'b0000_0000_0000_0000;
array[55312] <= 16'b0000_0000_0000_0000;
array[55313] <= 16'b0000_0000_0000_0000;
array[55314] <= 16'b0000_0000_0000_0000;
array[55315] <= 16'b0000_0000_0000_0000;
array[55316] <= 16'b0000_0000_0000_0000;
array[55317] <= 16'b0000_0000_0000_0000;
array[55318] <= 16'b0000_0000_0000_0000;
array[55319] <= 16'b0000_0000_0000_0000;
array[55320] <= 16'b0000_0000_0000_0000;
array[55321] <= 16'b0000_0000_0000_0000;
array[55322] <= 16'b0000_0000_0000_0000;
array[55323] <= 16'b0000_0000_0000_0000;
array[55324] <= 16'b0000_0000_0000_0000;
array[55325] <= 16'b0000_0000_0000_0000;
array[55326] <= 16'b0000_0000_0000_0000;
array[55327] <= 16'b0000_0000_0000_0000;
array[55328] <= 16'b0000_0000_0000_0000;
array[55329] <= 16'b0000_0000_0000_0000;
array[55330] <= 16'b0000_0000_0000_0000;
array[55331] <= 16'b0000_0000_0000_0000;
array[55332] <= 16'b0000_0000_0000_0000;
array[55333] <= 16'b0000_0000_0000_0000;
array[55334] <= 16'b0000_0000_0000_0000;
array[55335] <= 16'b0000_0000_0000_0000;
array[55336] <= 16'b0000_0000_0000_0000;
array[55337] <= 16'b0000_0000_0000_0000;
array[55338] <= 16'b0000_0000_0000_0000;
array[55339] <= 16'b0000_0000_0000_0000;
array[55340] <= 16'b0000_0000_0000_0000;
array[55341] <= 16'b0000_0000_0000_0000;
array[55342] <= 16'b0000_0000_0000_0000;
array[55343] <= 16'b0000_0000_0000_0000;
array[55344] <= 16'b0000_0000_0000_0000;
array[55345] <= 16'b0000_0000_0000_0000;
array[55346] <= 16'b0000_0000_0000_0000;
array[55347] <= 16'b0000_0000_0000_0000;
array[55348] <= 16'b0000_0000_0000_0000;
array[55349] <= 16'b0000_0000_0000_0000;
array[55350] <= 16'b0000_0000_0000_0000;
array[55351] <= 16'b0000_0000_0000_0000;
array[55352] <= 16'b0000_0000_0000_0000;
array[55353] <= 16'b0000_0000_0000_0000;
array[55354] <= 16'b0000_0000_0000_0000;
array[55355] <= 16'b0000_0000_0000_0000;
array[55356] <= 16'b0000_0000_0000_0000;
array[55357] <= 16'b0000_0000_0000_0000;
array[55358] <= 16'b0000_0000_0000_0000;
array[55359] <= 16'b0000_0000_0000_0000;
array[55360] <= 16'b0000_0000_0000_0000;
array[55361] <= 16'b0000_0000_0000_0000;
array[55362] <= 16'b0000_0000_0000_0000;
array[55363] <= 16'b0000_0000_0000_0000;
array[55364] <= 16'b0000_0000_0000_0000;
array[55365] <= 16'b0000_0000_0000_0000;
array[55366] <= 16'b0000_0000_0000_0000;
array[55367] <= 16'b0000_0000_0000_0000;
array[55368] <= 16'b0000_0000_0000_0000;
array[55369] <= 16'b0000_0000_0000_0000;
array[55370] <= 16'b0000_0000_0000_0000;
array[55371] <= 16'b0000_0000_0000_0000;
array[55372] <= 16'b0000_0000_0000_0000;
array[55373] <= 16'b0000_0000_0000_0000;
array[55374] <= 16'b0000_0000_0000_0000;
array[55375] <= 16'b0000_0000_0000_0000;
array[55376] <= 16'b0000_0000_0000_0000;
array[55377] <= 16'b0000_0000_0000_0000;
array[55378] <= 16'b0000_0000_0000_0000;
array[55379] <= 16'b0000_0000_0000_0000;
array[55380] <= 16'b0000_0000_0000_0000;
array[55381] <= 16'b0000_0000_0000_0000;
array[55382] <= 16'b0000_0000_0000_0000;
array[55383] <= 16'b0000_0000_0000_0000;
array[55384] <= 16'b0000_0000_0000_0000;
array[55385] <= 16'b0000_0000_0000_0000;
array[55386] <= 16'b0000_0000_0000_0000;
array[55387] <= 16'b0000_0000_0000_0000;
array[55388] <= 16'b0000_0000_0000_0000;
array[55389] <= 16'b0000_0000_0000_0000;
array[55390] <= 16'b0000_0000_0000_0000;
array[55391] <= 16'b0000_0000_0000_0000;
array[55392] <= 16'b0000_0000_0000_0000;
array[55393] <= 16'b0000_0000_0000_0000;
array[55394] <= 16'b0000_0000_0000_0000;
array[55395] <= 16'b0000_0000_0000_0000;
array[55396] <= 16'b0000_0000_0000_0000;
array[55397] <= 16'b0000_0000_0000_0000;
array[55398] <= 16'b0000_0000_0000_0000;
array[55399] <= 16'b0000_0000_0000_0000;
array[55400] <= 16'b0000_0000_0000_0000;
array[55401] <= 16'b0000_0000_0000_0000;
array[55402] <= 16'b0000_0000_0000_0000;
array[55403] <= 16'b0000_0000_0000_0000;
array[55404] <= 16'b0000_0000_0000_0000;
array[55405] <= 16'b0000_0000_0000_0000;
array[55406] <= 16'b0000_0000_0000_0000;
array[55407] <= 16'b0000_0000_0000_0000;
array[55408] <= 16'b0000_0000_0000_0000;
array[55409] <= 16'b0000_0000_0000_0000;
array[55410] <= 16'b0000_0000_0000_0000;
array[55411] <= 16'b0000_0000_0000_0000;
array[55412] <= 16'b0000_0000_0000_0000;
array[55413] <= 16'b0000_0000_0000_0000;
array[55414] <= 16'b0000_0000_0000_0000;
array[55415] <= 16'b0000_0000_0000_0000;
array[55416] <= 16'b0000_0000_0000_0000;
array[55417] <= 16'b0000_0000_0000_0000;
array[55418] <= 16'b0000_0000_0000_0000;
array[55419] <= 16'b0000_0000_0000_0000;
array[55420] <= 16'b0000_0000_0000_0000;
array[55421] <= 16'b0000_0000_0000_0000;
array[55422] <= 16'b0000_0000_0000_0000;
array[55423] <= 16'b0000_0000_0000_0000;
array[55424] <= 16'b0000_0000_0000_0000;
array[55425] <= 16'b0000_0000_0000_0000;
array[55426] <= 16'b0000_0000_0000_0000;
array[55427] <= 16'b0000_0000_0000_0000;
array[55428] <= 16'b0000_0000_0000_0000;
array[55429] <= 16'b0000_0000_0000_0000;
array[55430] <= 16'b0000_0000_0000_0000;
array[55431] <= 16'b0000_0000_0000_0000;
array[55432] <= 16'b0000_0000_0000_0000;
array[55433] <= 16'b0000_0000_0000_0000;
array[55434] <= 16'b0000_0000_0000_0000;
array[55435] <= 16'b0000_0000_0000_0000;
array[55436] <= 16'b0000_0000_0000_0000;
array[55437] <= 16'b0000_0000_0000_0000;
array[55438] <= 16'b0000_0000_0000_0000;
array[55439] <= 16'b0000_0000_0000_0000;
array[55440] <= 16'b0000_0000_0000_0000;
array[55441] <= 16'b0000_0000_0000_0000;
array[55442] <= 16'b0000_0000_0000_0000;
array[55443] <= 16'b0000_0000_0000_0000;
array[55444] <= 16'b0000_0000_0000_0000;
array[55445] <= 16'b0000_0000_0000_0000;
array[55446] <= 16'b0000_0000_0000_0000;
array[55447] <= 16'b0000_0000_0000_0000;
array[55448] <= 16'b0000_0000_0000_0000;
array[55449] <= 16'b0000_0000_0000_0000;
array[55450] <= 16'b0000_0000_0000_0000;
array[55451] <= 16'b0000_0000_0000_0000;
array[55452] <= 16'b0000_0000_0000_0000;
array[55453] <= 16'b0000_0000_0000_0000;
array[55454] <= 16'b0000_0000_0000_0000;
array[55455] <= 16'b0000_0000_0000_0000;
array[55456] <= 16'b0000_0000_0000_0000;
array[55457] <= 16'b0000_0000_0000_0000;
array[55458] <= 16'b0000_0000_0000_0000;
array[55459] <= 16'b0000_0000_0000_0000;
array[55460] <= 16'b0000_0000_0000_0000;
array[55461] <= 16'b0000_0000_0000_0000;
array[55462] <= 16'b0000_0000_0000_0000;
array[55463] <= 16'b0000_0000_0000_0000;
array[55464] <= 16'b0000_0000_0000_0000;
array[55465] <= 16'b0000_0000_0000_0000;
array[55466] <= 16'b0000_0000_0000_0000;
array[55467] <= 16'b0000_0000_0000_0000;
array[55468] <= 16'b0000_0000_0000_0000;
array[55469] <= 16'b0000_0000_0000_0000;
array[55470] <= 16'b0000_0000_0000_0000;
array[55471] <= 16'b0000_0000_0000_0000;
array[55472] <= 16'b0000_0000_0000_0000;
array[55473] <= 16'b0000_0000_0000_0000;
array[55474] <= 16'b0000_0000_0000_0000;
array[55475] <= 16'b0000_0000_0000_0000;
array[55476] <= 16'b0000_0000_0000_0000;
array[55477] <= 16'b0000_0000_0000_0000;
array[55478] <= 16'b0000_0000_0000_0000;
array[55479] <= 16'b0000_0000_0000_0000;
array[55480] <= 16'b0000_0000_0000_0000;
array[55481] <= 16'b0000_0000_0000_0000;
array[55482] <= 16'b0000_0000_0000_0000;
array[55483] <= 16'b0000_0000_0000_0000;
array[55484] <= 16'b0000_0000_0000_0000;
array[55485] <= 16'b0000_0000_0000_0000;
array[55486] <= 16'b0000_0000_0000_0000;
array[55487] <= 16'b0000_0000_0000_0000;
array[55488] <= 16'b0000_0000_0000_0000;
array[55489] <= 16'b0000_0000_0000_0000;
array[55490] <= 16'b0000_0000_0000_0000;
array[55491] <= 16'b0000_0000_0000_0000;
array[55492] <= 16'b0000_0000_0000_0000;
array[55493] <= 16'b0000_0000_0000_0000;
array[55494] <= 16'b0000_0000_0000_0000;
array[55495] <= 16'b0000_0000_0000_0000;
array[55496] <= 16'b0000_0000_0000_0000;
array[55497] <= 16'b0000_0000_0000_0000;
array[55498] <= 16'b0000_0000_0000_0000;
array[55499] <= 16'b0000_0000_0000_0000;
array[55500] <= 16'b0000_0000_0000_0000;
array[55501] <= 16'b0000_0000_0000_0000;
array[55502] <= 16'b0000_0000_0000_0000;
array[55503] <= 16'b0000_0000_0000_0000;
array[55504] <= 16'b0000_0000_0000_0000;
array[55505] <= 16'b0000_0000_0000_0000;
array[55506] <= 16'b0000_0000_0000_0000;
array[55507] <= 16'b0000_0000_0000_0000;
array[55508] <= 16'b0000_0000_0000_0000;
array[55509] <= 16'b0000_0000_0000_0000;
array[55510] <= 16'b0000_0000_0000_0000;
array[55511] <= 16'b0000_0000_0000_0000;
array[55512] <= 16'b0000_0000_0000_0000;
array[55513] <= 16'b0000_0000_0000_0000;
array[55514] <= 16'b0000_0000_0000_0000;
array[55515] <= 16'b0000_0000_0000_0000;
array[55516] <= 16'b0000_0000_0000_0000;
array[55517] <= 16'b0000_0000_0000_0000;
array[55518] <= 16'b0000_0000_0000_0000;
array[55519] <= 16'b0000_0000_0000_0000;
array[55520] <= 16'b0000_0000_0000_0000;
array[55521] <= 16'b0000_0000_0000_0000;
array[55522] <= 16'b0000_0000_0000_0000;
array[55523] <= 16'b0000_0000_0000_0000;
array[55524] <= 16'b0000_0000_0000_0000;
array[55525] <= 16'b0000_0000_0000_0000;
array[55526] <= 16'b0000_0000_0000_0000;
array[55527] <= 16'b0000_0000_0000_0000;
array[55528] <= 16'b0000_0000_0000_0000;
array[55529] <= 16'b0000_0000_0000_0000;
array[55530] <= 16'b0000_0000_0000_0000;
array[55531] <= 16'b0000_0000_0000_0000;
array[55532] <= 16'b0000_0000_0000_0000;
array[55533] <= 16'b0000_0000_0000_0000;
array[55534] <= 16'b0000_0000_0000_0000;
array[55535] <= 16'b0000_0000_0000_0000;
array[55536] <= 16'b0000_0000_0000_0000;
array[55537] <= 16'b0000_0000_0000_0000;
array[55538] <= 16'b0000_0000_0000_0000;
array[55539] <= 16'b0000_0000_0000_0000;
array[55540] <= 16'b0000_0000_0000_0000;
array[55541] <= 16'b0000_0000_0000_0000;
array[55542] <= 16'b0000_0000_0000_0000;
array[55543] <= 16'b0000_0000_0000_0000;
array[55544] <= 16'b0000_0000_0000_0000;
array[55545] <= 16'b0000_0000_0000_0000;
array[55546] <= 16'b0000_0000_0000_0000;
array[55547] <= 16'b0000_0000_0000_0000;
array[55548] <= 16'b0000_0000_0000_0000;
array[55549] <= 16'b0000_0000_0000_0000;
array[55550] <= 16'b0000_0000_0000_0000;
array[55551] <= 16'b0000_0000_0000_0000;
array[55552] <= 16'b0000_0000_0000_0000;
array[55553] <= 16'b0000_0000_0000_0000;
array[55554] <= 16'b0000_0000_0000_0000;
array[55555] <= 16'b0000_0000_0000_0000;
array[55556] <= 16'b0000_0000_0000_0000;
array[55557] <= 16'b0000_0000_0000_0000;
array[55558] <= 16'b0000_0000_0000_0000;
array[55559] <= 16'b0000_0000_0000_0000;
array[55560] <= 16'b0000_0000_0000_0000;
array[55561] <= 16'b0000_0000_0000_0000;
array[55562] <= 16'b0000_0000_0000_0000;
array[55563] <= 16'b0000_0000_0000_0000;
array[55564] <= 16'b0000_0000_0000_0000;
array[55565] <= 16'b0000_0000_0000_0000;
array[55566] <= 16'b0000_0000_0000_0000;
array[55567] <= 16'b0000_0000_0000_0000;
array[55568] <= 16'b0000_0000_0000_0000;
array[55569] <= 16'b0000_0000_0000_0000;
array[55570] <= 16'b0000_0000_0000_0000;
array[55571] <= 16'b0000_0000_0000_0000;
array[55572] <= 16'b0000_0000_0000_0000;
array[55573] <= 16'b0000_0000_0000_0000;
array[55574] <= 16'b0000_0000_0000_0000;
array[55575] <= 16'b0000_0000_0000_0000;
array[55576] <= 16'b0000_0000_0000_0000;
array[55577] <= 16'b0000_0000_0000_0000;
array[55578] <= 16'b0000_0000_0000_0000;
array[55579] <= 16'b0000_0000_0000_0000;
array[55580] <= 16'b0000_0000_0000_0000;
array[55581] <= 16'b0000_0000_0000_0000;
array[55582] <= 16'b0000_0000_0000_0000;
array[55583] <= 16'b0000_0000_0000_0000;
array[55584] <= 16'b0000_0000_0000_0000;
array[55585] <= 16'b0000_0000_0000_0000;
array[55586] <= 16'b0000_0000_0000_0000;
array[55587] <= 16'b0000_0000_0000_0000;
array[55588] <= 16'b0000_0000_0000_0000;
array[55589] <= 16'b0000_0000_0000_0000;
array[55590] <= 16'b0000_0000_0000_0000;
array[55591] <= 16'b0000_0000_0000_0000;
array[55592] <= 16'b0000_0000_0000_0000;
array[55593] <= 16'b0000_0000_0000_0000;
array[55594] <= 16'b0000_0000_0000_0000;
array[55595] <= 16'b0000_0000_0000_0000;
array[55596] <= 16'b0000_0000_0000_0000;
array[55597] <= 16'b0000_0000_0000_0000;
array[55598] <= 16'b0000_0000_0000_0000;
array[55599] <= 16'b0000_0000_0000_0000;
array[55600] <= 16'b0000_0000_0000_0000;
array[55601] <= 16'b0000_0000_0000_0000;
array[55602] <= 16'b0000_0000_0000_0000;
array[55603] <= 16'b0000_0000_0000_0000;
array[55604] <= 16'b0000_0000_0000_0000;
array[55605] <= 16'b0000_0000_0000_0000;
array[55606] <= 16'b0000_0000_0000_0000;
array[55607] <= 16'b0000_0000_0000_0000;
array[55608] <= 16'b0000_0000_0000_0000;
array[55609] <= 16'b0000_0000_0000_0000;
array[55610] <= 16'b0000_0000_0000_0000;
array[55611] <= 16'b0000_0000_0000_0000;
array[55612] <= 16'b0000_0000_0000_0000;
array[55613] <= 16'b0000_0000_0000_0000;
array[55614] <= 16'b0000_0000_0000_0000;
array[55615] <= 16'b0000_0000_0000_0000;
array[55616] <= 16'b0000_0000_0000_0000;
array[55617] <= 16'b0000_0000_0000_0000;
array[55618] <= 16'b0000_0000_0000_0000;
array[55619] <= 16'b0000_0000_0000_0000;
array[55620] <= 16'b0000_0000_0000_0000;
array[55621] <= 16'b0000_0000_0000_0000;
array[55622] <= 16'b0000_0000_0000_0000;
array[55623] <= 16'b0000_0000_0000_0000;
array[55624] <= 16'b0000_0000_0000_0000;
array[55625] <= 16'b0000_0000_0000_0000;
array[55626] <= 16'b0000_0000_0000_0000;
array[55627] <= 16'b0000_0000_0000_0000;
array[55628] <= 16'b0000_0000_0000_0000;
array[55629] <= 16'b0000_0000_0000_0000;
array[55630] <= 16'b0000_0000_0000_0000;
array[55631] <= 16'b0000_0000_0000_0000;
array[55632] <= 16'b0000_0000_0000_0000;
array[55633] <= 16'b0000_0000_0000_0000;
array[55634] <= 16'b0000_0000_0000_0000;
array[55635] <= 16'b0000_0000_0000_0000;
array[55636] <= 16'b0000_0000_0000_0000;
array[55637] <= 16'b0000_0000_0000_0000;
array[55638] <= 16'b0000_0000_0000_0000;
array[55639] <= 16'b0000_0000_0000_0000;
array[55640] <= 16'b0000_0000_0000_0000;
array[55641] <= 16'b0000_0000_0000_0000;
array[55642] <= 16'b0000_0000_0000_0000;
array[55643] <= 16'b0000_0000_0000_0000;
array[55644] <= 16'b0000_0000_0000_0000;
array[55645] <= 16'b0000_0000_0000_0000;
array[55646] <= 16'b0000_0000_0000_0000;
array[55647] <= 16'b0000_0000_0000_0000;
array[55648] <= 16'b0000_0000_0000_0000;
array[55649] <= 16'b0000_0000_0000_0000;
array[55650] <= 16'b0000_0000_0000_0000;
array[55651] <= 16'b0000_0000_0000_0000;
array[55652] <= 16'b0000_0000_0000_0000;
array[55653] <= 16'b0000_0000_0000_0000;
array[55654] <= 16'b0000_0000_0000_0000;
array[55655] <= 16'b0000_0000_0000_0000;
array[55656] <= 16'b0000_0000_0000_0000;
array[55657] <= 16'b0000_0000_0000_0000;
array[55658] <= 16'b0000_0000_0000_0000;
array[55659] <= 16'b0000_0000_0000_0000;
array[55660] <= 16'b0000_0000_0000_0000;
array[55661] <= 16'b0000_0000_0000_0000;
array[55662] <= 16'b0000_0000_0000_0000;
array[55663] <= 16'b0000_0000_0000_0000;
array[55664] <= 16'b0000_0000_0000_0000;
array[55665] <= 16'b0000_0000_0000_0000;
array[55666] <= 16'b0000_0000_0000_0000;
array[55667] <= 16'b0000_0000_0000_0000;
array[55668] <= 16'b0000_0000_0000_0000;
array[55669] <= 16'b0000_0000_0000_0000;
array[55670] <= 16'b0000_0000_0000_0000;
array[55671] <= 16'b0000_0000_0000_0000;
array[55672] <= 16'b0000_0000_0000_0000;
array[55673] <= 16'b0000_0000_0000_0000;
array[55674] <= 16'b0000_0000_0000_0000;
array[55675] <= 16'b0000_0000_0000_0000;
array[55676] <= 16'b0000_0000_0000_0000;
array[55677] <= 16'b0000_0000_0000_0000;
array[55678] <= 16'b0000_0000_0000_0000;
array[55679] <= 16'b0000_0000_0000_0000;
array[55680] <= 16'b0000_0000_0000_0000;
array[55681] <= 16'b0000_0000_0000_0000;
array[55682] <= 16'b0000_0000_0000_0000;
array[55683] <= 16'b0000_0000_0000_0000;
array[55684] <= 16'b0000_0000_0000_0000;
array[55685] <= 16'b0000_0000_0000_0000;
array[55686] <= 16'b0000_0000_0000_0000;
array[55687] <= 16'b0000_0000_0000_0000;
array[55688] <= 16'b0000_0000_0000_0000;
array[55689] <= 16'b0000_0000_0000_0000;
array[55690] <= 16'b0000_0000_0000_0000;
array[55691] <= 16'b0000_0000_0000_0000;
array[55692] <= 16'b0000_0000_0000_0000;
array[55693] <= 16'b0000_0000_0000_0000;
array[55694] <= 16'b0000_0000_0000_0000;
array[55695] <= 16'b0000_0000_0000_0000;
array[55696] <= 16'b0000_0000_0000_0000;
array[55697] <= 16'b0000_0000_0000_0000;
array[55698] <= 16'b0000_0000_0000_0000;
array[55699] <= 16'b0000_0000_0000_0000;
array[55700] <= 16'b0000_0000_0000_0000;
array[55701] <= 16'b0000_0000_0000_0000;
array[55702] <= 16'b0000_0000_0000_0000;
array[55703] <= 16'b0000_0000_0000_0000;
array[55704] <= 16'b0000_0000_0000_0000;
array[55705] <= 16'b0000_0000_0000_0000;
array[55706] <= 16'b0000_0000_0000_0000;
array[55707] <= 16'b0000_0000_0000_0000;
array[55708] <= 16'b0000_0000_0000_0000;
array[55709] <= 16'b0000_0000_0000_0000;
array[55710] <= 16'b0000_0000_0000_0000;
array[55711] <= 16'b0000_0000_0000_0000;
array[55712] <= 16'b0000_0000_0000_0000;
array[55713] <= 16'b0000_0000_0000_0000;
array[55714] <= 16'b0000_0000_0000_0000;
array[55715] <= 16'b0000_0000_0000_0000;
array[55716] <= 16'b0000_0000_0000_0000;
array[55717] <= 16'b0000_0000_0000_0000;
array[55718] <= 16'b0000_0000_0000_0000;
array[55719] <= 16'b0000_0000_0000_0000;
array[55720] <= 16'b0000_0000_0000_0000;
array[55721] <= 16'b0000_0000_0000_0000;
array[55722] <= 16'b0000_0000_0000_0000;
array[55723] <= 16'b0000_0000_0000_0000;
array[55724] <= 16'b0000_0000_0000_0000;
array[55725] <= 16'b0000_0000_0000_0000;
array[55726] <= 16'b0000_0000_0000_0000;
array[55727] <= 16'b0000_0000_0000_0000;
array[55728] <= 16'b0000_0000_0000_0000;
array[55729] <= 16'b0000_0000_0000_0000;
array[55730] <= 16'b0000_0000_0000_0000;
array[55731] <= 16'b0000_0000_0000_0000;
array[55732] <= 16'b0000_0000_0000_0000;
array[55733] <= 16'b0000_0000_0000_0000;
array[55734] <= 16'b0000_0000_0000_0000;
array[55735] <= 16'b0000_0000_0000_0000;
array[55736] <= 16'b0000_0000_0000_0000;
array[55737] <= 16'b0000_0000_0000_0000;
array[55738] <= 16'b0000_0000_0000_0000;
array[55739] <= 16'b0000_0000_0000_0000;
array[55740] <= 16'b0000_0000_0000_0000;
array[55741] <= 16'b0000_0000_0000_0000;
array[55742] <= 16'b0000_0000_0000_0000;
array[55743] <= 16'b0000_0000_0000_0000;
array[55744] <= 16'b0000_0000_0000_0000;
array[55745] <= 16'b0000_0000_0000_0000;
array[55746] <= 16'b0000_0000_0000_0000;
array[55747] <= 16'b0000_0000_0000_0000;
array[55748] <= 16'b0000_0000_0000_0000;
array[55749] <= 16'b0000_0000_0000_0000;
array[55750] <= 16'b0000_0000_0000_0000;
array[55751] <= 16'b0000_0000_0000_0000;
array[55752] <= 16'b0000_0000_0000_0000;
array[55753] <= 16'b0000_0000_0000_0000;
array[55754] <= 16'b0000_0000_0000_0000;
array[55755] <= 16'b0000_0000_0000_0000;
array[55756] <= 16'b0000_0000_0000_0000;
array[55757] <= 16'b0000_0000_0000_0000;
array[55758] <= 16'b0000_0000_0000_0000;
array[55759] <= 16'b0000_0000_0000_0000;
array[55760] <= 16'b0000_0000_0000_0000;
array[55761] <= 16'b0000_0000_0000_0000;
array[55762] <= 16'b0000_0000_0000_0000;
array[55763] <= 16'b0000_0000_0000_0000;
array[55764] <= 16'b0000_0000_0000_0000;
array[55765] <= 16'b0000_0000_0000_0000;
array[55766] <= 16'b0000_0000_0000_0000;
array[55767] <= 16'b0000_0000_0000_0000;
array[55768] <= 16'b0000_0000_0000_0000;
array[55769] <= 16'b0000_0000_0000_0000;
array[55770] <= 16'b0000_0000_0000_0000;
array[55771] <= 16'b0000_0000_0000_0000;
array[55772] <= 16'b0000_0000_0000_0000;
array[55773] <= 16'b0000_0000_0000_0000;
array[55774] <= 16'b0000_0000_0000_0000;
array[55775] <= 16'b0000_0000_0000_0000;
array[55776] <= 16'b0000_0000_0000_0000;
array[55777] <= 16'b0000_0000_0000_0000;
array[55778] <= 16'b0000_0000_0000_0000;
array[55779] <= 16'b0000_0000_0000_0000;
array[55780] <= 16'b0000_0000_0000_0000;
array[55781] <= 16'b0000_0000_0000_0000;
array[55782] <= 16'b0000_0000_0000_0000;
array[55783] <= 16'b0000_0000_0000_0000;
array[55784] <= 16'b0000_0000_0000_0000;
array[55785] <= 16'b0000_0000_0000_0000;
array[55786] <= 16'b0000_0000_0000_0000;
array[55787] <= 16'b0000_0000_0000_0000;
array[55788] <= 16'b0000_0000_0000_0000;
array[55789] <= 16'b0000_0000_0000_0000;
array[55790] <= 16'b0000_0000_0000_0000;
array[55791] <= 16'b0000_0000_0000_0000;
array[55792] <= 16'b0000_0000_0000_0000;
array[55793] <= 16'b0000_0000_0000_0000;
array[55794] <= 16'b0000_0000_0000_0000;
array[55795] <= 16'b0000_0000_0000_0000;
array[55796] <= 16'b0000_0000_0000_0000;
array[55797] <= 16'b0000_0000_0000_0000;
array[55798] <= 16'b0000_0000_0000_0000;
array[55799] <= 16'b0000_0000_0000_0000;
array[55800] <= 16'b0000_0000_0000_0000;
array[55801] <= 16'b0000_0000_0000_0000;
array[55802] <= 16'b0000_0000_0000_0000;
array[55803] <= 16'b0000_0000_0000_0000;
array[55804] <= 16'b0000_0000_0000_0000;
array[55805] <= 16'b0000_0000_0000_0000;
array[55806] <= 16'b0000_0000_0000_0000;
array[55807] <= 16'b0000_0000_0000_0000;
array[55808] <= 16'b0000_0000_0000_0000;
array[55809] <= 16'b0000_0000_0000_0000;
array[55810] <= 16'b0000_0000_0000_0000;
array[55811] <= 16'b0000_0000_0000_0000;
array[55812] <= 16'b0000_0000_0000_0000;
array[55813] <= 16'b0000_0000_0000_0000;
array[55814] <= 16'b0000_0000_0000_0000;
array[55815] <= 16'b0000_0000_0000_0000;
array[55816] <= 16'b0000_0000_0000_0000;
array[55817] <= 16'b0000_0000_0000_0000;
array[55818] <= 16'b0000_0000_0000_0000;
array[55819] <= 16'b0000_0000_0000_0000;
array[55820] <= 16'b0000_0000_0000_0000;
array[55821] <= 16'b0000_0000_0000_0000;
array[55822] <= 16'b0000_0000_0000_0000;
array[55823] <= 16'b0000_0000_0000_0000;
array[55824] <= 16'b0000_0000_0000_0000;
array[55825] <= 16'b0000_0000_0000_0000;
array[55826] <= 16'b0000_0000_0000_0000;
array[55827] <= 16'b0000_0000_0000_0000;
array[55828] <= 16'b0000_0000_0000_0000;
array[55829] <= 16'b0000_0000_0000_0000;
array[55830] <= 16'b0000_0000_0000_0000;
array[55831] <= 16'b0000_0000_0000_0000;
array[55832] <= 16'b0000_0000_0000_0000;
array[55833] <= 16'b0000_0000_0000_0000;
array[55834] <= 16'b0000_0000_0000_0000;
array[55835] <= 16'b0000_0000_0000_0000;
array[55836] <= 16'b0000_0000_0000_0000;
array[55837] <= 16'b0000_0000_0000_0000;
array[55838] <= 16'b0000_0000_0000_0000;
array[55839] <= 16'b0000_0000_0000_0000;
array[55840] <= 16'b0000_0000_0000_0000;
array[55841] <= 16'b0000_0000_0000_0000;
array[55842] <= 16'b0000_0000_0000_0000;
array[55843] <= 16'b0000_0000_0000_0000;
array[55844] <= 16'b0000_0000_0000_0000;
array[55845] <= 16'b0000_0000_0000_0000;
array[55846] <= 16'b0000_0000_0000_0000;
array[55847] <= 16'b0000_0000_0000_0000;
array[55848] <= 16'b0000_0000_0000_0000;
array[55849] <= 16'b0000_0000_0000_0000;
array[55850] <= 16'b0000_0000_0000_0000;
array[55851] <= 16'b0000_0000_0000_0000;
array[55852] <= 16'b0000_0000_0000_0000;
array[55853] <= 16'b0000_0000_0000_0000;
array[55854] <= 16'b0000_0000_0000_0000;
array[55855] <= 16'b0000_0000_0000_0000;
array[55856] <= 16'b0000_0000_0000_0000;
array[55857] <= 16'b0000_0000_0000_0000;
array[55858] <= 16'b0000_0000_0000_0000;
array[55859] <= 16'b0000_0000_0000_0000;
array[55860] <= 16'b0000_0000_0000_0000;
array[55861] <= 16'b0000_0000_0000_0000;
array[55862] <= 16'b0000_0000_0000_0000;
array[55863] <= 16'b0000_0000_0000_0000;
array[55864] <= 16'b0000_0000_0000_0000;
array[55865] <= 16'b0000_0000_0000_0000;
array[55866] <= 16'b0000_0000_0000_0000;
array[55867] <= 16'b0000_0000_0000_0000;
array[55868] <= 16'b0000_0000_0000_0000;
array[55869] <= 16'b0000_0000_0000_0000;
array[55870] <= 16'b0000_0000_0000_0000;
array[55871] <= 16'b0000_0000_0000_0000;
array[55872] <= 16'b0000_0000_0000_0000;
array[55873] <= 16'b0000_0000_0000_0000;
array[55874] <= 16'b0000_0000_0000_0000;
array[55875] <= 16'b0000_0000_0000_0000;
array[55876] <= 16'b0000_0000_0000_0000;
array[55877] <= 16'b0000_0000_0000_0000;
array[55878] <= 16'b0000_0000_0000_0000;
array[55879] <= 16'b0000_0000_0000_0000;
array[55880] <= 16'b0000_0000_0000_0000;
array[55881] <= 16'b0000_0000_0000_0000;
array[55882] <= 16'b0000_0000_0000_0000;
array[55883] <= 16'b0000_0000_0000_0000;
array[55884] <= 16'b0000_0000_0000_0000;
array[55885] <= 16'b0000_0000_0000_0000;
array[55886] <= 16'b0000_0000_0000_0000;
array[55887] <= 16'b0000_0000_0000_0000;
array[55888] <= 16'b0000_0000_0000_0000;
array[55889] <= 16'b0000_0000_0000_0000;
array[55890] <= 16'b0000_0000_0000_0000;
array[55891] <= 16'b0000_0000_0000_0000;
array[55892] <= 16'b0000_0000_0000_0000;
array[55893] <= 16'b0000_0000_0000_0000;
array[55894] <= 16'b0000_0000_0000_0000;
array[55895] <= 16'b0000_0000_0000_0000;
array[55896] <= 16'b0000_0000_0000_0000;
array[55897] <= 16'b0000_0000_0000_0000;
array[55898] <= 16'b0000_0000_0000_0000;
array[55899] <= 16'b0000_0000_0000_0000;
array[55900] <= 16'b0000_0000_0000_0000;
array[55901] <= 16'b0000_0000_0000_0000;
array[55902] <= 16'b0000_0000_0000_0000;
array[55903] <= 16'b0000_0000_0000_0000;
array[55904] <= 16'b0000_0000_0000_0000;
array[55905] <= 16'b0000_0000_0000_0000;
array[55906] <= 16'b0000_0000_0000_0000;
array[55907] <= 16'b0000_0000_0000_0000;
array[55908] <= 16'b0000_0000_0000_0000;
array[55909] <= 16'b0000_0000_0000_0000;
array[55910] <= 16'b0000_0000_0000_0000;
array[55911] <= 16'b0000_0000_0000_0000;
array[55912] <= 16'b0000_0000_0000_0000;
array[55913] <= 16'b0000_0000_0000_0000;
array[55914] <= 16'b0000_0000_0000_0000;
array[55915] <= 16'b0000_0000_0000_0000;
array[55916] <= 16'b0000_0000_0000_0000;
array[55917] <= 16'b0000_0000_0000_0000;
array[55918] <= 16'b0000_0000_0000_0000;
array[55919] <= 16'b0000_0000_0000_0000;
array[55920] <= 16'b0000_0000_0000_0000;
array[55921] <= 16'b0000_0000_0000_0000;
array[55922] <= 16'b0000_0000_0000_0000;
array[55923] <= 16'b0000_0000_0000_0000;
array[55924] <= 16'b0000_0000_0000_0000;
array[55925] <= 16'b0000_0000_0000_0000;
array[55926] <= 16'b0000_0000_0000_0000;
array[55927] <= 16'b0000_0000_0000_0000;
array[55928] <= 16'b0000_0000_0000_0000;
array[55929] <= 16'b0000_0000_0000_0000;
array[55930] <= 16'b0000_0000_0000_0000;
array[55931] <= 16'b0000_0000_0000_0000;
array[55932] <= 16'b0000_0000_0000_0000;
array[55933] <= 16'b0000_0000_0000_0000;
array[55934] <= 16'b0000_0000_0000_0000;
array[55935] <= 16'b0000_0000_0000_0000;
array[55936] <= 16'b0000_0000_0000_0000;
array[55937] <= 16'b0000_0000_0000_0000;
array[55938] <= 16'b0000_0000_0000_0000;
array[55939] <= 16'b0000_0000_0000_0000;
array[55940] <= 16'b0000_0000_0000_0000;
array[55941] <= 16'b0000_0000_0000_0000;
array[55942] <= 16'b0000_0000_0000_0000;
array[55943] <= 16'b0000_0000_0000_0000;
array[55944] <= 16'b0000_0000_0000_0000;
array[55945] <= 16'b0000_0000_0000_0000;
array[55946] <= 16'b0000_0000_0000_0000;
array[55947] <= 16'b0000_0000_0000_0000;
array[55948] <= 16'b0000_0000_0000_0000;
array[55949] <= 16'b0000_0000_0000_0000;
array[55950] <= 16'b0000_0000_0000_0000;
array[55951] <= 16'b0000_0000_0000_0000;
array[55952] <= 16'b0000_0000_0000_0000;
array[55953] <= 16'b0000_0000_0000_0000;
array[55954] <= 16'b0000_0000_0000_0000;
array[55955] <= 16'b0000_0000_0000_0000;
array[55956] <= 16'b0000_0000_0000_0000;
array[55957] <= 16'b0000_0000_0000_0000;
array[55958] <= 16'b0000_0000_0000_0000;
array[55959] <= 16'b0000_0000_0000_0000;
array[55960] <= 16'b0000_0000_0000_0000;
array[55961] <= 16'b0000_0000_0000_0000;
array[55962] <= 16'b0000_0000_0000_0000;
array[55963] <= 16'b0000_0000_0000_0000;
array[55964] <= 16'b0000_0000_0000_0000;
array[55965] <= 16'b0000_0000_0000_0000;
array[55966] <= 16'b0000_0000_0000_0000;
array[55967] <= 16'b0000_0000_0000_0000;
array[55968] <= 16'b0000_0000_0000_0000;
array[55969] <= 16'b0000_0000_0000_0000;
array[55970] <= 16'b0000_0000_0000_0000;
array[55971] <= 16'b0000_0000_0000_0000;
array[55972] <= 16'b0000_0000_0000_0000;
array[55973] <= 16'b0000_0000_0000_0000;
array[55974] <= 16'b0000_0000_0000_0000;
array[55975] <= 16'b0000_0000_0000_0000;
array[55976] <= 16'b0000_0000_0000_0000;
array[55977] <= 16'b0000_0000_0000_0000;
array[55978] <= 16'b0000_0000_0000_0000;
array[55979] <= 16'b0000_0000_0000_0000;
array[55980] <= 16'b0000_0000_0000_0000;
array[55981] <= 16'b0000_0000_0000_0000;
array[55982] <= 16'b0000_0000_0000_0000;
array[55983] <= 16'b0000_0000_0000_0000;
array[55984] <= 16'b0000_0000_0000_0000;
array[55985] <= 16'b0000_0000_0000_0000;
array[55986] <= 16'b0000_0000_0000_0000;
array[55987] <= 16'b0000_0000_0000_0000;
array[55988] <= 16'b0000_0000_0000_0000;
array[55989] <= 16'b0000_0000_0000_0000;
array[55990] <= 16'b0000_0000_0000_0000;
array[55991] <= 16'b0000_0000_0000_0000;
array[55992] <= 16'b0000_0000_0000_0000;
array[55993] <= 16'b0000_0000_0000_0000;
array[55994] <= 16'b0000_0000_0000_0000;
array[55995] <= 16'b0000_0000_0000_0000;
array[55996] <= 16'b0000_0000_0000_0000;
array[55997] <= 16'b0000_0000_0000_0000;
array[55998] <= 16'b0000_0000_0000_0000;
array[55999] <= 16'b0000_0000_0000_0000;
array[56000] <= 16'b0000_0000_0000_0000;
array[56001] <= 16'b0000_0000_0000_0000;
array[56002] <= 16'b0000_0000_0000_0000;
array[56003] <= 16'b0000_0000_0000_0000;
array[56004] <= 16'b0000_0000_0000_0000;
array[56005] <= 16'b0000_0000_0000_0000;
array[56006] <= 16'b0000_0000_0000_0000;
array[56007] <= 16'b0000_0000_0000_0000;
array[56008] <= 16'b0000_0000_0000_0000;
array[56009] <= 16'b0000_0000_0000_0000;
array[56010] <= 16'b0000_0000_0000_0000;
array[56011] <= 16'b0000_0000_0000_0000;
array[56012] <= 16'b0000_0000_0000_0000;
array[56013] <= 16'b0000_0000_0000_0000;
array[56014] <= 16'b0000_0000_0000_0000;
array[56015] <= 16'b0000_0000_0000_0000;
array[56016] <= 16'b0000_0000_0000_0000;
array[56017] <= 16'b0000_0000_0000_0000;
array[56018] <= 16'b0000_0000_0000_0000;
array[56019] <= 16'b0000_0000_0000_0000;
array[56020] <= 16'b0000_0000_0000_0000;
array[56021] <= 16'b0000_0000_0000_0000;
array[56022] <= 16'b0000_0000_0000_0000;
array[56023] <= 16'b0000_0000_0000_0000;
array[56024] <= 16'b0000_0000_0000_0000;
array[56025] <= 16'b0000_0000_0000_0000;
array[56026] <= 16'b0000_0000_0000_0000;
array[56027] <= 16'b0000_0000_0000_0000;
array[56028] <= 16'b0000_0000_0000_0000;
array[56029] <= 16'b0000_0000_0000_0000;
array[56030] <= 16'b0000_0000_0000_0000;
array[56031] <= 16'b0000_0000_0000_0000;
array[56032] <= 16'b0000_0000_0000_0000;
array[56033] <= 16'b0000_0000_0000_0000;
array[56034] <= 16'b0000_0000_0000_0000;
array[56035] <= 16'b0000_0000_0000_0000;
array[56036] <= 16'b0000_0000_0000_0000;
array[56037] <= 16'b0000_0000_0000_0000;
array[56038] <= 16'b0000_0000_0000_0000;
array[56039] <= 16'b0000_0000_0000_0000;
array[56040] <= 16'b0000_0000_0000_0000;
array[56041] <= 16'b0000_0000_0000_0000;
array[56042] <= 16'b0000_0000_0000_0000;
array[56043] <= 16'b0000_0000_0000_0000;
array[56044] <= 16'b0000_0000_0000_0000;
array[56045] <= 16'b0000_0000_0000_0000;
array[56046] <= 16'b0000_0000_0000_0000;
array[56047] <= 16'b0000_0000_0000_0000;
array[56048] <= 16'b0000_0000_0000_0000;
array[56049] <= 16'b0000_0000_0000_0000;
array[56050] <= 16'b0000_0000_0000_0000;
array[56051] <= 16'b0000_0000_0000_0000;
array[56052] <= 16'b0000_0000_0000_0000;
array[56053] <= 16'b0000_0000_0000_0000;
array[56054] <= 16'b0000_0000_0000_0000;
array[56055] <= 16'b0000_0000_0000_0000;
array[56056] <= 16'b0000_0000_0000_0000;
array[56057] <= 16'b0000_0000_0000_0000;
array[56058] <= 16'b0000_0000_0000_0000;
array[56059] <= 16'b0000_0000_0000_0000;
array[56060] <= 16'b0000_0000_0000_0000;
array[56061] <= 16'b0000_0000_0000_0000;
array[56062] <= 16'b0000_0000_0000_0000;
array[56063] <= 16'b0000_0000_0000_0000;
array[56064] <= 16'b0000_0000_0000_0000;
array[56065] <= 16'b0000_0000_0000_0000;
array[56066] <= 16'b0000_0000_0000_0000;
array[56067] <= 16'b0000_0000_0000_0000;
array[56068] <= 16'b0000_0000_0000_0000;
array[56069] <= 16'b0000_0000_0000_0000;
array[56070] <= 16'b0000_0000_0000_0000;
array[56071] <= 16'b0000_0000_0000_0000;
array[56072] <= 16'b0000_0000_0000_0000;
array[56073] <= 16'b0000_0000_0000_0000;
array[56074] <= 16'b0000_0000_0000_0000;
array[56075] <= 16'b0000_0000_0000_0000;
array[56076] <= 16'b0000_0000_0000_0000;
array[56077] <= 16'b0000_0000_0000_0000;
array[56078] <= 16'b0000_0000_0000_0000;
array[56079] <= 16'b0000_0000_0000_0000;
array[56080] <= 16'b0000_0000_0000_0000;
array[56081] <= 16'b0000_0000_0000_0000;
array[56082] <= 16'b0000_0000_0000_0000;
array[56083] <= 16'b0000_0000_0000_0000;
array[56084] <= 16'b0000_0000_0000_0000;
array[56085] <= 16'b0000_0000_0000_0000;
array[56086] <= 16'b0000_0000_0000_0000;
array[56087] <= 16'b0000_0000_0000_0000;
array[56088] <= 16'b0000_0000_0000_0000;
array[56089] <= 16'b0000_0000_0000_0000;
array[56090] <= 16'b0000_0000_0000_0000;
array[56091] <= 16'b0000_0000_0000_0000;
array[56092] <= 16'b0000_0000_0000_0000;
array[56093] <= 16'b0000_0000_0000_0000;
array[56094] <= 16'b0000_0000_0000_0000;
array[56095] <= 16'b0000_0000_0000_0000;
array[56096] <= 16'b0000_0000_0000_0000;
array[56097] <= 16'b0000_0000_0000_0000;
array[56098] <= 16'b0000_0000_0000_0000;
array[56099] <= 16'b0000_0000_0000_0000;
array[56100] <= 16'b0000_0000_0000_0000;
array[56101] <= 16'b0000_0000_0000_0000;
array[56102] <= 16'b0000_0000_0000_0000;
array[56103] <= 16'b0000_0000_0000_0000;
array[56104] <= 16'b0000_0000_0000_0000;
array[56105] <= 16'b0000_0000_0000_0000;
array[56106] <= 16'b0000_0000_0000_0000;
array[56107] <= 16'b0000_0000_0000_0000;
array[56108] <= 16'b0000_0000_0000_0000;
array[56109] <= 16'b0000_0000_0000_0000;
array[56110] <= 16'b0000_0000_0000_0000;
array[56111] <= 16'b0000_0000_0000_0000;
array[56112] <= 16'b0000_0000_0000_0000;
array[56113] <= 16'b0000_0000_0000_0000;
array[56114] <= 16'b0000_0000_0000_0000;
array[56115] <= 16'b0000_0000_0000_0000;
array[56116] <= 16'b0000_0000_0000_0000;
array[56117] <= 16'b0000_0000_0000_0000;
array[56118] <= 16'b0000_0000_0000_0000;
array[56119] <= 16'b0000_0000_0000_0000;
array[56120] <= 16'b0000_0000_0000_0000;
array[56121] <= 16'b0000_0000_0000_0000;
array[56122] <= 16'b0000_0000_0000_0000;
array[56123] <= 16'b0000_0000_0000_0000;
array[56124] <= 16'b0000_0000_0000_0000;
array[56125] <= 16'b0000_0000_0000_0000;
array[56126] <= 16'b0000_0000_0000_0000;
array[56127] <= 16'b0000_0000_0000_0000;
array[56128] <= 16'b0000_0000_0000_0000;
array[56129] <= 16'b0000_0000_0000_0000;
array[56130] <= 16'b0000_0000_0000_0000;
array[56131] <= 16'b0000_0000_0000_0000;
array[56132] <= 16'b0000_0000_0000_0000;
array[56133] <= 16'b0000_0000_0000_0000;
array[56134] <= 16'b0000_0000_0000_0000;
array[56135] <= 16'b0000_0000_0000_0000;
array[56136] <= 16'b0000_0000_0000_0000;
array[56137] <= 16'b0000_0000_0000_0000;
array[56138] <= 16'b0000_0000_0000_0000;
array[56139] <= 16'b0000_0000_0000_0000;
array[56140] <= 16'b0000_0000_0000_0000;
array[56141] <= 16'b0000_0000_0000_0000;
array[56142] <= 16'b0000_0000_0000_0000;
array[56143] <= 16'b0000_0000_0000_0000;
array[56144] <= 16'b0000_0000_0000_0000;
array[56145] <= 16'b0000_0000_0000_0000;
array[56146] <= 16'b0000_0000_0000_0000;
array[56147] <= 16'b0000_0000_0000_0000;
array[56148] <= 16'b0000_0000_0000_0000;
array[56149] <= 16'b0000_0000_0000_0000;
array[56150] <= 16'b0000_0000_0000_0000;
array[56151] <= 16'b0000_0000_0000_0000;
array[56152] <= 16'b0000_0000_0000_0000;
array[56153] <= 16'b0000_0000_0000_0000;
array[56154] <= 16'b0000_0000_0000_0000;
array[56155] <= 16'b0000_0000_0000_0000;
array[56156] <= 16'b0000_0000_0000_0000;
array[56157] <= 16'b0000_0000_0000_0000;
array[56158] <= 16'b0000_0000_0000_0000;
array[56159] <= 16'b0000_0000_0000_0000;
array[56160] <= 16'b0000_0000_0000_0000;
array[56161] <= 16'b0000_0000_0000_0000;
array[56162] <= 16'b0000_0000_0000_0000;
array[56163] <= 16'b0000_0000_0000_0000;
array[56164] <= 16'b0000_0000_0000_0000;
array[56165] <= 16'b0000_0000_0000_0000;
array[56166] <= 16'b0000_0000_0000_0000;
array[56167] <= 16'b0000_0000_0000_0000;
array[56168] <= 16'b0000_0000_0000_0000;
array[56169] <= 16'b0000_0000_0000_0000;
array[56170] <= 16'b0000_0000_0000_0000;
array[56171] <= 16'b0000_0000_0000_0000;
array[56172] <= 16'b0000_0000_0000_0000;
array[56173] <= 16'b0000_0000_0000_0000;
array[56174] <= 16'b0000_0000_0000_0000;
array[56175] <= 16'b0000_0000_0000_0000;
array[56176] <= 16'b0000_0000_0000_0000;
array[56177] <= 16'b0000_0000_0000_0000;
array[56178] <= 16'b0000_0000_0000_0000;
array[56179] <= 16'b0000_0000_0000_0000;
array[56180] <= 16'b0000_0000_0000_0000;
array[56181] <= 16'b0000_0000_0000_0000;
array[56182] <= 16'b0000_0000_0000_0000;
array[56183] <= 16'b0000_0000_0000_0000;
array[56184] <= 16'b0000_0000_0000_0000;
array[56185] <= 16'b0000_0000_0000_0000;
array[56186] <= 16'b0000_0000_0000_0000;
array[56187] <= 16'b0000_0000_0000_0000;
array[56188] <= 16'b0000_0000_0000_0000;
array[56189] <= 16'b0000_0000_0000_0000;
array[56190] <= 16'b0000_0000_0000_0000;
array[56191] <= 16'b0000_0000_0000_0000;
array[56192] <= 16'b0000_0000_0000_0000;
array[56193] <= 16'b0000_0000_0000_0000;
array[56194] <= 16'b0000_0000_0000_0000;
array[56195] <= 16'b0000_0000_0000_0000;
array[56196] <= 16'b0000_0000_0000_0000;
array[56197] <= 16'b0000_0000_0000_0000;
array[56198] <= 16'b0000_0000_0000_0000;
array[56199] <= 16'b0000_0000_0000_0000;
array[56200] <= 16'b0000_0000_0000_0000;
array[56201] <= 16'b0000_0000_0000_0000;
array[56202] <= 16'b0000_0000_0000_0000;
array[56203] <= 16'b0000_0000_0000_0000;
array[56204] <= 16'b0000_0000_0000_0000;
array[56205] <= 16'b0000_0000_0000_0000;
array[56206] <= 16'b0000_0000_0000_0000;
array[56207] <= 16'b0000_0000_0000_0000;
array[56208] <= 16'b0000_0000_0000_0000;
array[56209] <= 16'b0000_0000_0000_0000;
array[56210] <= 16'b0000_0000_0000_0000;
array[56211] <= 16'b0000_0000_0000_0000;
array[56212] <= 16'b0000_0000_0000_0000;
array[56213] <= 16'b0000_0000_0000_0000;
array[56214] <= 16'b0000_0000_0000_0000;
array[56215] <= 16'b0000_0000_0000_0000;
array[56216] <= 16'b0000_0000_0000_0000;
array[56217] <= 16'b0000_0000_0000_0000;
array[56218] <= 16'b0000_0000_0000_0000;
array[56219] <= 16'b0000_0000_0000_0000;
array[56220] <= 16'b0000_0000_0000_0000;
array[56221] <= 16'b0000_0000_0000_0000;
array[56222] <= 16'b0000_0000_0000_0000;
array[56223] <= 16'b0000_0000_0000_0000;
array[56224] <= 16'b0000_0000_0000_0000;
array[56225] <= 16'b0000_0000_0000_0000;
array[56226] <= 16'b0000_0000_0000_0000;
array[56227] <= 16'b0000_0000_0000_0000;
array[56228] <= 16'b0000_0000_0000_0000;
array[56229] <= 16'b0000_0000_0000_0000;
array[56230] <= 16'b0000_0000_0000_0000;
array[56231] <= 16'b0000_0000_0000_0000;
array[56232] <= 16'b0000_0000_0000_0000;
array[56233] <= 16'b0000_0000_0000_0000;
array[56234] <= 16'b0000_0000_0000_0000;
array[56235] <= 16'b0000_0000_0000_0000;
array[56236] <= 16'b0000_0000_0000_0000;
array[56237] <= 16'b0000_0000_0000_0000;
array[56238] <= 16'b0000_0000_0000_0000;
array[56239] <= 16'b0000_0000_0000_0000;
array[56240] <= 16'b0000_0000_0000_0000;
array[56241] <= 16'b0000_0000_0000_0000;
array[56242] <= 16'b0000_0000_0000_0000;
array[56243] <= 16'b0000_0000_0000_0000;
array[56244] <= 16'b0000_0000_0000_0000;
array[56245] <= 16'b0000_0000_0000_0000;
array[56246] <= 16'b0000_0000_0000_0000;
array[56247] <= 16'b0000_0000_0000_0000;
array[56248] <= 16'b0000_0000_0000_0000;
array[56249] <= 16'b0000_0000_0000_0000;
array[56250] <= 16'b0000_0000_0000_0000;
array[56251] <= 16'b0000_0000_0000_0000;
array[56252] <= 16'b0000_0000_0000_0000;
array[56253] <= 16'b0000_0000_0000_0000;
array[56254] <= 16'b0000_0000_0000_0000;
array[56255] <= 16'b0000_0000_0000_0000;
array[56256] <= 16'b0000_0000_0000_0000;
array[56257] <= 16'b0000_0000_0000_0000;
array[56258] <= 16'b0000_0000_0000_0000;
array[56259] <= 16'b0000_0000_0000_0000;
array[56260] <= 16'b0000_0000_0000_0000;
array[56261] <= 16'b0000_0000_0000_0000;
array[56262] <= 16'b0000_0000_0000_0000;
array[56263] <= 16'b0000_0000_0000_0000;
array[56264] <= 16'b0000_0000_0000_0000;
array[56265] <= 16'b0000_0000_0000_0000;
array[56266] <= 16'b0000_0000_0000_0000;
array[56267] <= 16'b0000_0000_0000_0000;
array[56268] <= 16'b0000_0000_0000_0000;
array[56269] <= 16'b0000_0000_0000_0000;
array[56270] <= 16'b0000_0000_0000_0000;
array[56271] <= 16'b0000_0000_0000_0000;
array[56272] <= 16'b0000_0000_0000_0000;
array[56273] <= 16'b0000_0000_0000_0000;
array[56274] <= 16'b0000_0000_0000_0000;
array[56275] <= 16'b0000_0000_0000_0000;
array[56276] <= 16'b0000_0000_0000_0000;
array[56277] <= 16'b0000_0000_0000_0000;
array[56278] <= 16'b0000_0000_0000_0000;
array[56279] <= 16'b0000_0000_0000_0000;
array[56280] <= 16'b0000_0000_0000_0000;
array[56281] <= 16'b0000_0000_0000_0000;
array[56282] <= 16'b0000_0000_0000_0000;
array[56283] <= 16'b0000_0000_0000_0000;
array[56284] <= 16'b0000_0000_0000_0000;
array[56285] <= 16'b0000_0000_0000_0000;
array[56286] <= 16'b0000_0000_0000_0000;
array[56287] <= 16'b0000_0000_0000_0000;
array[56288] <= 16'b0000_0000_0000_0000;
array[56289] <= 16'b0000_0000_0000_0000;
array[56290] <= 16'b0000_0000_0000_0000;
array[56291] <= 16'b0000_0000_0000_0000;
array[56292] <= 16'b0000_0000_0000_0000;
array[56293] <= 16'b0000_0000_0000_0000;
array[56294] <= 16'b0000_0000_0000_0000;
array[56295] <= 16'b0000_0000_0000_0000;
array[56296] <= 16'b0000_0000_0000_0000;
array[56297] <= 16'b0000_0000_0000_0000;
array[56298] <= 16'b0000_0000_0000_0000;
array[56299] <= 16'b0000_0000_0000_0000;
array[56300] <= 16'b0000_0000_0000_0000;
array[56301] <= 16'b0000_0000_0000_0000;
array[56302] <= 16'b0000_0000_0000_0000;
array[56303] <= 16'b0000_0000_0000_0000;
array[56304] <= 16'b0000_0000_0000_0000;
array[56305] <= 16'b0000_0000_0000_0000;
array[56306] <= 16'b0000_0000_0000_0000;
array[56307] <= 16'b0000_0000_0000_0000;
array[56308] <= 16'b0000_0000_0000_0000;
array[56309] <= 16'b0000_0000_0000_0000;
array[56310] <= 16'b0000_0000_0000_0000;
array[56311] <= 16'b0000_0000_0000_0000;
array[56312] <= 16'b0000_0000_0000_0000;
array[56313] <= 16'b0000_0000_0000_0000;
array[56314] <= 16'b0000_0000_0000_0000;
array[56315] <= 16'b0000_0000_0000_0000;
array[56316] <= 16'b0000_0000_0000_0000;
array[56317] <= 16'b0000_0000_0000_0000;
array[56318] <= 16'b0000_0000_0000_0000;
array[56319] <= 16'b0000_0000_0000_0000;
array[56320] <= 16'b0000_0000_0000_0000;
array[56321] <= 16'b0000_0000_0000_0000;
array[56322] <= 16'b0000_0000_0000_0000;
array[56323] <= 16'b0000_0000_0000_0000;
array[56324] <= 16'b0000_0000_0000_0000;
array[56325] <= 16'b0000_0000_0000_0000;
array[56326] <= 16'b0000_0000_0000_0000;
array[56327] <= 16'b0000_0000_0000_0000;
array[56328] <= 16'b0000_0000_0000_0000;
array[56329] <= 16'b0000_0000_0000_0000;
array[56330] <= 16'b0000_0000_0000_0000;
array[56331] <= 16'b0000_0000_0000_0000;
array[56332] <= 16'b0000_0000_0000_0000;
array[56333] <= 16'b0000_0000_0000_0000;
array[56334] <= 16'b0000_0000_0000_0000;
array[56335] <= 16'b0000_0000_0000_0000;
array[56336] <= 16'b0000_0000_0000_0000;
array[56337] <= 16'b0000_0000_0000_0000;
array[56338] <= 16'b0000_0000_0000_0000;
array[56339] <= 16'b0000_0000_0000_0000;
array[56340] <= 16'b0000_0000_0000_0000;
array[56341] <= 16'b0000_0000_0000_0000;
array[56342] <= 16'b0000_0000_0000_0000;
array[56343] <= 16'b0000_0000_0000_0000;
array[56344] <= 16'b0000_0000_0000_0000;
array[56345] <= 16'b0000_0000_0000_0000;
array[56346] <= 16'b0000_0000_0000_0000;
array[56347] <= 16'b0000_0000_0000_0000;
array[56348] <= 16'b0000_0000_0000_0000;
array[56349] <= 16'b0000_0000_0000_0000;
array[56350] <= 16'b0000_0000_0000_0000;
array[56351] <= 16'b0000_0000_0000_0000;
array[56352] <= 16'b0000_0000_0000_0000;
array[56353] <= 16'b0000_0000_0000_0000;
array[56354] <= 16'b0000_0000_0000_0000;
array[56355] <= 16'b0000_0000_0000_0000;
array[56356] <= 16'b0000_0000_0000_0000;
array[56357] <= 16'b0000_0000_0000_0000;
array[56358] <= 16'b0000_0000_0000_0000;
array[56359] <= 16'b0000_0000_0000_0000;
array[56360] <= 16'b0000_0000_0000_0000;
array[56361] <= 16'b0000_0000_0000_0000;
array[56362] <= 16'b0000_0000_0000_0000;
array[56363] <= 16'b0000_0000_0000_0000;
array[56364] <= 16'b0000_0000_0000_0000;
array[56365] <= 16'b0000_0000_0000_0000;
array[56366] <= 16'b0000_0000_0000_0000;
array[56367] <= 16'b0000_0000_0000_0000;
array[56368] <= 16'b0000_0000_0000_0000;
array[56369] <= 16'b0000_0000_0000_0000;
array[56370] <= 16'b0000_0000_0000_0000;
array[56371] <= 16'b0000_0000_0000_0000;
array[56372] <= 16'b0000_0000_0000_0000;
array[56373] <= 16'b0000_0000_0000_0000;
array[56374] <= 16'b0000_0000_0000_0000;
array[56375] <= 16'b0000_0000_0000_0000;
array[56376] <= 16'b0000_0000_0000_0000;
array[56377] <= 16'b0000_0000_0000_0000;
array[56378] <= 16'b0000_0000_0000_0000;
array[56379] <= 16'b0000_0000_0000_0000;
array[56380] <= 16'b0000_0000_0000_0000;
array[56381] <= 16'b0000_0000_0000_0000;
array[56382] <= 16'b0000_0000_0000_0000;
array[56383] <= 16'b0000_0000_0000_0000;
array[56384] <= 16'b0000_0000_0000_0000;
array[56385] <= 16'b0000_0000_0000_0000;
array[56386] <= 16'b0000_0000_0000_0000;
array[56387] <= 16'b0000_0000_0000_0000;
array[56388] <= 16'b0000_0000_0000_0000;
array[56389] <= 16'b0000_0000_0000_0000;
array[56390] <= 16'b0000_0000_0000_0000;
array[56391] <= 16'b0000_0000_0000_0000;
array[56392] <= 16'b0000_0000_0000_0000;
array[56393] <= 16'b0000_0000_0000_0000;
array[56394] <= 16'b0000_0000_0000_0000;
array[56395] <= 16'b0000_0000_0000_0000;
array[56396] <= 16'b0000_0000_0000_0000;
array[56397] <= 16'b0000_0000_0000_0000;
array[56398] <= 16'b0000_0000_0000_0000;
array[56399] <= 16'b0000_0000_0000_0000;
array[56400] <= 16'b0000_0000_0000_0000;
array[56401] <= 16'b0000_0000_0000_0000;
array[56402] <= 16'b0000_0000_0000_0000;
array[56403] <= 16'b0000_0000_0000_0000;
array[56404] <= 16'b0000_0000_0000_0000;
array[56405] <= 16'b0000_0000_0000_0000;
array[56406] <= 16'b0000_0000_0000_0000;
array[56407] <= 16'b0000_0000_0000_0000;
array[56408] <= 16'b0000_0000_0000_0000;
array[56409] <= 16'b0000_0000_0000_0000;
array[56410] <= 16'b0000_0000_0000_0000;
array[56411] <= 16'b0000_0000_0000_0000;
array[56412] <= 16'b0000_0000_0000_0000;
array[56413] <= 16'b0000_0000_0000_0000;
array[56414] <= 16'b0000_0000_0000_0000;
array[56415] <= 16'b0000_0000_0000_0000;
array[56416] <= 16'b0000_0000_0000_0000;
array[56417] <= 16'b0000_0000_0000_0000;
array[56418] <= 16'b0000_0000_0000_0000;
array[56419] <= 16'b0000_0000_0000_0000;
array[56420] <= 16'b0000_0000_0000_0000;
array[56421] <= 16'b0000_0000_0000_0000;
array[56422] <= 16'b0000_0000_0000_0000;
array[56423] <= 16'b0000_0000_0000_0000;
array[56424] <= 16'b0000_0000_0000_0000;
array[56425] <= 16'b0000_0000_0000_0000;
array[56426] <= 16'b0000_0000_0000_0000;
array[56427] <= 16'b0000_0000_0000_0000;
array[56428] <= 16'b0000_0000_0000_0000;
array[56429] <= 16'b0000_0000_0000_0000;
array[56430] <= 16'b0000_0000_0000_0000;
array[56431] <= 16'b0000_0000_0000_0000;
array[56432] <= 16'b0000_0000_0000_0000;
array[56433] <= 16'b0000_0000_0000_0000;
array[56434] <= 16'b0000_0000_0000_0000;
array[56435] <= 16'b0000_0000_0000_0000;
array[56436] <= 16'b0000_0000_0000_0000;
array[56437] <= 16'b0000_0000_0000_0000;
array[56438] <= 16'b0000_0000_0000_0000;
array[56439] <= 16'b0000_0000_0000_0000;
array[56440] <= 16'b0000_0000_0000_0000;
array[56441] <= 16'b0000_0000_0000_0000;
array[56442] <= 16'b0000_0000_0000_0000;
array[56443] <= 16'b0000_0000_0000_0000;
array[56444] <= 16'b0000_0000_0000_0000;
array[56445] <= 16'b0000_0000_0000_0000;
array[56446] <= 16'b0000_0000_0000_0000;
array[56447] <= 16'b0000_0000_0000_0000;
array[56448] <= 16'b0000_0000_0000_0000;
array[56449] <= 16'b0000_0000_0000_0000;
array[56450] <= 16'b0000_0000_0000_0000;
array[56451] <= 16'b0000_0000_0000_0000;
array[56452] <= 16'b0000_0000_0000_0000;
array[56453] <= 16'b0000_0000_0000_0000;
array[56454] <= 16'b0000_0000_0000_0000;
array[56455] <= 16'b0000_0000_0000_0000;
array[56456] <= 16'b0000_0000_0000_0000;
array[56457] <= 16'b0000_0000_0000_0000;
array[56458] <= 16'b0000_0000_0000_0000;
array[56459] <= 16'b0000_0000_0000_0000;
array[56460] <= 16'b0000_0000_0000_0000;
array[56461] <= 16'b0000_0000_0000_0000;
array[56462] <= 16'b0000_0000_0000_0000;
array[56463] <= 16'b0000_0000_0000_0000;
array[56464] <= 16'b0000_0000_0000_0000;
array[56465] <= 16'b0000_0000_0000_0000;
array[56466] <= 16'b0000_0000_0000_0000;
array[56467] <= 16'b0000_0000_0000_0000;
array[56468] <= 16'b0000_0000_0000_0000;
array[56469] <= 16'b0000_0000_0000_0000;
array[56470] <= 16'b0000_0000_0000_0000;
array[56471] <= 16'b0000_0000_0000_0000;
array[56472] <= 16'b0000_0000_0000_0000;
array[56473] <= 16'b0000_0000_0000_0000;
array[56474] <= 16'b0000_0000_0000_0000;
array[56475] <= 16'b0000_0000_0000_0000;
array[56476] <= 16'b0000_0000_0000_0000;
array[56477] <= 16'b0000_0000_0000_0000;
array[56478] <= 16'b0000_0000_0000_0000;
array[56479] <= 16'b0000_0000_0000_0000;
array[56480] <= 16'b0000_0000_0000_0000;
array[56481] <= 16'b0000_0000_0000_0000;
array[56482] <= 16'b0000_0000_0000_0000;
array[56483] <= 16'b0000_0000_0000_0000;
array[56484] <= 16'b0000_0000_0000_0000;
array[56485] <= 16'b0000_0000_0000_0000;
array[56486] <= 16'b0000_0000_0000_0000;
array[56487] <= 16'b0000_0000_0000_0000;
array[56488] <= 16'b0000_0000_0000_0000;
array[56489] <= 16'b0000_0000_0000_0000;
array[56490] <= 16'b0000_0000_0000_0000;
array[56491] <= 16'b0000_0000_0000_0000;
array[56492] <= 16'b0000_0000_0000_0000;
array[56493] <= 16'b0000_0000_0000_0000;
array[56494] <= 16'b0000_0000_0000_0000;
array[56495] <= 16'b0000_0000_0000_0000;
array[56496] <= 16'b0000_0000_0000_0000;
array[56497] <= 16'b0000_0000_0000_0000;
array[56498] <= 16'b0000_0000_0000_0000;
array[56499] <= 16'b0000_0000_0000_0000;
array[56500] <= 16'b0000_0000_0000_0000;
array[56501] <= 16'b0000_0000_0000_0000;
array[56502] <= 16'b0000_0000_0000_0000;
array[56503] <= 16'b0000_0000_0000_0000;
array[56504] <= 16'b0000_0000_0000_0000;
array[56505] <= 16'b0000_0000_0000_0000;
array[56506] <= 16'b0000_0000_0000_0000;
array[56507] <= 16'b0000_0000_0000_0000;
array[56508] <= 16'b0000_0000_0000_0000;
array[56509] <= 16'b0000_0000_0000_0000;
array[56510] <= 16'b0000_0000_0000_0000;
array[56511] <= 16'b0000_0000_0000_0000;
array[56512] <= 16'b0000_0000_0000_0000;
array[56513] <= 16'b0000_0000_0000_0000;
array[56514] <= 16'b0000_0000_0000_0000;
array[56515] <= 16'b0000_0000_0000_0000;
array[56516] <= 16'b0000_0000_0000_0000;
array[56517] <= 16'b0000_0000_0000_0000;
array[56518] <= 16'b0000_0000_0000_0000;
array[56519] <= 16'b0000_0000_0000_0000;
array[56520] <= 16'b0000_0000_0000_0000;
array[56521] <= 16'b0000_0000_0000_0000;
array[56522] <= 16'b0000_0000_0000_0000;
array[56523] <= 16'b0000_0000_0000_0000;
array[56524] <= 16'b0000_0000_0000_0000;
array[56525] <= 16'b0000_0000_0000_0000;
array[56526] <= 16'b0000_0000_0000_0000;
array[56527] <= 16'b0000_0000_0000_0000;
array[56528] <= 16'b0000_0000_0000_0000;
array[56529] <= 16'b0000_0000_0000_0000;
array[56530] <= 16'b0000_0000_0000_0000;
array[56531] <= 16'b0000_0000_0000_0000;
array[56532] <= 16'b0000_0000_0000_0000;
array[56533] <= 16'b0000_0000_0000_0000;
array[56534] <= 16'b0000_0000_0000_0000;
array[56535] <= 16'b0000_0000_0000_0000;
array[56536] <= 16'b0000_0000_0000_0000;
array[56537] <= 16'b0000_0000_0000_0000;
array[56538] <= 16'b0000_0000_0000_0000;
array[56539] <= 16'b0000_0000_0000_0000;
array[56540] <= 16'b0000_0000_0000_0000;
array[56541] <= 16'b0000_0000_0000_0000;
array[56542] <= 16'b0000_0000_0000_0000;
array[56543] <= 16'b0000_0000_0000_0000;
array[56544] <= 16'b0000_0000_0000_0000;
array[56545] <= 16'b0000_0000_0000_0000;
array[56546] <= 16'b0000_0000_0000_0000;
array[56547] <= 16'b0000_0000_0000_0000;
array[56548] <= 16'b0000_0000_0000_0000;
array[56549] <= 16'b0000_0000_0000_0000;
array[56550] <= 16'b0000_0000_0000_0000;
array[56551] <= 16'b0000_0000_0000_0000;
array[56552] <= 16'b0000_0000_0000_0000;
array[56553] <= 16'b0000_0000_0000_0000;
array[56554] <= 16'b0000_0000_0000_0000;
array[56555] <= 16'b0000_0000_0000_0000;
array[56556] <= 16'b0000_0000_0000_0000;
array[56557] <= 16'b0000_0000_0000_0000;
array[56558] <= 16'b0000_0000_0000_0000;
array[56559] <= 16'b0000_0000_0000_0000;
array[56560] <= 16'b0000_0000_0000_0000;
array[56561] <= 16'b0000_0000_0000_0000;
array[56562] <= 16'b0000_0000_0000_0000;
array[56563] <= 16'b0000_0000_0000_0000;
array[56564] <= 16'b0000_0000_0000_0000;
array[56565] <= 16'b0000_0000_0000_0000;
array[56566] <= 16'b0000_0000_0000_0000;
array[56567] <= 16'b0000_0000_0000_0000;
array[56568] <= 16'b0000_0000_0000_0000;
array[56569] <= 16'b0000_0000_0000_0000;
array[56570] <= 16'b0000_0000_0000_0000;
array[56571] <= 16'b0000_0000_0000_0000;
array[56572] <= 16'b0000_0000_0000_0000;
array[56573] <= 16'b0000_0000_0000_0000;
array[56574] <= 16'b0000_0000_0000_0000;
array[56575] <= 16'b0000_0000_0000_0000;
array[56576] <= 16'b0000_0000_0000_0000;
array[56577] <= 16'b0000_0000_0000_0000;
array[56578] <= 16'b0000_0000_0000_0000;
array[56579] <= 16'b0000_0000_0000_0000;
array[56580] <= 16'b0000_0000_0000_0000;
array[56581] <= 16'b0000_0000_0000_0000;
array[56582] <= 16'b0000_0000_0000_0000;
array[56583] <= 16'b0000_0000_0000_0000;
array[56584] <= 16'b0000_0000_0000_0000;
array[56585] <= 16'b0000_0000_0000_0000;
array[56586] <= 16'b0000_0000_0000_0000;
array[56587] <= 16'b0000_0000_0000_0000;
array[56588] <= 16'b0000_0000_0000_0000;
array[56589] <= 16'b0000_0000_0000_0000;
array[56590] <= 16'b0000_0000_0000_0000;
array[56591] <= 16'b0000_0000_0000_0000;
array[56592] <= 16'b0000_0000_0000_0000;
array[56593] <= 16'b0000_0000_0000_0000;
array[56594] <= 16'b0000_0000_0000_0000;
array[56595] <= 16'b0000_0000_0000_0000;
array[56596] <= 16'b0000_0000_0000_0000;
array[56597] <= 16'b0000_0000_0000_0000;
array[56598] <= 16'b0000_0000_0000_0000;
array[56599] <= 16'b0000_0000_0000_0000;
array[56600] <= 16'b0000_0000_0000_0000;
array[56601] <= 16'b0000_0000_0000_0000;
array[56602] <= 16'b0000_0000_0000_0000;
array[56603] <= 16'b0000_0000_0000_0000;
array[56604] <= 16'b0000_0000_0000_0000;
array[56605] <= 16'b0000_0000_0000_0000;
array[56606] <= 16'b0000_0000_0000_0000;
array[56607] <= 16'b0000_0000_0000_0000;
array[56608] <= 16'b0000_0000_0000_0000;
array[56609] <= 16'b0000_0000_0000_0000;
array[56610] <= 16'b0000_0000_0000_0000;
array[56611] <= 16'b0000_0000_0000_0000;
array[56612] <= 16'b0000_0000_0000_0000;
array[56613] <= 16'b0000_0000_0000_0000;
array[56614] <= 16'b0000_0000_0000_0000;
array[56615] <= 16'b0000_0000_0000_0000;
array[56616] <= 16'b0000_0000_0000_0000;
array[56617] <= 16'b0000_0000_0000_0000;
array[56618] <= 16'b0000_0000_0000_0000;
array[56619] <= 16'b0000_0000_0000_0000;
array[56620] <= 16'b0000_0000_0000_0000;
array[56621] <= 16'b0000_0000_0000_0000;
array[56622] <= 16'b0000_0000_0000_0000;
array[56623] <= 16'b0000_0000_0000_0000;
array[56624] <= 16'b0000_0000_0000_0000;
array[56625] <= 16'b0000_0000_0000_0000;
array[56626] <= 16'b0000_0000_0000_0000;
array[56627] <= 16'b0000_0000_0000_0000;
array[56628] <= 16'b0000_0000_0000_0000;
array[56629] <= 16'b0000_0000_0000_0000;
array[56630] <= 16'b0000_0000_0000_0000;
array[56631] <= 16'b0000_0000_0000_0000;
array[56632] <= 16'b0000_0000_0000_0000;
array[56633] <= 16'b0000_0000_0000_0000;
array[56634] <= 16'b0000_0000_0000_0000;
array[56635] <= 16'b0000_0000_0000_0000;
array[56636] <= 16'b0000_0000_0000_0000;
array[56637] <= 16'b0000_0000_0000_0000;
array[56638] <= 16'b0000_0000_0000_0000;
array[56639] <= 16'b0000_0000_0000_0000;
array[56640] <= 16'b0000_0000_0000_0000;
array[56641] <= 16'b0000_0000_0000_0000;
array[56642] <= 16'b0000_0000_0000_0000;
array[56643] <= 16'b0000_0000_0000_0000;
array[56644] <= 16'b0000_0000_0000_0000;
array[56645] <= 16'b0000_0000_0000_0000;
array[56646] <= 16'b0000_0000_0000_0000;
array[56647] <= 16'b0000_0000_0000_0000;
array[56648] <= 16'b0000_0000_0000_0000;
array[56649] <= 16'b0000_0000_0000_0000;
array[56650] <= 16'b0000_0000_0000_0000;
array[56651] <= 16'b0000_0000_0000_0000;
array[56652] <= 16'b0000_0000_0000_0000;
array[56653] <= 16'b0000_0000_0000_0000;
array[56654] <= 16'b0000_0000_0000_0000;
array[56655] <= 16'b0000_0000_0000_0000;
array[56656] <= 16'b0000_0000_0000_0000;
array[56657] <= 16'b0000_0000_0000_0000;
array[56658] <= 16'b0000_0000_0000_0000;
array[56659] <= 16'b0000_0000_0000_0000;
array[56660] <= 16'b0000_0000_0000_0000;
array[56661] <= 16'b0000_0000_0000_0000;
array[56662] <= 16'b0000_0000_0000_0000;
array[56663] <= 16'b0000_0000_0000_0000;
array[56664] <= 16'b0000_0000_0000_0000;
array[56665] <= 16'b0000_0000_0000_0000;
array[56666] <= 16'b0000_0000_0000_0000;
array[56667] <= 16'b0000_0000_0000_0000;
array[56668] <= 16'b0000_0000_0000_0000;
array[56669] <= 16'b0000_0000_0000_0000;
array[56670] <= 16'b0000_0000_0000_0000;
array[56671] <= 16'b0000_0000_0000_0000;
array[56672] <= 16'b0000_0000_0000_0000;
array[56673] <= 16'b0000_0000_0000_0000;
array[56674] <= 16'b0000_0000_0000_0000;
array[56675] <= 16'b0000_0000_0000_0000;
array[56676] <= 16'b0000_0000_0000_0000;
array[56677] <= 16'b0000_0000_0000_0000;
array[56678] <= 16'b0000_0000_0000_0000;
array[56679] <= 16'b0000_0000_0000_0000;
array[56680] <= 16'b0000_0000_0000_0000;
array[56681] <= 16'b0000_0000_0000_0000;
array[56682] <= 16'b0000_0000_0000_0000;
array[56683] <= 16'b0000_0000_0000_0000;
array[56684] <= 16'b0000_0000_0000_0000;
array[56685] <= 16'b0000_0000_0000_0000;
array[56686] <= 16'b0000_0000_0000_0000;
array[56687] <= 16'b0000_0000_0000_0000;
array[56688] <= 16'b0000_0000_0000_0000;
array[56689] <= 16'b0000_0000_0000_0000;
array[56690] <= 16'b0000_0000_0000_0000;
array[56691] <= 16'b0000_0000_0000_0000;
array[56692] <= 16'b0000_0000_0000_0000;
array[56693] <= 16'b0000_0000_0000_0000;
array[56694] <= 16'b0000_0000_0000_0000;
array[56695] <= 16'b0000_0000_0000_0000;
array[56696] <= 16'b0000_0000_0000_0000;
array[56697] <= 16'b0000_0000_0000_0000;
array[56698] <= 16'b0000_0000_0000_0000;
array[56699] <= 16'b0000_0000_0000_0000;
array[56700] <= 16'b0000_0000_0000_0000;
array[56701] <= 16'b0000_0000_0000_0000;
array[56702] <= 16'b0000_0000_0000_0000;
array[56703] <= 16'b0000_0000_0000_0000;
array[56704] <= 16'b0000_0000_0000_0000;
array[56705] <= 16'b0000_0000_0000_0000;
array[56706] <= 16'b0000_0000_0000_0000;
array[56707] <= 16'b0000_0000_0000_0000;
array[56708] <= 16'b0000_0000_0000_0000;
array[56709] <= 16'b0000_0000_0000_0000;
array[56710] <= 16'b0000_0000_0000_0000;
array[56711] <= 16'b0000_0000_0000_0000;
array[56712] <= 16'b0000_0000_0000_0000;
array[56713] <= 16'b0000_0000_0000_0000;
array[56714] <= 16'b0000_0000_0000_0000;
array[56715] <= 16'b0000_0000_0000_0000;
array[56716] <= 16'b0000_0000_0000_0000;
array[56717] <= 16'b0000_0000_0000_0000;
array[56718] <= 16'b0000_0000_0000_0000;
array[56719] <= 16'b0000_0000_0000_0000;
array[56720] <= 16'b0000_0000_0000_0000;
array[56721] <= 16'b0000_0000_0000_0000;
array[56722] <= 16'b0000_0000_0000_0000;
array[56723] <= 16'b0000_0000_0000_0000;
array[56724] <= 16'b0000_0000_0000_0000;
array[56725] <= 16'b0000_0000_0000_0000;
array[56726] <= 16'b0000_0000_0000_0000;
array[56727] <= 16'b0000_0000_0000_0000;
array[56728] <= 16'b0000_0000_0000_0000;
array[56729] <= 16'b0000_0000_0000_0000;
array[56730] <= 16'b0000_0000_0000_0000;
array[56731] <= 16'b0000_0000_0000_0000;
array[56732] <= 16'b0000_0000_0000_0000;
array[56733] <= 16'b0000_0000_0000_0000;
array[56734] <= 16'b0000_0000_0000_0000;
array[56735] <= 16'b0000_0000_0000_0000;
array[56736] <= 16'b0000_0000_0000_0000;
array[56737] <= 16'b0000_0000_0000_0000;
array[56738] <= 16'b0000_0000_0000_0000;
array[56739] <= 16'b0000_0000_0000_0000;
array[56740] <= 16'b0000_0000_0000_0000;
array[56741] <= 16'b0000_0000_0000_0000;
array[56742] <= 16'b0000_0000_0000_0000;
array[56743] <= 16'b0000_0000_0000_0000;
array[56744] <= 16'b0000_0000_0000_0000;
array[56745] <= 16'b0000_0000_0000_0000;
array[56746] <= 16'b0000_0000_0000_0000;
array[56747] <= 16'b0000_0000_0000_0000;
array[56748] <= 16'b0000_0000_0000_0000;
array[56749] <= 16'b0000_0000_0000_0000;
array[56750] <= 16'b0000_0000_0000_0000;
array[56751] <= 16'b0000_0000_0000_0000;
array[56752] <= 16'b0000_0000_0000_0000;
array[56753] <= 16'b0000_0000_0000_0000;
array[56754] <= 16'b0000_0000_0000_0000;
array[56755] <= 16'b0000_0000_0000_0000;
array[56756] <= 16'b0000_0000_0000_0000;
array[56757] <= 16'b0000_0000_0000_0000;
array[56758] <= 16'b0000_0000_0000_0000;
array[56759] <= 16'b0000_0000_0000_0000;
array[56760] <= 16'b0000_0000_0000_0000;
array[56761] <= 16'b0000_0000_0000_0000;
array[56762] <= 16'b0000_0000_0000_0000;
array[56763] <= 16'b0000_0000_0000_0000;
array[56764] <= 16'b0000_0000_0000_0000;
array[56765] <= 16'b0000_0000_0000_0000;
array[56766] <= 16'b0000_0000_0000_0000;
array[56767] <= 16'b0000_0000_0000_0000;
array[56768] <= 16'b0000_0000_0000_0000;
array[56769] <= 16'b0000_0000_0000_0000;
array[56770] <= 16'b0000_0000_0000_0000;
array[56771] <= 16'b0000_0000_0000_0000;
array[56772] <= 16'b0000_0000_0000_0000;
array[56773] <= 16'b0000_0000_0000_0000;
array[56774] <= 16'b0000_0000_0000_0000;
array[56775] <= 16'b0000_0000_0000_0000;
array[56776] <= 16'b0000_0000_0000_0000;
array[56777] <= 16'b0000_0000_0000_0000;
array[56778] <= 16'b0000_0000_0000_0000;
array[56779] <= 16'b0000_0000_0000_0000;
array[56780] <= 16'b0000_0000_0000_0000;
array[56781] <= 16'b0000_0000_0000_0000;
array[56782] <= 16'b0000_0000_0000_0000;
array[56783] <= 16'b0000_0000_0000_0000;
array[56784] <= 16'b0000_0000_0000_0000;
array[56785] <= 16'b0000_0000_0000_0000;
array[56786] <= 16'b0000_0000_0000_0000;
array[56787] <= 16'b0000_0000_0000_0000;
array[56788] <= 16'b0000_0000_0000_0000;
array[56789] <= 16'b0000_0000_0000_0000;
array[56790] <= 16'b0000_0000_0000_0000;
array[56791] <= 16'b0000_0000_0000_0000;
array[56792] <= 16'b0000_0000_0000_0000;
array[56793] <= 16'b0000_0000_0000_0000;
array[56794] <= 16'b0000_0000_0000_0000;
array[56795] <= 16'b0000_0000_0000_0000;
array[56796] <= 16'b0000_0000_0000_0000;
array[56797] <= 16'b0000_0000_0000_0000;
array[56798] <= 16'b0000_0000_0000_0000;
array[56799] <= 16'b0000_0000_0000_0000;
array[56800] <= 16'b0000_0000_0000_0000;
array[56801] <= 16'b0000_0000_0000_0000;
array[56802] <= 16'b0000_0000_0000_0000;
array[56803] <= 16'b0000_0000_0000_0000;
array[56804] <= 16'b0000_0000_0000_0000;
array[56805] <= 16'b0000_0000_0000_0000;
array[56806] <= 16'b0000_0000_0000_0000;
array[56807] <= 16'b0000_0000_0000_0000;
array[56808] <= 16'b0000_0000_0000_0000;
array[56809] <= 16'b0000_0000_0000_0000;
array[56810] <= 16'b0000_0000_0000_0000;
array[56811] <= 16'b0000_0000_0000_0000;
array[56812] <= 16'b0000_0000_0000_0000;
array[56813] <= 16'b0000_0000_0000_0000;
array[56814] <= 16'b0000_0000_0000_0000;
array[56815] <= 16'b0000_0000_0000_0000;
array[56816] <= 16'b0000_0000_0000_0000;
array[56817] <= 16'b0000_0000_0000_0000;
array[56818] <= 16'b0000_0000_0000_0000;
array[56819] <= 16'b0000_0000_0000_0000;
array[56820] <= 16'b0000_0000_0000_0000;
array[56821] <= 16'b0000_0000_0000_0000;
array[56822] <= 16'b0000_0000_0000_0000;
array[56823] <= 16'b0000_0000_0000_0000;
array[56824] <= 16'b0000_0000_0000_0000;
array[56825] <= 16'b0000_0000_0000_0000;
array[56826] <= 16'b0000_0000_0000_0000;
array[56827] <= 16'b0000_0000_0000_0000;
array[56828] <= 16'b0000_0000_0000_0000;
array[56829] <= 16'b0000_0000_0000_0000;
array[56830] <= 16'b0000_0000_0000_0000;
array[56831] <= 16'b0000_0000_0000_0000;
array[56832] <= 16'b0000_0000_0000_0000;
array[56833] <= 16'b0000_0000_0000_0000;
array[56834] <= 16'b0000_0000_0000_0000;
array[56835] <= 16'b0000_0000_0000_0000;
array[56836] <= 16'b0000_0000_0000_0000;
array[56837] <= 16'b0000_0000_0000_0000;
array[56838] <= 16'b0000_0000_0000_0000;
array[56839] <= 16'b0000_0000_0000_0000;
array[56840] <= 16'b0000_0000_0000_0000;
array[56841] <= 16'b0000_0000_0000_0000;
array[56842] <= 16'b0000_0000_0000_0000;
array[56843] <= 16'b0000_0000_0000_0000;
array[56844] <= 16'b0000_0000_0000_0000;
array[56845] <= 16'b0000_0000_0000_0000;
array[56846] <= 16'b0000_0000_0000_0000;
array[56847] <= 16'b0000_0000_0000_0000;
array[56848] <= 16'b0000_0000_0000_0000;
array[56849] <= 16'b0000_0000_0000_0000;
array[56850] <= 16'b0000_0000_0000_0000;
array[56851] <= 16'b0000_0000_0000_0000;
array[56852] <= 16'b0000_0000_0000_0000;
array[56853] <= 16'b0000_0000_0000_0000;
array[56854] <= 16'b0000_0000_0000_0000;
array[56855] <= 16'b0000_0000_0000_0000;
array[56856] <= 16'b0000_0000_0000_0000;
array[56857] <= 16'b0000_0000_0000_0000;
array[56858] <= 16'b0000_0000_0000_0000;
array[56859] <= 16'b0000_0000_0000_0000;
array[56860] <= 16'b0000_0000_0000_0000;
array[56861] <= 16'b0000_0000_0000_0000;
array[56862] <= 16'b0000_0000_0000_0000;
array[56863] <= 16'b0000_0000_0000_0000;
array[56864] <= 16'b0000_0000_0000_0000;
array[56865] <= 16'b0000_0000_0000_0000;
array[56866] <= 16'b0000_0000_0000_0000;
array[56867] <= 16'b0000_0000_0000_0000;
array[56868] <= 16'b0000_0000_0000_0000;
array[56869] <= 16'b0000_0000_0000_0000;
array[56870] <= 16'b0000_0000_0000_0000;
array[56871] <= 16'b0000_0000_0000_0000;
array[56872] <= 16'b0000_0000_0000_0000;
array[56873] <= 16'b0000_0000_0000_0000;
array[56874] <= 16'b0000_0000_0000_0000;
array[56875] <= 16'b0000_0000_0000_0000;
array[56876] <= 16'b0000_0000_0000_0000;
array[56877] <= 16'b0000_0000_0000_0000;
array[56878] <= 16'b0000_0000_0000_0000;
array[56879] <= 16'b0000_0000_0000_0000;
array[56880] <= 16'b0000_0000_0000_0000;
array[56881] <= 16'b0000_0000_0000_0000;
array[56882] <= 16'b0000_0000_0000_0000;
array[56883] <= 16'b0000_0000_0000_0000;
array[56884] <= 16'b0000_0000_0000_0000;
array[56885] <= 16'b0000_0000_0000_0000;
array[56886] <= 16'b0000_0000_0000_0000;
array[56887] <= 16'b0000_0000_0000_0000;
array[56888] <= 16'b0000_0000_0000_0000;
array[56889] <= 16'b0000_0000_0000_0000;
array[56890] <= 16'b0000_0000_0000_0000;
array[56891] <= 16'b0000_0000_0000_0000;
array[56892] <= 16'b0000_0000_0000_0000;
array[56893] <= 16'b0000_0000_0000_0000;
array[56894] <= 16'b0000_0000_0000_0000;
array[56895] <= 16'b0000_0000_0000_0000;
array[56896] <= 16'b0000_0000_0000_0000;
array[56897] <= 16'b0000_0000_0000_0000;
array[56898] <= 16'b0000_0000_0000_0000;
array[56899] <= 16'b0000_0000_0000_0000;
array[56900] <= 16'b0000_0000_0000_0000;
array[56901] <= 16'b0000_0000_0000_0000;
array[56902] <= 16'b0000_0000_0000_0000;
array[56903] <= 16'b0000_0000_0000_0000;
array[56904] <= 16'b0000_0000_0000_0000;
array[56905] <= 16'b0000_0000_0000_0000;
array[56906] <= 16'b0000_0000_0000_0000;
array[56907] <= 16'b0000_0000_0000_0000;
array[56908] <= 16'b0000_0000_0000_0000;
array[56909] <= 16'b0000_0000_0000_0000;
array[56910] <= 16'b0000_0000_0000_0000;
array[56911] <= 16'b0000_0000_0000_0000;
array[56912] <= 16'b0000_0000_0000_0000;
array[56913] <= 16'b0000_0000_0000_0000;
array[56914] <= 16'b0000_0000_0000_0000;
array[56915] <= 16'b0000_0000_0000_0000;
array[56916] <= 16'b0000_0000_0000_0000;
array[56917] <= 16'b0000_0000_0000_0000;
array[56918] <= 16'b0000_0000_0000_0000;
array[56919] <= 16'b0000_0000_0000_0000;
array[56920] <= 16'b0000_0000_0000_0000;
array[56921] <= 16'b0000_0000_0000_0000;
array[56922] <= 16'b0000_0000_0000_0000;
array[56923] <= 16'b0000_0000_0000_0000;
array[56924] <= 16'b0000_0000_0000_0000;
array[56925] <= 16'b0000_0000_0000_0000;
array[56926] <= 16'b0000_0000_0000_0000;
array[56927] <= 16'b0000_0000_0000_0000;
array[56928] <= 16'b0000_0000_0000_0000;
array[56929] <= 16'b0000_0000_0000_0000;
array[56930] <= 16'b0000_0000_0000_0000;
array[56931] <= 16'b0000_0000_0000_0000;
array[56932] <= 16'b0000_0000_0000_0000;
array[56933] <= 16'b0000_0000_0000_0000;
array[56934] <= 16'b0000_0000_0000_0000;
array[56935] <= 16'b0000_0000_0000_0000;
array[56936] <= 16'b0000_0000_0000_0000;
array[56937] <= 16'b0000_0000_0000_0000;
array[56938] <= 16'b0000_0000_0000_0000;
array[56939] <= 16'b0000_0000_0000_0000;
array[56940] <= 16'b0000_0000_0000_0000;
array[56941] <= 16'b0000_0000_0000_0000;
array[56942] <= 16'b0000_0000_0000_0000;
array[56943] <= 16'b0000_0000_0000_0000;
array[56944] <= 16'b0000_0000_0000_0000;
array[56945] <= 16'b0000_0000_0000_0000;
array[56946] <= 16'b0000_0000_0000_0000;
array[56947] <= 16'b0000_0000_0000_0000;
array[56948] <= 16'b0000_0000_0000_0000;
array[56949] <= 16'b0000_0000_0000_0000;
array[56950] <= 16'b0000_0000_0000_0000;
array[56951] <= 16'b0000_0000_0000_0000;
array[56952] <= 16'b0000_0000_0000_0000;
array[56953] <= 16'b0000_0000_0000_0000;
array[56954] <= 16'b0000_0000_0000_0000;
array[56955] <= 16'b0000_0000_0000_0000;
array[56956] <= 16'b0000_0000_0000_0000;
array[56957] <= 16'b0000_0000_0000_0000;
array[56958] <= 16'b0000_0000_0000_0000;
array[56959] <= 16'b0000_0000_0000_0000;
array[56960] <= 16'b0000_0000_0000_0000;
array[56961] <= 16'b0000_0000_0000_0000;
array[56962] <= 16'b0000_0000_0000_0000;
array[56963] <= 16'b0000_0000_0000_0000;
array[56964] <= 16'b0000_0000_0000_0000;
array[56965] <= 16'b0000_0000_0000_0000;
array[56966] <= 16'b0000_0000_0000_0000;
array[56967] <= 16'b0000_0000_0000_0000;
array[56968] <= 16'b0000_0000_0000_0000;
array[56969] <= 16'b0000_0000_0000_0000;
array[56970] <= 16'b0000_0000_0000_0000;
array[56971] <= 16'b0000_0000_0000_0000;
array[56972] <= 16'b0000_0000_0000_0000;
array[56973] <= 16'b0000_0000_0000_0000;
array[56974] <= 16'b0000_0000_0000_0000;
array[56975] <= 16'b0000_0000_0000_0000;
array[56976] <= 16'b0000_0000_0000_0000;
array[56977] <= 16'b0000_0000_0000_0000;
array[56978] <= 16'b0000_0000_0000_0000;
array[56979] <= 16'b0000_0000_0000_0000;
array[56980] <= 16'b0000_0000_0000_0000;
array[56981] <= 16'b0000_0000_0000_0000;
array[56982] <= 16'b0000_0000_0000_0000;
array[56983] <= 16'b0000_0000_0000_0000;
array[56984] <= 16'b0000_0000_0000_0000;
array[56985] <= 16'b0000_0000_0000_0000;
array[56986] <= 16'b0000_0000_0000_0000;
array[56987] <= 16'b0000_0000_0000_0000;
array[56988] <= 16'b0000_0000_0000_0000;
array[56989] <= 16'b0000_0000_0000_0000;
array[56990] <= 16'b0000_0000_0000_0000;
array[56991] <= 16'b0000_0000_0000_0000;
array[56992] <= 16'b0000_0000_0000_0000;
array[56993] <= 16'b0000_0000_0000_0000;
array[56994] <= 16'b0000_0000_0000_0000;
array[56995] <= 16'b0000_0000_0000_0000;
array[56996] <= 16'b0000_0000_0000_0000;
array[56997] <= 16'b0000_0000_0000_0000;
array[56998] <= 16'b0000_0000_0000_0000;
array[56999] <= 16'b0000_0000_0000_0000;
array[57000] <= 16'b0000_0000_0000_0000;
array[57001] <= 16'b0000_0000_0000_0000;
array[57002] <= 16'b0000_0000_0000_0000;
array[57003] <= 16'b0000_0000_0000_0000;
array[57004] <= 16'b0000_0000_0000_0000;
array[57005] <= 16'b0000_0000_0000_0000;
array[57006] <= 16'b0000_0000_0000_0000;
array[57007] <= 16'b0000_0000_0000_0000;
array[57008] <= 16'b0000_0000_0000_0000;
array[57009] <= 16'b0000_0000_0000_0000;
array[57010] <= 16'b0000_0000_0000_0000;
array[57011] <= 16'b0000_0000_0000_0000;
array[57012] <= 16'b0000_0000_0000_0000;
array[57013] <= 16'b0000_0000_0000_0000;
array[57014] <= 16'b0000_0000_0000_0000;
array[57015] <= 16'b0000_0000_0000_0000;
array[57016] <= 16'b0000_0000_0000_0000;
array[57017] <= 16'b0000_0000_0000_0000;
array[57018] <= 16'b0000_0000_0000_0000;
array[57019] <= 16'b0000_0000_0000_0000;
array[57020] <= 16'b0000_0000_0000_0000;
array[57021] <= 16'b0000_0000_0000_0000;
array[57022] <= 16'b0000_0000_0000_0000;
array[57023] <= 16'b0000_0000_0000_0000;
array[57024] <= 16'b0000_0000_0000_0000;
array[57025] <= 16'b0000_0000_0000_0000;
array[57026] <= 16'b0000_0000_0000_0000;
array[57027] <= 16'b0000_0000_0000_0000;
array[57028] <= 16'b0000_0000_0000_0000;
array[57029] <= 16'b0000_0000_0000_0000;
array[57030] <= 16'b0000_0000_0000_0000;
array[57031] <= 16'b0000_0000_0000_0000;
array[57032] <= 16'b0000_0000_0000_0000;
array[57033] <= 16'b0000_0000_0000_0000;
array[57034] <= 16'b0000_0000_0000_0000;
array[57035] <= 16'b0000_0000_0000_0000;
array[57036] <= 16'b0000_0000_0000_0000;
array[57037] <= 16'b0000_0000_0000_0000;
array[57038] <= 16'b0000_0000_0000_0000;
array[57039] <= 16'b0000_0000_0000_0000;
array[57040] <= 16'b0000_0000_0000_0000;
array[57041] <= 16'b0000_0000_0000_0000;
array[57042] <= 16'b0000_0000_0000_0000;
array[57043] <= 16'b0000_0000_0000_0000;
array[57044] <= 16'b0000_0000_0000_0000;
array[57045] <= 16'b0000_0000_0000_0000;
array[57046] <= 16'b0000_0000_0000_0000;
array[57047] <= 16'b0000_0000_0000_0000;
array[57048] <= 16'b0000_0000_0000_0000;
array[57049] <= 16'b0000_0000_0000_0000;
array[57050] <= 16'b0000_0000_0000_0000;
array[57051] <= 16'b0000_0000_0000_0000;
array[57052] <= 16'b0000_0000_0000_0000;
array[57053] <= 16'b0000_0000_0000_0000;
array[57054] <= 16'b0000_0000_0000_0000;
array[57055] <= 16'b0000_0000_0000_0000;
array[57056] <= 16'b0000_0000_0000_0000;
array[57057] <= 16'b0000_0000_0000_0000;
array[57058] <= 16'b0000_0000_0000_0000;
array[57059] <= 16'b0000_0000_0000_0000;
array[57060] <= 16'b0000_0000_0000_0000;
array[57061] <= 16'b0000_0000_0000_0000;
array[57062] <= 16'b0000_0000_0000_0000;
array[57063] <= 16'b0000_0000_0000_0000;
array[57064] <= 16'b0000_0000_0000_0000;
array[57065] <= 16'b0000_0000_0000_0000;
array[57066] <= 16'b0000_0000_0000_0000;
array[57067] <= 16'b0000_0000_0000_0000;
array[57068] <= 16'b0000_0000_0000_0000;
array[57069] <= 16'b0000_0000_0000_0000;
array[57070] <= 16'b0000_0000_0000_0000;
array[57071] <= 16'b0000_0000_0000_0000;
array[57072] <= 16'b0000_0000_0000_0000;
array[57073] <= 16'b0000_0000_0000_0000;
array[57074] <= 16'b0000_0000_0000_0000;
array[57075] <= 16'b0000_0000_0000_0000;
array[57076] <= 16'b0000_0000_0000_0000;
array[57077] <= 16'b0000_0000_0000_0000;
array[57078] <= 16'b0000_0000_0000_0000;
array[57079] <= 16'b0000_0000_0000_0000;
array[57080] <= 16'b0000_0000_0000_0000;
array[57081] <= 16'b0000_0000_0000_0000;
array[57082] <= 16'b0000_0000_0000_0000;
array[57083] <= 16'b0000_0000_0000_0000;
array[57084] <= 16'b0000_0000_0000_0000;
array[57085] <= 16'b0000_0000_0000_0000;
array[57086] <= 16'b0000_0000_0000_0000;
array[57087] <= 16'b0000_0000_0000_0000;
array[57088] <= 16'b0000_0000_0000_0000;
array[57089] <= 16'b0000_0000_0000_0000;
array[57090] <= 16'b0000_0000_0000_0000;
array[57091] <= 16'b0000_0000_0000_0000;
array[57092] <= 16'b0000_0000_0000_0000;
array[57093] <= 16'b0000_0000_0000_0000;
array[57094] <= 16'b0000_0000_0000_0000;
array[57095] <= 16'b0000_0000_0000_0000;
array[57096] <= 16'b0000_0000_0000_0000;
array[57097] <= 16'b0000_0000_0000_0000;
array[57098] <= 16'b0000_0000_0000_0000;
array[57099] <= 16'b0000_0000_0000_0000;
array[57100] <= 16'b0000_0000_0000_0000;
array[57101] <= 16'b0000_0000_0000_0000;
array[57102] <= 16'b0000_0000_0000_0000;
array[57103] <= 16'b0000_0000_0000_0000;
array[57104] <= 16'b0000_0000_0000_0000;
array[57105] <= 16'b0000_0000_0000_0000;
array[57106] <= 16'b0000_0000_0000_0000;
array[57107] <= 16'b0000_0000_0000_0000;
array[57108] <= 16'b0000_0000_0000_0000;
array[57109] <= 16'b0000_0000_0000_0000;
array[57110] <= 16'b0000_0000_0000_0000;
array[57111] <= 16'b0000_0000_0000_0000;
array[57112] <= 16'b0000_0000_0000_0000;
array[57113] <= 16'b0000_0000_0000_0000;
array[57114] <= 16'b0000_0000_0000_0000;
array[57115] <= 16'b0000_0000_0000_0000;
array[57116] <= 16'b0000_0000_0000_0000;
array[57117] <= 16'b0000_0000_0000_0000;
array[57118] <= 16'b0000_0000_0000_0000;
array[57119] <= 16'b0000_0000_0000_0000;
array[57120] <= 16'b0000_0000_0000_0000;
array[57121] <= 16'b0000_0000_0000_0000;
array[57122] <= 16'b0000_0000_0000_0000;
array[57123] <= 16'b0000_0000_0000_0000;
array[57124] <= 16'b0000_0000_0000_0000;
array[57125] <= 16'b0000_0000_0000_0000;
array[57126] <= 16'b0000_0000_0000_0000;
array[57127] <= 16'b0000_0000_0000_0000;
array[57128] <= 16'b0000_0000_0000_0000;
array[57129] <= 16'b0000_0000_0000_0000;
array[57130] <= 16'b0000_0000_0000_0000;
array[57131] <= 16'b0000_0000_0000_0000;
array[57132] <= 16'b0000_0000_0000_0000;
array[57133] <= 16'b0000_0000_0000_0000;
array[57134] <= 16'b0000_0000_0000_0000;
array[57135] <= 16'b0000_0000_0000_0000;
array[57136] <= 16'b0000_0000_0000_0000;
array[57137] <= 16'b0000_0000_0000_0000;
array[57138] <= 16'b0000_0000_0000_0000;
array[57139] <= 16'b0000_0000_0000_0000;
array[57140] <= 16'b0000_0000_0000_0000;
array[57141] <= 16'b0000_0000_0000_0000;
array[57142] <= 16'b0000_0000_0000_0000;
array[57143] <= 16'b0000_0000_0000_0000;
array[57144] <= 16'b0000_0000_0000_0000;
array[57145] <= 16'b0000_0000_0000_0000;
array[57146] <= 16'b0000_0000_0000_0000;
array[57147] <= 16'b0000_0000_0000_0000;
array[57148] <= 16'b0000_0000_0000_0000;
array[57149] <= 16'b0000_0000_0000_0000;
array[57150] <= 16'b0000_0000_0000_0000;
array[57151] <= 16'b0000_0000_0000_0000;
array[57152] <= 16'b0000_0000_0000_0000;
array[57153] <= 16'b0000_0000_0000_0000;
array[57154] <= 16'b0000_0000_0000_0000;
array[57155] <= 16'b0000_0000_0000_0000;
array[57156] <= 16'b0000_0000_0000_0000;
array[57157] <= 16'b0000_0000_0000_0000;
array[57158] <= 16'b0000_0000_0000_0000;
array[57159] <= 16'b0000_0000_0000_0000;
array[57160] <= 16'b0000_0000_0000_0000;
array[57161] <= 16'b0000_0000_0000_0000;
array[57162] <= 16'b0000_0000_0000_0000;
array[57163] <= 16'b0000_0000_0000_0000;
array[57164] <= 16'b0000_0000_0000_0000;
array[57165] <= 16'b0000_0000_0000_0000;
array[57166] <= 16'b0000_0000_0000_0000;
array[57167] <= 16'b0000_0000_0000_0000;
array[57168] <= 16'b0000_0000_0000_0000;
array[57169] <= 16'b0000_0000_0000_0000;
array[57170] <= 16'b0000_0000_0000_0000;
array[57171] <= 16'b0000_0000_0000_0000;
array[57172] <= 16'b0000_0000_0000_0000;
array[57173] <= 16'b0000_0000_0000_0000;
array[57174] <= 16'b0000_0000_0000_0000;
array[57175] <= 16'b0000_0000_0000_0000;
array[57176] <= 16'b0000_0000_0000_0000;
array[57177] <= 16'b0000_0000_0000_0000;
array[57178] <= 16'b0000_0000_0000_0000;
array[57179] <= 16'b0000_0000_0000_0000;
array[57180] <= 16'b0000_0000_0000_0000;
array[57181] <= 16'b0000_0000_0000_0000;
array[57182] <= 16'b0000_0000_0000_0000;
array[57183] <= 16'b0000_0000_0000_0000;
array[57184] <= 16'b0000_0000_0000_0000;
array[57185] <= 16'b0000_0000_0000_0000;
array[57186] <= 16'b0000_0000_0000_0000;
array[57187] <= 16'b0000_0000_0000_0000;
array[57188] <= 16'b0000_0000_0000_0000;
array[57189] <= 16'b0000_0000_0000_0000;
array[57190] <= 16'b0000_0000_0000_0000;
array[57191] <= 16'b0000_0000_0000_0000;
array[57192] <= 16'b0000_0000_0000_0000;
array[57193] <= 16'b0000_0000_0000_0000;
array[57194] <= 16'b0000_0000_0000_0000;
array[57195] <= 16'b0000_0000_0000_0000;
array[57196] <= 16'b0000_0000_0000_0000;
array[57197] <= 16'b0000_0000_0000_0000;
array[57198] <= 16'b0000_0000_0000_0000;
array[57199] <= 16'b0000_0000_0000_0000;
array[57200] <= 16'b0000_0000_0000_0000;
array[57201] <= 16'b0000_0000_0000_0000;
array[57202] <= 16'b0000_0000_0000_0000;
array[57203] <= 16'b0000_0000_0000_0000;
array[57204] <= 16'b0000_0000_0000_0000;
array[57205] <= 16'b0000_0000_0000_0000;
array[57206] <= 16'b0000_0000_0000_0000;
array[57207] <= 16'b0000_0000_0000_0000;
array[57208] <= 16'b0000_0000_0000_0000;
array[57209] <= 16'b0000_0000_0000_0000;
array[57210] <= 16'b0000_0000_0000_0000;
array[57211] <= 16'b0000_0000_0000_0000;
array[57212] <= 16'b0000_0000_0000_0000;
array[57213] <= 16'b0000_0000_0000_0000;
array[57214] <= 16'b0000_0000_0000_0000;
array[57215] <= 16'b0000_0000_0000_0000;
array[57216] <= 16'b0000_0000_0000_0000;
array[57217] <= 16'b0000_0000_0000_0000;
array[57218] <= 16'b0000_0000_0000_0000;
array[57219] <= 16'b0000_0000_0000_0000;
array[57220] <= 16'b0000_0000_0000_0000;
array[57221] <= 16'b0000_0000_0000_0000;
array[57222] <= 16'b0000_0000_0000_0000;
array[57223] <= 16'b0000_0000_0000_0000;
array[57224] <= 16'b0000_0000_0000_0000;
array[57225] <= 16'b0000_0000_0000_0000;
array[57226] <= 16'b0000_0000_0000_0000;
array[57227] <= 16'b0000_0000_0000_0000;
array[57228] <= 16'b0000_0000_0000_0000;
array[57229] <= 16'b0000_0000_0000_0000;
array[57230] <= 16'b0000_0000_0000_0000;
array[57231] <= 16'b0000_0000_0000_0000;
array[57232] <= 16'b0000_0000_0000_0000;
array[57233] <= 16'b0000_0000_0000_0000;
array[57234] <= 16'b0000_0000_0000_0000;
array[57235] <= 16'b0000_0000_0000_0000;
array[57236] <= 16'b0000_0000_0000_0000;
array[57237] <= 16'b0000_0000_0000_0000;
array[57238] <= 16'b0000_0000_0000_0000;
array[57239] <= 16'b0000_0000_0000_0000;
array[57240] <= 16'b0000_0000_0000_0000;
array[57241] <= 16'b0000_0000_0000_0000;
array[57242] <= 16'b0000_0000_0000_0000;
array[57243] <= 16'b0000_0000_0000_0000;
array[57244] <= 16'b0000_0000_0000_0000;
array[57245] <= 16'b0000_0000_0000_0000;
array[57246] <= 16'b0000_0000_0000_0000;
array[57247] <= 16'b0000_0000_0000_0000;
array[57248] <= 16'b0000_0000_0000_0000;
array[57249] <= 16'b0000_0000_0000_0000;
array[57250] <= 16'b0000_0000_0000_0000;
array[57251] <= 16'b0000_0000_0000_0000;
array[57252] <= 16'b0000_0000_0000_0000;
array[57253] <= 16'b0000_0000_0000_0000;
array[57254] <= 16'b0000_0000_0000_0000;
array[57255] <= 16'b0000_0000_0000_0000;
array[57256] <= 16'b0000_0000_0000_0000;
array[57257] <= 16'b0000_0000_0000_0000;
array[57258] <= 16'b0000_0000_0000_0000;
array[57259] <= 16'b0000_0000_0000_0000;
array[57260] <= 16'b0000_0000_0000_0000;
array[57261] <= 16'b0000_0000_0000_0000;
array[57262] <= 16'b0000_0000_0000_0000;
array[57263] <= 16'b0000_0000_0000_0000;
array[57264] <= 16'b0000_0000_0000_0000;
array[57265] <= 16'b0000_0000_0000_0000;
array[57266] <= 16'b0000_0000_0000_0000;
array[57267] <= 16'b0000_0000_0000_0000;
array[57268] <= 16'b0000_0000_0000_0000;
array[57269] <= 16'b0000_0000_0000_0000;
array[57270] <= 16'b0000_0000_0000_0000;
array[57271] <= 16'b0000_0000_0000_0000;
array[57272] <= 16'b0000_0000_0000_0000;
array[57273] <= 16'b0000_0000_0000_0000;
array[57274] <= 16'b0000_0000_0000_0000;
array[57275] <= 16'b0000_0000_0000_0000;
array[57276] <= 16'b0000_0000_0000_0000;
array[57277] <= 16'b0000_0000_0000_0000;
array[57278] <= 16'b0000_0000_0000_0000;
array[57279] <= 16'b0000_0000_0000_0000;
array[57280] <= 16'b0000_0000_0000_0000;
array[57281] <= 16'b0000_0000_0000_0000;
array[57282] <= 16'b0000_0000_0000_0000;
array[57283] <= 16'b0000_0000_0000_0000;
array[57284] <= 16'b0000_0000_0000_0000;
array[57285] <= 16'b0000_0000_0000_0000;
array[57286] <= 16'b0000_0000_0000_0000;
array[57287] <= 16'b0000_0000_0000_0000;
array[57288] <= 16'b0000_0000_0000_0000;
array[57289] <= 16'b0000_0000_0000_0000;
array[57290] <= 16'b0000_0000_0000_0000;
array[57291] <= 16'b0000_0000_0000_0000;
array[57292] <= 16'b0000_0000_0000_0000;
array[57293] <= 16'b0000_0000_0000_0000;
array[57294] <= 16'b0000_0000_0000_0000;
array[57295] <= 16'b0000_0000_0000_0000;
array[57296] <= 16'b0000_0000_0000_0000;
array[57297] <= 16'b0000_0000_0000_0000;
array[57298] <= 16'b0000_0000_0000_0000;
array[57299] <= 16'b0000_0000_0000_0000;
array[57300] <= 16'b0000_0000_0000_0000;
array[57301] <= 16'b0000_0000_0000_0000;
array[57302] <= 16'b0000_0000_0000_0000;
array[57303] <= 16'b0000_0000_0000_0000;
array[57304] <= 16'b0000_0000_0000_0000;
array[57305] <= 16'b0000_0000_0000_0000;
array[57306] <= 16'b0000_0000_0000_0000;
array[57307] <= 16'b0000_0000_0000_0000;
array[57308] <= 16'b0000_0000_0000_0000;
array[57309] <= 16'b0000_0000_0000_0000;
array[57310] <= 16'b0000_0000_0000_0000;
array[57311] <= 16'b0000_0000_0000_0000;
array[57312] <= 16'b0000_0000_0000_0000;
array[57313] <= 16'b0000_0000_0000_0000;
array[57314] <= 16'b0000_0000_0000_0000;
array[57315] <= 16'b0000_0000_0000_0000;
array[57316] <= 16'b0000_0000_0000_0000;
array[57317] <= 16'b0000_0000_0000_0000;
array[57318] <= 16'b0000_0000_0000_0000;
array[57319] <= 16'b0000_0000_0000_0000;
array[57320] <= 16'b0000_0000_0000_0000;
array[57321] <= 16'b0000_0000_0000_0000;
array[57322] <= 16'b0000_0000_0000_0000;
array[57323] <= 16'b0000_0000_0000_0000;
array[57324] <= 16'b0000_0000_0000_0000;
array[57325] <= 16'b0000_0000_0000_0000;
array[57326] <= 16'b0000_0000_0000_0000;
array[57327] <= 16'b0000_0000_0000_0000;
array[57328] <= 16'b0000_0000_0000_0000;
array[57329] <= 16'b0000_0000_0000_0000;
array[57330] <= 16'b0000_0000_0000_0000;
array[57331] <= 16'b0000_0000_0000_0000;
array[57332] <= 16'b0000_0000_0000_0000;
array[57333] <= 16'b0000_0000_0000_0000;
array[57334] <= 16'b0000_0000_0000_0000;
array[57335] <= 16'b0000_0000_0000_0000;
array[57336] <= 16'b0000_0000_0000_0000;
array[57337] <= 16'b0000_0000_0000_0000;
array[57338] <= 16'b0000_0000_0000_0000;
array[57339] <= 16'b0000_0000_0000_0000;
array[57340] <= 16'b0000_0000_0000_0000;
array[57341] <= 16'b0000_0000_0000_0000;
array[57342] <= 16'b0000_0000_0000_0000;
array[57343] <= 16'b0000_0000_0000_0000;
array[57344] <= 16'b0000_0000_0000_0000;
array[57345] <= 16'b0000_0000_0000_0000;
array[57346] <= 16'b0000_0000_0000_0000;
array[57347] <= 16'b0000_0000_0000_0000;
array[57348] <= 16'b0000_0000_0000_0000;
array[57349] <= 16'b0000_0000_0000_0000;
array[57350] <= 16'b0000_0000_0000_0000;
array[57351] <= 16'b0000_0000_0000_0000;
array[57352] <= 16'b0000_0000_0000_0000;
array[57353] <= 16'b0000_0000_0000_0000;
array[57354] <= 16'b0000_0000_0000_0000;
array[57355] <= 16'b0000_0000_0000_0000;
array[57356] <= 16'b0000_0000_0000_0000;
array[57357] <= 16'b0000_0000_0000_0000;
array[57358] <= 16'b0000_0000_0000_0000;
array[57359] <= 16'b0000_0000_0000_0000;
array[57360] <= 16'b0000_0000_0000_0000;
array[57361] <= 16'b0000_0000_0000_0000;
array[57362] <= 16'b0000_0000_0000_0000;
array[57363] <= 16'b0000_0000_0000_0000;
array[57364] <= 16'b0000_0000_0000_0000;
array[57365] <= 16'b0000_0000_0000_0000;
array[57366] <= 16'b0000_0000_0000_0000;
array[57367] <= 16'b0000_0000_0000_0000;
array[57368] <= 16'b0000_0000_0000_0000;
array[57369] <= 16'b0000_0000_0000_0000;
array[57370] <= 16'b0000_0000_0000_0000;
array[57371] <= 16'b0000_0000_0000_0000;
array[57372] <= 16'b0000_0000_0000_0000;
array[57373] <= 16'b0000_0000_0000_0000;
array[57374] <= 16'b0000_0000_0000_0000;
array[57375] <= 16'b0000_0000_0000_0000;
array[57376] <= 16'b0000_0000_0000_0000;
array[57377] <= 16'b0000_0000_0000_0000;
array[57378] <= 16'b0000_0000_0000_0000;
array[57379] <= 16'b0000_0000_0000_0000;
array[57380] <= 16'b0000_0000_0000_0000;
array[57381] <= 16'b0000_0000_0000_0000;
array[57382] <= 16'b0000_0000_0000_0000;
array[57383] <= 16'b0000_0000_0000_0000;
array[57384] <= 16'b0000_0000_0000_0000;
array[57385] <= 16'b0000_0000_0000_0000;
array[57386] <= 16'b0000_0000_0000_0000;
array[57387] <= 16'b0000_0000_0000_0000;
array[57388] <= 16'b0000_0000_0000_0000;
array[57389] <= 16'b0000_0000_0000_0000;
array[57390] <= 16'b0000_0000_0000_0000;
array[57391] <= 16'b0000_0000_0000_0000;
array[57392] <= 16'b0000_0000_0000_0000;
array[57393] <= 16'b0000_0000_0000_0000;
array[57394] <= 16'b0000_0000_0000_0000;
array[57395] <= 16'b0000_0000_0000_0000;
array[57396] <= 16'b0000_0000_0000_0000;
array[57397] <= 16'b0000_0000_0000_0000;
array[57398] <= 16'b0000_0000_0000_0000;
array[57399] <= 16'b0000_0000_0000_0000;
array[57400] <= 16'b0000_0000_0000_0000;
array[57401] <= 16'b0000_0000_0000_0000;
array[57402] <= 16'b0000_0000_0000_0000;
array[57403] <= 16'b0000_0000_0000_0000;
array[57404] <= 16'b0000_0000_0000_0000;
array[57405] <= 16'b0000_0000_0000_0000;
array[57406] <= 16'b0000_0000_0000_0000;
array[57407] <= 16'b0000_0000_0000_0000;
array[57408] <= 16'b0000_0000_0000_0000;
array[57409] <= 16'b0000_0000_0000_0000;
array[57410] <= 16'b0000_0000_0000_0000;
array[57411] <= 16'b0000_0000_0000_0000;
array[57412] <= 16'b0000_0000_0000_0000;
array[57413] <= 16'b0000_0000_0000_0000;
array[57414] <= 16'b0000_0000_0000_0000;
array[57415] <= 16'b0000_0000_0000_0000;
array[57416] <= 16'b0000_0000_0000_0000;
array[57417] <= 16'b0000_0000_0000_0000;
array[57418] <= 16'b0000_0000_0000_0000;
array[57419] <= 16'b0000_0000_0000_0000;
array[57420] <= 16'b0000_0000_0000_0000;
array[57421] <= 16'b0000_0000_0000_0000;
array[57422] <= 16'b0000_0000_0000_0000;
array[57423] <= 16'b0000_0000_0000_0000;
array[57424] <= 16'b0000_0000_0000_0000;
array[57425] <= 16'b0000_0000_0000_0000;
array[57426] <= 16'b0000_0000_0000_0000;
array[57427] <= 16'b0000_0000_0000_0000;
array[57428] <= 16'b0000_0000_0000_0000;
array[57429] <= 16'b0000_0000_0000_0000;
array[57430] <= 16'b0000_0000_0000_0000;
array[57431] <= 16'b0000_0000_0000_0000;
array[57432] <= 16'b0000_0000_0000_0000;
array[57433] <= 16'b0000_0000_0000_0000;
array[57434] <= 16'b0000_0000_0000_0000;
array[57435] <= 16'b0000_0000_0000_0000;
array[57436] <= 16'b0000_0000_0000_0000;
array[57437] <= 16'b0000_0000_0000_0000;
array[57438] <= 16'b0000_0000_0000_0000;
array[57439] <= 16'b0000_0000_0000_0000;
array[57440] <= 16'b0000_0000_0000_0000;
array[57441] <= 16'b0000_0000_0000_0000;
array[57442] <= 16'b0000_0000_0000_0000;
array[57443] <= 16'b0000_0000_0000_0000;
array[57444] <= 16'b0000_0000_0000_0000;
array[57445] <= 16'b0000_0000_0000_0000;
array[57446] <= 16'b0000_0000_0000_0000;
array[57447] <= 16'b0000_0000_0000_0000;
array[57448] <= 16'b0000_0000_0000_0000;
array[57449] <= 16'b0000_0000_0000_0000;
array[57450] <= 16'b0000_0000_0000_0000;
array[57451] <= 16'b0000_0000_0000_0000;
array[57452] <= 16'b0000_0000_0000_0000;
array[57453] <= 16'b0000_0000_0000_0000;
array[57454] <= 16'b0000_0000_0000_0000;
array[57455] <= 16'b0000_0000_0000_0000;
array[57456] <= 16'b0000_0000_0000_0000;
array[57457] <= 16'b0000_0000_0000_0000;
array[57458] <= 16'b0000_0000_0000_0000;
array[57459] <= 16'b0000_0000_0000_0000;
array[57460] <= 16'b0000_0000_0000_0000;
array[57461] <= 16'b0000_0000_0000_0000;
array[57462] <= 16'b0000_0000_0000_0000;
array[57463] <= 16'b0000_0000_0000_0000;
array[57464] <= 16'b0000_0000_0000_0000;
array[57465] <= 16'b0000_0000_0000_0000;
array[57466] <= 16'b0000_0000_0000_0000;
array[57467] <= 16'b0000_0000_0000_0000;
array[57468] <= 16'b0000_0000_0000_0000;
array[57469] <= 16'b0000_0000_0000_0000;
array[57470] <= 16'b0000_0000_0000_0000;
array[57471] <= 16'b0000_0000_0000_0000;
array[57472] <= 16'b0000_0000_0000_0000;
array[57473] <= 16'b0000_0000_0000_0000;
array[57474] <= 16'b0000_0000_0000_0000;
array[57475] <= 16'b0000_0000_0000_0000;
array[57476] <= 16'b0000_0000_0000_0000;
array[57477] <= 16'b0000_0000_0000_0000;
array[57478] <= 16'b0000_0000_0000_0000;
array[57479] <= 16'b0000_0000_0000_0000;
array[57480] <= 16'b0000_0000_0000_0000;
array[57481] <= 16'b0000_0000_0000_0000;
array[57482] <= 16'b0000_0000_0000_0000;
array[57483] <= 16'b0000_0000_0000_0000;
array[57484] <= 16'b0000_0000_0000_0000;
array[57485] <= 16'b0000_0000_0000_0000;
array[57486] <= 16'b0000_0000_0000_0000;
array[57487] <= 16'b0000_0000_0000_0000;
array[57488] <= 16'b0000_0000_0000_0000;
array[57489] <= 16'b0000_0000_0000_0000;
array[57490] <= 16'b0000_0000_0000_0000;
array[57491] <= 16'b0000_0000_0000_0000;
array[57492] <= 16'b0000_0000_0000_0000;
array[57493] <= 16'b0000_0000_0000_0000;
array[57494] <= 16'b0000_0000_0000_0000;
array[57495] <= 16'b0000_0000_0000_0000;
array[57496] <= 16'b0000_0000_0000_0000;
array[57497] <= 16'b0000_0000_0000_0000;
array[57498] <= 16'b0000_0000_0000_0000;
array[57499] <= 16'b0000_0000_0000_0000;
array[57500] <= 16'b0000_0000_0000_0000;
array[57501] <= 16'b0000_0000_0000_0000;
array[57502] <= 16'b0000_0000_0000_0000;
array[57503] <= 16'b0000_0000_0000_0000;
array[57504] <= 16'b0000_0000_0000_0000;
array[57505] <= 16'b0000_0000_0000_0000;
array[57506] <= 16'b0000_0000_0000_0000;
array[57507] <= 16'b0000_0000_0000_0000;
array[57508] <= 16'b0000_0000_0000_0000;
array[57509] <= 16'b0000_0000_0000_0000;
array[57510] <= 16'b0000_0000_0000_0000;
array[57511] <= 16'b0000_0000_0000_0000;
array[57512] <= 16'b0000_0000_0000_0000;
array[57513] <= 16'b0000_0000_0000_0000;
array[57514] <= 16'b0000_0000_0000_0000;
array[57515] <= 16'b0000_0000_0000_0000;
array[57516] <= 16'b0000_0000_0000_0000;
array[57517] <= 16'b0000_0000_0000_0000;
array[57518] <= 16'b0000_0000_0000_0000;
array[57519] <= 16'b0000_0000_0000_0000;
array[57520] <= 16'b0000_0000_0000_0000;
array[57521] <= 16'b0000_0000_0000_0000;
array[57522] <= 16'b0000_0000_0000_0000;
array[57523] <= 16'b0000_0000_0000_0000;
array[57524] <= 16'b0000_0000_0000_0000;
array[57525] <= 16'b0000_0000_0000_0000;
array[57526] <= 16'b0000_0000_0000_0000;
array[57527] <= 16'b0000_0000_0000_0000;
array[57528] <= 16'b0000_0000_0000_0000;
array[57529] <= 16'b0000_0000_0000_0000;
array[57530] <= 16'b0000_0000_0000_0000;
array[57531] <= 16'b0000_0000_0000_0000;
array[57532] <= 16'b0000_0000_0000_0000;
array[57533] <= 16'b0000_0000_0000_0000;
array[57534] <= 16'b0000_0000_0000_0000;
array[57535] <= 16'b0000_0000_0000_0000;
array[57536] <= 16'b0000_0000_0000_0000;
array[57537] <= 16'b0000_0000_0000_0000;
array[57538] <= 16'b0000_0000_0000_0000;
array[57539] <= 16'b0000_0000_0000_0000;
array[57540] <= 16'b0000_0000_0000_0000;
array[57541] <= 16'b0000_0000_0000_0000;
array[57542] <= 16'b0000_0000_0000_0000;
array[57543] <= 16'b0000_0000_0000_0000;
array[57544] <= 16'b0000_0000_0000_0000;
array[57545] <= 16'b0000_0000_0000_0000;
array[57546] <= 16'b0000_0000_0000_0000;
array[57547] <= 16'b0000_0000_0000_0000;
array[57548] <= 16'b0000_0000_0000_0000;
array[57549] <= 16'b0000_0000_0000_0000;
array[57550] <= 16'b0000_0000_0000_0000;
array[57551] <= 16'b0000_0000_0000_0000;
array[57552] <= 16'b0000_0000_0000_0000;
array[57553] <= 16'b0000_0000_0000_0000;
array[57554] <= 16'b0000_0000_0000_0000;
array[57555] <= 16'b0000_0000_0000_0000;
array[57556] <= 16'b0000_0000_0000_0000;
array[57557] <= 16'b0000_0000_0000_0000;
array[57558] <= 16'b0000_0000_0000_0000;
array[57559] <= 16'b0000_0000_0000_0000;
array[57560] <= 16'b0000_0000_0000_0000;
array[57561] <= 16'b0000_0000_0000_0000;
array[57562] <= 16'b0000_0000_0000_0000;
array[57563] <= 16'b0000_0000_0000_0000;
array[57564] <= 16'b0000_0000_0000_0000;
array[57565] <= 16'b0000_0000_0000_0000;
array[57566] <= 16'b0000_0000_0000_0000;
array[57567] <= 16'b0000_0000_0000_0000;
array[57568] <= 16'b0000_0000_0000_0000;
array[57569] <= 16'b0000_0000_0000_0000;
array[57570] <= 16'b0000_0000_0000_0000;
array[57571] <= 16'b0000_0000_0000_0000;
array[57572] <= 16'b0000_0000_0000_0000;
array[57573] <= 16'b0000_0000_0000_0000;
array[57574] <= 16'b0000_0000_0000_0000;
array[57575] <= 16'b0000_0000_0000_0000;
array[57576] <= 16'b0000_0000_0000_0000;
array[57577] <= 16'b0000_0000_0000_0000;
array[57578] <= 16'b0000_0000_0000_0000;
array[57579] <= 16'b0000_0000_0000_0000;
array[57580] <= 16'b0000_0000_0000_0000;
array[57581] <= 16'b0000_0000_0000_0000;
array[57582] <= 16'b0000_0000_0000_0000;
array[57583] <= 16'b0000_0000_0000_0000;
array[57584] <= 16'b0000_0000_0000_0000;
array[57585] <= 16'b0000_0000_0000_0000;
array[57586] <= 16'b0000_0000_0000_0000;
array[57587] <= 16'b0000_0000_0000_0000;
array[57588] <= 16'b0000_0000_0000_0000;
array[57589] <= 16'b0000_0000_0000_0000;
array[57590] <= 16'b0000_0000_0000_0000;
array[57591] <= 16'b0000_0000_0000_0000;
array[57592] <= 16'b0000_0000_0000_0000;
array[57593] <= 16'b0000_0000_0000_0000;
array[57594] <= 16'b0000_0000_0000_0000;
array[57595] <= 16'b0000_0000_0000_0000;
array[57596] <= 16'b0000_0000_0000_0000;
array[57597] <= 16'b0000_0000_0000_0000;
array[57598] <= 16'b0000_0000_0000_0000;
array[57599] <= 16'b0000_0000_0000_0000;
array[57600] <= 16'b0000_0000_0000_0000;
array[57601] <= 16'b0000_0000_0000_0000;
array[57602] <= 16'b0000_0000_0000_0000;
array[57603] <= 16'b0000_0000_0000_0000;
array[57604] <= 16'b0000_0000_0000_0000;
array[57605] <= 16'b0000_0000_0000_0000;
array[57606] <= 16'b0000_0000_0000_0000;
array[57607] <= 16'b0000_0000_0000_0000;
array[57608] <= 16'b0000_0000_0000_0000;
array[57609] <= 16'b0000_0000_0000_0000;
array[57610] <= 16'b0000_0000_0000_0000;
array[57611] <= 16'b0000_0000_0000_0000;
array[57612] <= 16'b0000_0000_0000_0000;
array[57613] <= 16'b0000_0000_0000_0000;
array[57614] <= 16'b0000_0000_0000_0000;
array[57615] <= 16'b0000_0000_0000_0000;
array[57616] <= 16'b0000_0000_0000_0000;
array[57617] <= 16'b0000_0000_0000_0000;
array[57618] <= 16'b0000_0000_0000_0000;
array[57619] <= 16'b0000_0000_0000_0000;
array[57620] <= 16'b0000_0000_0000_0000;
array[57621] <= 16'b0000_0000_0000_0000;
array[57622] <= 16'b0000_0000_0000_0000;
array[57623] <= 16'b0000_0000_0000_0000;
array[57624] <= 16'b0000_0000_0000_0000;
array[57625] <= 16'b0000_0000_0000_0000;
array[57626] <= 16'b0000_0000_0000_0000;
array[57627] <= 16'b0000_0000_0000_0000;
array[57628] <= 16'b0000_0000_0000_0000;
array[57629] <= 16'b0000_0000_0000_0000;
array[57630] <= 16'b0000_0000_0000_0000;
array[57631] <= 16'b0000_0000_0000_0000;
array[57632] <= 16'b0000_0000_0000_0000;
array[57633] <= 16'b0000_0000_0000_0000;
array[57634] <= 16'b0000_0000_0000_0000;
array[57635] <= 16'b0000_0000_0000_0000;
array[57636] <= 16'b0000_0000_0000_0000;
array[57637] <= 16'b0000_0000_0000_0000;
array[57638] <= 16'b0000_0000_0000_0000;
array[57639] <= 16'b0000_0000_0000_0000;
array[57640] <= 16'b0000_0000_0000_0000;
array[57641] <= 16'b0000_0000_0000_0000;
array[57642] <= 16'b0000_0000_0000_0000;
array[57643] <= 16'b0000_0000_0000_0000;
array[57644] <= 16'b0000_0000_0000_0000;
array[57645] <= 16'b0000_0000_0000_0000;
array[57646] <= 16'b0000_0000_0000_0000;
array[57647] <= 16'b0000_0000_0000_0000;
array[57648] <= 16'b0000_0000_0000_0000;
array[57649] <= 16'b0000_0000_0000_0000;
array[57650] <= 16'b0000_0000_0000_0000;
array[57651] <= 16'b0000_0000_0000_0000;
array[57652] <= 16'b0000_0000_0000_0000;
array[57653] <= 16'b0000_0000_0000_0000;
array[57654] <= 16'b0000_0000_0000_0000;
array[57655] <= 16'b0000_0000_0000_0000;
array[57656] <= 16'b0000_0000_0000_0000;
array[57657] <= 16'b0000_0000_0000_0000;
array[57658] <= 16'b0000_0000_0000_0000;
array[57659] <= 16'b0000_0000_0000_0000;
array[57660] <= 16'b0000_0000_0000_0000;
array[57661] <= 16'b0000_0000_0000_0000;
array[57662] <= 16'b0000_0000_0000_0000;
array[57663] <= 16'b0000_0000_0000_0000;
array[57664] <= 16'b0000_0000_0000_0000;
array[57665] <= 16'b0000_0000_0000_0000;
array[57666] <= 16'b0000_0000_0000_0000;
array[57667] <= 16'b0000_0000_0000_0000;
array[57668] <= 16'b0000_0000_0000_0000;
array[57669] <= 16'b0000_0000_0000_0000;
array[57670] <= 16'b0000_0000_0000_0000;
array[57671] <= 16'b0000_0000_0000_0000;
array[57672] <= 16'b0000_0000_0000_0000;
array[57673] <= 16'b0000_0000_0000_0000;
array[57674] <= 16'b0000_0000_0000_0000;
array[57675] <= 16'b0000_0000_0000_0000;
array[57676] <= 16'b0000_0000_0000_0000;
array[57677] <= 16'b0000_0000_0000_0000;
array[57678] <= 16'b0000_0000_0000_0000;
array[57679] <= 16'b0000_0000_0000_0000;
array[57680] <= 16'b0000_0000_0000_0000;
array[57681] <= 16'b0000_0000_0000_0000;
array[57682] <= 16'b0000_0000_0000_0000;
array[57683] <= 16'b0000_0000_0000_0000;
array[57684] <= 16'b0000_0000_0000_0000;
array[57685] <= 16'b0000_0000_0000_0000;
array[57686] <= 16'b0000_0000_0000_0000;
array[57687] <= 16'b0000_0000_0000_0000;
array[57688] <= 16'b0000_0000_0000_0000;
array[57689] <= 16'b0000_0000_0000_0000;
array[57690] <= 16'b0000_0000_0000_0000;
array[57691] <= 16'b0000_0000_0000_0000;
array[57692] <= 16'b0000_0000_0000_0000;
array[57693] <= 16'b0000_0000_0000_0000;
array[57694] <= 16'b0000_0000_0000_0000;
array[57695] <= 16'b0000_0000_0000_0000;
array[57696] <= 16'b0000_0000_0000_0000;
array[57697] <= 16'b0000_0000_0000_0000;
array[57698] <= 16'b0000_0000_0000_0000;
array[57699] <= 16'b0000_0000_0000_0000;
array[57700] <= 16'b0000_0000_0000_0000;
array[57701] <= 16'b0000_0000_0000_0000;
array[57702] <= 16'b0000_0000_0000_0000;
array[57703] <= 16'b0000_0000_0000_0000;
array[57704] <= 16'b0000_0000_0000_0000;
array[57705] <= 16'b0000_0000_0000_0000;
array[57706] <= 16'b0000_0000_0000_0000;
array[57707] <= 16'b0000_0000_0000_0000;
array[57708] <= 16'b0000_0000_0000_0000;
array[57709] <= 16'b0000_0000_0000_0000;
array[57710] <= 16'b0000_0000_0000_0000;
array[57711] <= 16'b0000_0000_0000_0000;
array[57712] <= 16'b0000_0000_0000_0000;
array[57713] <= 16'b0000_0000_0000_0000;
array[57714] <= 16'b0000_0000_0000_0000;
array[57715] <= 16'b0000_0000_0000_0000;
array[57716] <= 16'b0000_0000_0000_0000;
array[57717] <= 16'b0000_0000_0000_0000;
array[57718] <= 16'b0000_0000_0000_0000;
array[57719] <= 16'b0000_0000_0000_0000;
array[57720] <= 16'b0000_0000_0000_0000;
array[57721] <= 16'b0000_0000_0000_0000;
array[57722] <= 16'b0000_0000_0000_0000;
array[57723] <= 16'b0000_0000_0000_0000;
array[57724] <= 16'b0000_0000_0000_0000;
array[57725] <= 16'b0000_0000_0000_0000;
array[57726] <= 16'b0000_0000_0000_0000;
array[57727] <= 16'b0000_0000_0000_0000;
array[57728] <= 16'b0000_0000_0000_0000;
array[57729] <= 16'b0000_0000_0000_0000;
array[57730] <= 16'b0000_0000_0000_0000;
array[57731] <= 16'b0000_0000_0000_0000;
array[57732] <= 16'b0000_0000_0000_0000;
array[57733] <= 16'b0000_0000_0000_0000;
array[57734] <= 16'b0000_0000_0000_0000;
array[57735] <= 16'b0000_0000_0000_0000;
array[57736] <= 16'b0000_0000_0000_0000;
array[57737] <= 16'b0000_0000_0000_0000;
array[57738] <= 16'b0000_0000_0000_0000;
array[57739] <= 16'b0000_0000_0000_0000;
array[57740] <= 16'b0000_0000_0000_0000;
array[57741] <= 16'b0000_0000_0000_0000;
array[57742] <= 16'b0000_0000_0000_0000;
array[57743] <= 16'b0000_0000_0000_0000;
array[57744] <= 16'b0000_0000_0000_0000;
array[57745] <= 16'b0000_0000_0000_0000;
array[57746] <= 16'b0000_0000_0000_0000;
array[57747] <= 16'b0000_0000_0000_0000;
array[57748] <= 16'b0000_0000_0000_0000;
array[57749] <= 16'b0000_0000_0000_0000;
array[57750] <= 16'b0000_0000_0000_0000;
array[57751] <= 16'b0000_0000_0000_0000;
array[57752] <= 16'b0000_0000_0000_0000;
array[57753] <= 16'b0000_0000_0000_0000;
array[57754] <= 16'b0000_0000_0000_0000;
array[57755] <= 16'b0000_0000_0000_0000;
array[57756] <= 16'b0000_0000_0000_0000;
array[57757] <= 16'b0000_0000_0000_0000;
array[57758] <= 16'b0000_0000_0000_0000;
array[57759] <= 16'b0000_0000_0000_0000;
array[57760] <= 16'b0000_0000_0000_0000;
array[57761] <= 16'b0000_0000_0000_0000;
array[57762] <= 16'b0000_0000_0000_0000;
array[57763] <= 16'b0000_0000_0000_0000;
array[57764] <= 16'b0000_0000_0000_0000;
array[57765] <= 16'b0000_0000_0000_0000;
array[57766] <= 16'b0000_0000_0000_0000;
array[57767] <= 16'b0000_0000_0000_0000;
array[57768] <= 16'b0000_0000_0000_0000;
array[57769] <= 16'b0000_0000_0000_0000;
array[57770] <= 16'b0000_0000_0000_0000;
array[57771] <= 16'b0000_0000_0000_0000;
array[57772] <= 16'b0000_0000_0000_0000;
array[57773] <= 16'b0000_0000_0000_0000;
array[57774] <= 16'b0000_0000_0000_0000;
array[57775] <= 16'b0000_0000_0000_0000;
array[57776] <= 16'b0000_0000_0000_0000;
array[57777] <= 16'b0000_0000_0000_0000;
array[57778] <= 16'b0000_0000_0000_0000;
array[57779] <= 16'b0000_0000_0000_0000;
array[57780] <= 16'b0000_0000_0000_0000;
array[57781] <= 16'b0000_0000_0000_0000;
array[57782] <= 16'b0000_0000_0000_0000;
array[57783] <= 16'b0000_0000_0000_0000;
array[57784] <= 16'b0000_0000_0000_0000;
array[57785] <= 16'b0000_0000_0000_0000;
array[57786] <= 16'b0000_0000_0000_0000;
array[57787] <= 16'b0000_0000_0000_0000;
array[57788] <= 16'b0000_0000_0000_0000;
array[57789] <= 16'b0000_0000_0000_0000;
array[57790] <= 16'b0000_0000_0000_0000;
array[57791] <= 16'b0000_0000_0000_0000;
array[57792] <= 16'b0000_0000_0000_0000;
array[57793] <= 16'b0000_0000_0000_0000;
array[57794] <= 16'b0000_0000_0000_0000;
array[57795] <= 16'b0000_0000_0000_0000;
array[57796] <= 16'b0000_0000_0000_0000;
array[57797] <= 16'b0000_0000_0000_0000;
array[57798] <= 16'b0000_0000_0000_0000;
array[57799] <= 16'b0000_0000_0000_0000;
array[57800] <= 16'b0000_0000_0000_0000;
array[57801] <= 16'b0000_0000_0000_0000;
array[57802] <= 16'b0000_0000_0000_0000;
array[57803] <= 16'b0000_0000_0000_0000;
array[57804] <= 16'b0000_0000_0000_0000;
array[57805] <= 16'b0000_0000_0000_0000;
array[57806] <= 16'b0000_0000_0000_0000;
array[57807] <= 16'b0000_0000_0000_0000;
array[57808] <= 16'b0000_0000_0000_0000;
array[57809] <= 16'b0000_0000_0000_0000;
array[57810] <= 16'b0000_0000_0000_0000;
array[57811] <= 16'b0000_0000_0000_0000;
array[57812] <= 16'b0000_0000_0000_0000;
array[57813] <= 16'b0000_0000_0000_0000;
array[57814] <= 16'b0000_0000_0000_0000;
array[57815] <= 16'b0000_0000_0000_0000;
array[57816] <= 16'b0000_0000_0000_0000;
array[57817] <= 16'b0000_0000_0000_0000;
array[57818] <= 16'b0000_0000_0000_0000;
array[57819] <= 16'b0000_0000_0000_0000;
array[57820] <= 16'b0000_0000_0000_0000;
array[57821] <= 16'b0000_0000_0000_0000;
array[57822] <= 16'b0000_0000_0000_0000;
array[57823] <= 16'b0000_0000_0000_0000;
array[57824] <= 16'b0000_0000_0000_0000;
array[57825] <= 16'b0000_0000_0000_0000;
array[57826] <= 16'b0000_0000_0000_0000;
array[57827] <= 16'b0000_0000_0000_0000;
array[57828] <= 16'b0000_0000_0000_0000;
array[57829] <= 16'b0000_0000_0000_0000;
array[57830] <= 16'b0000_0000_0000_0000;
array[57831] <= 16'b0000_0000_0000_0000;
array[57832] <= 16'b0000_0000_0000_0000;
array[57833] <= 16'b0000_0000_0000_0000;
array[57834] <= 16'b0000_0000_0000_0000;
array[57835] <= 16'b0000_0000_0000_0000;
array[57836] <= 16'b0000_0000_0000_0000;
array[57837] <= 16'b0000_0000_0000_0000;
array[57838] <= 16'b0000_0000_0000_0000;
array[57839] <= 16'b0000_0000_0000_0000;
array[57840] <= 16'b0000_0000_0000_0000;
array[57841] <= 16'b0000_0000_0000_0000;
array[57842] <= 16'b0000_0000_0000_0000;
array[57843] <= 16'b0000_0000_0000_0000;
array[57844] <= 16'b0000_0000_0000_0000;
array[57845] <= 16'b0000_0000_0000_0000;
array[57846] <= 16'b0000_0000_0000_0000;
array[57847] <= 16'b0000_0000_0000_0000;
array[57848] <= 16'b0000_0000_0000_0000;
array[57849] <= 16'b0000_0000_0000_0000;
array[57850] <= 16'b0000_0000_0000_0000;
array[57851] <= 16'b0000_0000_0000_0000;
array[57852] <= 16'b0000_0000_0000_0000;
array[57853] <= 16'b0000_0000_0000_0000;
array[57854] <= 16'b0000_0000_0000_0000;
array[57855] <= 16'b0000_0000_0000_0000;
array[57856] <= 16'b0000_0000_0000_0000;
array[57857] <= 16'b0000_0000_0000_0000;
array[57858] <= 16'b0000_0000_0000_0000;
array[57859] <= 16'b0000_0000_0000_0000;
array[57860] <= 16'b0000_0000_0000_0000;
array[57861] <= 16'b0000_0000_0000_0000;
array[57862] <= 16'b0000_0000_0000_0000;
array[57863] <= 16'b0000_0000_0000_0000;
array[57864] <= 16'b0000_0000_0000_0000;
array[57865] <= 16'b0000_0000_0000_0000;
array[57866] <= 16'b0000_0000_0000_0000;
array[57867] <= 16'b0000_0000_0000_0000;
array[57868] <= 16'b0000_0000_0000_0000;
array[57869] <= 16'b0000_0000_0000_0000;
array[57870] <= 16'b0000_0000_0000_0000;
array[57871] <= 16'b0000_0000_0000_0000;
array[57872] <= 16'b0000_0000_0000_0000;
array[57873] <= 16'b0000_0000_0000_0000;
array[57874] <= 16'b0000_0000_0000_0000;
array[57875] <= 16'b0000_0000_0000_0000;
array[57876] <= 16'b0000_0000_0000_0000;
array[57877] <= 16'b0000_0000_0000_0000;
array[57878] <= 16'b0000_0000_0000_0000;
array[57879] <= 16'b0000_0000_0000_0000;
array[57880] <= 16'b0000_0000_0000_0000;
array[57881] <= 16'b0000_0000_0000_0000;
array[57882] <= 16'b0000_0000_0000_0000;
array[57883] <= 16'b0000_0000_0000_0000;
array[57884] <= 16'b0000_0000_0000_0000;
array[57885] <= 16'b0000_0000_0000_0000;
array[57886] <= 16'b0000_0000_0000_0000;
array[57887] <= 16'b0000_0000_0000_0000;
array[57888] <= 16'b0000_0000_0000_0000;
array[57889] <= 16'b0000_0000_0000_0000;
array[57890] <= 16'b0000_0000_0000_0000;
array[57891] <= 16'b0000_0000_0000_0000;
array[57892] <= 16'b0000_0000_0000_0000;
array[57893] <= 16'b0000_0000_0000_0000;
array[57894] <= 16'b0000_0000_0000_0000;
array[57895] <= 16'b0000_0000_0000_0000;
array[57896] <= 16'b0000_0000_0000_0000;
array[57897] <= 16'b0000_0000_0000_0000;
array[57898] <= 16'b0000_0000_0000_0000;
array[57899] <= 16'b0000_0000_0000_0000;
array[57900] <= 16'b0000_0000_0000_0000;
array[57901] <= 16'b0000_0000_0000_0000;
array[57902] <= 16'b0000_0000_0000_0000;
array[57903] <= 16'b0000_0000_0000_0000;
array[57904] <= 16'b0000_0000_0000_0000;
array[57905] <= 16'b0000_0000_0000_0000;
array[57906] <= 16'b0000_0000_0000_0000;
array[57907] <= 16'b0000_0000_0000_0000;
array[57908] <= 16'b0000_0000_0000_0000;
array[57909] <= 16'b0000_0000_0000_0000;
array[57910] <= 16'b0000_0000_0000_0000;
array[57911] <= 16'b0000_0000_0000_0000;
array[57912] <= 16'b0000_0000_0000_0000;
array[57913] <= 16'b0000_0000_0000_0000;
array[57914] <= 16'b0000_0000_0000_0000;
array[57915] <= 16'b0000_0000_0000_0000;
array[57916] <= 16'b0000_0000_0000_0000;
array[57917] <= 16'b0000_0000_0000_0000;
array[57918] <= 16'b0000_0000_0000_0000;
array[57919] <= 16'b0000_0000_0000_0000;
array[57920] <= 16'b0000_0000_0000_0000;
array[57921] <= 16'b0000_0000_0000_0000;
array[57922] <= 16'b0000_0000_0000_0000;
array[57923] <= 16'b0000_0000_0000_0000;
array[57924] <= 16'b0000_0000_0000_0000;
array[57925] <= 16'b0000_0000_0000_0000;
array[57926] <= 16'b0000_0000_0000_0000;
array[57927] <= 16'b0000_0000_0000_0000;
array[57928] <= 16'b0000_0000_0000_0000;
array[57929] <= 16'b0000_0000_0000_0000;
array[57930] <= 16'b0000_0000_0000_0000;
array[57931] <= 16'b0000_0000_0000_0000;
array[57932] <= 16'b0000_0000_0000_0000;
array[57933] <= 16'b0000_0000_0000_0000;
array[57934] <= 16'b0000_0000_0000_0000;
array[57935] <= 16'b0000_0000_0000_0000;
array[57936] <= 16'b0000_0000_0000_0000;
array[57937] <= 16'b0000_0000_0000_0000;
array[57938] <= 16'b0000_0000_0000_0000;
array[57939] <= 16'b0000_0000_0000_0000;
array[57940] <= 16'b0000_0000_0000_0000;
array[57941] <= 16'b0000_0000_0000_0000;
array[57942] <= 16'b0000_0000_0000_0000;
array[57943] <= 16'b0000_0000_0000_0000;
array[57944] <= 16'b0000_0000_0000_0000;
array[57945] <= 16'b0000_0000_0000_0000;
array[57946] <= 16'b0000_0000_0000_0000;
array[57947] <= 16'b0000_0000_0000_0000;
array[57948] <= 16'b0000_0000_0000_0000;
array[57949] <= 16'b0000_0000_0000_0000;
array[57950] <= 16'b0000_0000_0000_0000;
array[57951] <= 16'b0000_0000_0000_0000;
array[57952] <= 16'b0000_0000_0000_0000;
array[57953] <= 16'b0000_0000_0000_0000;
array[57954] <= 16'b0000_0000_0000_0000;
array[57955] <= 16'b0000_0000_0000_0000;
array[57956] <= 16'b0000_0000_0000_0000;
array[57957] <= 16'b0000_0000_0000_0000;
array[57958] <= 16'b0000_0000_0000_0000;
array[57959] <= 16'b0000_0000_0000_0000;
array[57960] <= 16'b0000_0000_0000_0000;
array[57961] <= 16'b0000_0000_0000_0000;
array[57962] <= 16'b0000_0000_0000_0000;
array[57963] <= 16'b0000_0000_0000_0000;
array[57964] <= 16'b0000_0000_0000_0000;
array[57965] <= 16'b0000_0000_0000_0000;
array[57966] <= 16'b0000_0000_0000_0000;
array[57967] <= 16'b0000_0000_0000_0000;
array[57968] <= 16'b0000_0000_0000_0000;
array[57969] <= 16'b0000_0000_0000_0000;
array[57970] <= 16'b0000_0000_0000_0000;
array[57971] <= 16'b0000_0000_0000_0000;
array[57972] <= 16'b0000_0000_0000_0000;
array[57973] <= 16'b0000_0000_0000_0000;
array[57974] <= 16'b0000_0000_0000_0000;
array[57975] <= 16'b0000_0000_0000_0000;
array[57976] <= 16'b0000_0000_0000_0000;
array[57977] <= 16'b0000_0000_0000_0000;
array[57978] <= 16'b0000_0000_0000_0000;
array[57979] <= 16'b0000_0000_0000_0000;
array[57980] <= 16'b0000_0000_0000_0000;
array[57981] <= 16'b0000_0000_0000_0000;
array[57982] <= 16'b0000_0000_0000_0000;
array[57983] <= 16'b0000_0000_0000_0000;
array[57984] <= 16'b0000_0000_0000_0000;
array[57985] <= 16'b0000_0000_0000_0000;
array[57986] <= 16'b0000_0000_0000_0000;
array[57987] <= 16'b0000_0000_0000_0000;
array[57988] <= 16'b0000_0000_0000_0000;
array[57989] <= 16'b0000_0000_0000_0000;
array[57990] <= 16'b0000_0000_0000_0000;
array[57991] <= 16'b0000_0000_0000_0000;
array[57992] <= 16'b0000_0000_0000_0000;
array[57993] <= 16'b0000_0000_0000_0000;
array[57994] <= 16'b0000_0000_0000_0000;
array[57995] <= 16'b0000_0000_0000_0000;
array[57996] <= 16'b0000_0000_0000_0000;
array[57997] <= 16'b0000_0000_0000_0000;
array[57998] <= 16'b0000_0000_0000_0000;
array[57999] <= 16'b0000_0000_0000_0000;
array[58000] <= 16'b0000_0000_0000_0000;
array[58001] <= 16'b0000_0000_0000_0000;
array[58002] <= 16'b0000_0000_0000_0000;
array[58003] <= 16'b0000_0000_0000_0000;
array[58004] <= 16'b0000_0000_0000_0000;
array[58005] <= 16'b0000_0000_0000_0000;
array[58006] <= 16'b0000_0000_0000_0000;
array[58007] <= 16'b0000_0000_0000_0000;
array[58008] <= 16'b0000_0000_0000_0000;
array[58009] <= 16'b0000_0000_0000_0000;
array[58010] <= 16'b0000_0000_0000_0000;
array[58011] <= 16'b0000_0000_0000_0000;
array[58012] <= 16'b0000_0000_0000_0000;
array[58013] <= 16'b0000_0000_0000_0000;
array[58014] <= 16'b0000_0000_0000_0000;
array[58015] <= 16'b0000_0000_0000_0000;
array[58016] <= 16'b0000_0000_0000_0000;
array[58017] <= 16'b0000_0000_0000_0000;
array[58018] <= 16'b0000_0000_0000_0000;
array[58019] <= 16'b0000_0000_0000_0000;
array[58020] <= 16'b0000_0000_0000_0000;
array[58021] <= 16'b0000_0000_0000_0000;
array[58022] <= 16'b0000_0000_0000_0000;
array[58023] <= 16'b0000_0000_0000_0000;
array[58024] <= 16'b0000_0000_0000_0000;
array[58025] <= 16'b0000_0000_0000_0000;
array[58026] <= 16'b0000_0000_0000_0000;
array[58027] <= 16'b0000_0000_0000_0000;
array[58028] <= 16'b0000_0000_0000_0000;
array[58029] <= 16'b0000_0000_0000_0000;
array[58030] <= 16'b0000_0000_0000_0000;
array[58031] <= 16'b0000_0000_0000_0000;
array[58032] <= 16'b0000_0000_0000_0000;
array[58033] <= 16'b0000_0000_0000_0000;
array[58034] <= 16'b0000_0000_0000_0000;
array[58035] <= 16'b0000_0000_0000_0000;
array[58036] <= 16'b0000_0000_0000_0000;
array[58037] <= 16'b0000_0000_0000_0000;
array[58038] <= 16'b0000_0000_0000_0000;
array[58039] <= 16'b0000_0000_0000_0000;
array[58040] <= 16'b0000_0000_0000_0000;
array[58041] <= 16'b0000_0000_0000_0000;
array[58042] <= 16'b0000_0000_0000_0000;
array[58043] <= 16'b0000_0000_0000_0000;
array[58044] <= 16'b0000_0000_0000_0000;
array[58045] <= 16'b0000_0000_0000_0000;
array[58046] <= 16'b0000_0000_0000_0000;
array[58047] <= 16'b0000_0000_0000_0000;
array[58048] <= 16'b0000_0000_0000_0000;
array[58049] <= 16'b0000_0000_0000_0000;
array[58050] <= 16'b0000_0000_0000_0000;
array[58051] <= 16'b0000_0000_0000_0000;
array[58052] <= 16'b0000_0000_0000_0000;
array[58053] <= 16'b0000_0000_0000_0000;
array[58054] <= 16'b0000_0000_0000_0000;
array[58055] <= 16'b0000_0000_0000_0000;
array[58056] <= 16'b0000_0000_0000_0000;
array[58057] <= 16'b0000_0000_0000_0000;
array[58058] <= 16'b0000_0000_0000_0000;
array[58059] <= 16'b0000_0000_0000_0000;
array[58060] <= 16'b0000_0000_0000_0000;
array[58061] <= 16'b0000_0000_0000_0000;
array[58062] <= 16'b0000_0000_0000_0000;
array[58063] <= 16'b0000_0000_0000_0000;
array[58064] <= 16'b0000_0000_0000_0000;
array[58065] <= 16'b0000_0000_0000_0000;
array[58066] <= 16'b0000_0000_0000_0000;
array[58067] <= 16'b0000_0000_0000_0000;
array[58068] <= 16'b0000_0000_0000_0000;
array[58069] <= 16'b0000_0000_0000_0000;
array[58070] <= 16'b0000_0000_0000_0000;
array[58071] <= 16'b0000_0000_0000_0000;
array[58072] <= 16'b0000_0000_0000_0000;
array[58073] <= 16'b0000_0000_0000_0000;
array[58074] <= 16'b0000_0000_0000_0000;
array[58075] <= 16'b0000_0000_0000_0000;
array[58076] <= 16'b0000_0000_0000_0000;
array[58077] <= 16'b0000_0000_0000_0000;
array[58078] <= 16'b0000_0000_0000_0000;
array[58079] <= 16'b0000_0000_0000_0000;
array[58080] <= 16'b0000_0000_0000_0000;
array[58081] <= 16'b0000_0000_0000_0000;
array[58082] <= 16'b0000_0000_0000_0000;
array[58083] <= 16'b0000_0000_0000_0000;
array[58084] <= 16'b0000_0000_0000_0000;
array[58085] <= 16'b0000_0000_0000_0000;
array[58086] <= 16'b0000_0000_0000_0000;
array[58087] <= 16'b0000_0000_0000_0000;
array[58088] <= 16'b0000_0000_0000_0000;
array[58089] <= 16'b0000_0000_0000_0000;
array[58090] <= 16'b0000_0000_0000_0000;
array[58091] <= 16'b0000_0000_0000_0000;
array[58092] <= 16'b0000_0000_0000_0000;
array[58093] <= 16'b0000_0000_0000_0000;
array[58094] <= 16'b0000_0000_0000_0000;
array[58095] <= 16'b0000_0000_0000_0000;
array[58096] <= 16'b0000_0000_0000_0000;
array[58097] <= 16'b0000_0000_0000_0000;
array[58098] <= 16'b0000_0000_0000_0000;
array[58099] <= 16'b0000_0000_0000_0000;
array[58100] <= 16'b0000_0000_0000_0000;
array[58101] <= 16'b0000_0000_0000_0000;
array[58102] <= 16'b0000_0000_0000_0000;
array[58103] <= 16'b0000_0000_0000_0000;
array[58104] <= 16'b0000_0000_0000_0000;
array[58105] <= 16'b0000_0000_0000_0000;
array[58106] <= 16'b0000_0000_0000_0000;
array[58107] <= 16'b0000_0000_0000_0000;
array[58108] <= 16'b0000_0000_0000_0000;
array[58109] <= 16'b0000_0000_0000_0000;
array[58110] <= 16'b0000_0000_0000_0000;
array[58111] <= 16'b0000_0000_0000_0000;
array[58112] <= 16'b0000_0000_0000_0000;
array[58113] <= 16'b0000_0000_0000_0000;
array[58114] <= 16'b0000_0000_0000_0000;
array[58115] <= 16'b0000_0000_0000_0000;
array[58116] <= 16'b0000_0000_0000_0000;
array[58117] <= 16'b0000_0000_0000_0000;
array[58118] <= 16'b0000_0000_0000_0000;
array[58119] <= 16'b0000_0000_0000_0000;
array[58120] <= 16'b0000_0000_0000_0000;
array[58121] <= 16'b0000_0000_0000_0000;
array[58122] <= 16'b0000_0000_0000_0000;
array[58123] <= 16'b0000_0000_0000_0000;
array[58124] <= 16'b0000_0000_0000_0000;
array[58125] <= 16'b0000_0000_0000_0000;
array[58126] <= 16'b0000_0000_0000_0000;
array[58127] <= 16'b0000_0000_0000_0000;
array[58128] <= 16'b0000_0000_0000_0000;
array[58129] <= 16'b0000_0000_0000_0000;
array[58130] <= 16'b0000_0000_0000_0000;
array[58131] <= 16'b0000_0000_0000_0000;
array[58132] <= 16'b0000_0000_0000_0000;
array[58133] <= 16'b0000_0000_0000_0000;
array[58134] <= 16'b0000_0000_0000_0000;
array[58135] <= 16'b0000_0000_0000_0000;
array[58136] <= 16'b0000_0000_0000_0000;
array[58137] <= 16'b0000_0000_0000_0000;
array[58138] <= 16'b0000_0000_0000_0000;
array[58139] <= 16'b0000_0000_0000_0000;
array[58140] <= 16'b0000_0000_0000_0000;
array[58141] <= 16'b0000_0000_0000_0000;
array[58142] <= 16'b0000_0000_0000_0000;
array[58143] <= 16'b0000_0000_0000_0000;
array[58144] <= 16'b0000_0000_0000_0000;
array[58145] <= 16'b0000_0000_0000_0000;
array[58146] <= 16'b0000_0000_0000_0000;
array[58147] <= 16'b0000_0000_0000_0000;
array[58148] <= 16'b0000_0000_0000_0000;
array[58149] <= 16'b0000_0000_0000_0000;
array[58150] <= 16'b0000_0000_0000_0000;
array[58151] <= 16'b0000_0000_0000_0000;
array[58152] <= 16'b0000_0000_0000_0000;
array[58153] <= 16'b0000_0000_0000_0000;
array[58154] <= 16'b0000_0000_0000_0000;
array[58155] <= 16'b0000_0000_0000_0000;
array[58156] <= 16'b0000_0000_0000_0000;
array[58157] <= 16'b0000_0000_0000_0000;
array[58158] <= 16'b0000_0000_0000_0000;
array[58159] <= 16'b0000_0000_0000_0000;
array[58160] <= 16'b0000_0000_0000_0000;
array[58161] <= 16'b0000_0000_0000_0000;
array[58162] <= 16'b0000_0000_0000_0000;
array[58163] <= 16'b0000_0000_0000_0000;
array[58164] <= 16'b0000_0000_0000_0000;
array[58165] <= 16'b0000_0000_0000_0000;
array[58166] <= 16'b0000_0000_0000_0000;
array[58167] <= 16'b0000_0000_0000_0000;
array[58168] <= 16'b0000_0000_0000_0000;
array[58169] <= 16'b0000_0000_0000_0000;
array[58170] <= 16'b0000_0000_0000_0000;
array[58171] <= 16'b0000_0000_0000_0000;
array[58172] <= 16'b0000_0000_0000_0000;
array[58173] <= 16'b0000_0000_0000_0000;
array[58174] <= 16'b0000_0000_0000_0000;
array[58175] <= 16'b0000_0000_0000_0000;
array[58176] <= 16'b0000_0000_0000_0000;
array[58177] <= 16'b0000_0000_0000_0000;
array[58178] <= 16'b0000_0000_0000_0000;
array[58179] <= 16'b0000_0000_0000_0000;
array[58180] <= 16'b0000_0000_0000_0000;
array[58181] <= 16'b0000_0000_0000_0000;
array[58182] <= 16'b0000_0000_0000_0000;
array[58183] <= 16'b0000_0000_0000_0000;
array[58184] <= 16'b0000_0000_0000_0000;
array[58185] <= 16'b0000_0000_0000_0000;
array[58186] <= 16'b0000_0000_0000_0000;
array[58187] <= 16'b0000_0000_0000_0000;
array[58188] <= 16'b0000_0000_0000_0000;
array[58189] <= 16'b0000_0000_0000_0000;
array[58190] <= 16'b0000_0000_0000_0000;
array[58191] <= 16'b0000_0000_0000_0000;
array[58192] <= 16'b0000_0000_0000_0000;
array[58193] <= 16'b0000_0000_0000_0000;
array[58194] <= 16'b0000_0000_0000_0000;
array[58195] <= 16'b0000_0000_0000_0000;
array[58196] <= 16'b0000_0000_0000_0000;
array[58197] <= 16'b0000_0000_0000_0000;
array[58198] <= 16'b0000_0000_0000_0000;
array[58199] <= 16'b0000_0000_0000_0000;
array[58200] <= 16'b0000_0000_0000_0000;
array[58201] <= 16'b0000_0000_0000_0000;
array[58202] <= 16'b0000_0000_0000_0000;
array[58203] <= 16'b0000_0000_0000_0000;
array[58204] <= 16'b0000_0000_0000_0000;
array[58205] <= 16'b0000_0000_0000_0000;
array[58206] <= 16'b0000_0000_0000_0000;
array[58207] <= 16'b0000_0000_0000_0000;
array[58208] <= 16'b0000_0000_0000_0000;
array[58209] <= 16'b0000_0000_0000_0000;
array[58210] <= 16'b0000_0000_0000_0000;
array[58211] <= 16'b0000_0000_0000_0000;
array[58212] <= 16'b0000_0000_0000_0000;
array[58213] <= 16'b0000_0000_0000_0000;
array[58214] <= 16'b0000_0000_0000_0000;
array[58215] <= 16'b0000_0000_0000_0000;
array[58216] <= 16'b0000_0000_0000_0000;
array[58217] <= 16'b0000_0000_0000_0000;
array[58218] <= 16'b0000_0000_0000_0000;
array[58219] <= 16'b0000_0000_0000_0000;
array[58220] <= 16'b0000_0000_0000_0000;
array[58221] <= 16'b0000_0000_0000_0000;
array[58222] <= 16'b0000_0000_0000_0000;
array[58223] <= 16'b0000_0000_0000_0000;
array[58224] <= 16'b0000_0000_0000_0000;
array[58225] <= 16'b0000_0000_0000_0000;
array[58226] <= 16'b0000_0000_0000_0000;
array[58227] <= 16'b0000_0000_0000_0000;
array[58228] <= 16'b0000_0000_0000_0000;
array[58229] <= 16'b0000_0000_0000_0000;
array[58230] <= 16'b0000_0000_0000_0000;
array[58231] <= 16'b0000_0000_0000_0000;
array[58232] <= 16'b0000_0000_0000_0000;
array[58233] <= 16'b0000_0000_0000_0000;
array[58234] <= 16'b0000_0000_0000_0000;
array[58235] <= 16'b0000_0000_0000_0000;
array[58236] <= 16'b0000_0000_0000_0000;
array[58237] <= 16'b0000_0000_0000_0000;
array[58238] <= 16'b0000_0000_0000_0000;
array[58239] <= 16'b0000_0000_0000_0000;
array[58240] <= 16'b0000_0000_0000_0000;
array[58241] <= 16'b0000_0000_0000_0000;
array[58242] <= 16'b0000_0000_0000_0000;
array[58243] <= 16'b0000_0000_0000_0000;
array[58244] <= 16'b0000_0000_0000_0000;
array[58245] <= 16'b0000_0000_0000_0000;
array[58246] <= 16'b0000_0000_0000_0000;
array[58247] <= 16'b0000_0000_0000_0000;
array[58248] <= 16'b0000_0000_0000_0000;
array[58249] <= 16'b0000_0000_0000_0000;
array[58250] <= 16'b0000_0000_0000_0000;
array[58251] <= 16'b0000_0000_0000_0000;
array[58252] <= 16'b0000_0000_0000_0000;
array[58253] <= 16'b0000_0000_0000_0000;
array[58254] <= 16'b0000_0000_0000_0000;
array[58255] <= 16'b0000_0000_0000_0000;
array[58256] <= 16'b0000_0000_0000_0000;
array[58257] <= 16'b0000_0000_0000_0000;
array[58258] <= 16'b0000_0000_0000_0000;
array[58259] <= 16'b0000_0000_0000_0000;
array[58260] <= 16'b0000_0000_0000_0000;
array[58261] <= 16'b0000_0000_0000_0000;
array[58262] <= 16'b0000_0000_0000_0000;
array[58263] <= 16'b0000_0000_0000_0000;
array[58264] <= 16'b0000_0000_0000_0000;
array[58265] <= 16'b0000_0000_0000_0000;
array[58266] <= 16'b0000_0000_0000_0000;
array[58267] <= 16'b0000_0000_0000_0000;
array[58268] <= 16'b0000_0000_0000_0000;
array[58269] <= 16'b0000_0000_0000_0000;
array[58270] <= 16'b0000_0000_0000_0000;
array[58271] <= 16'b0000_0000_0000_0000;
array[58272] <= 16'b0000_0000_0000_0000;
array[58273] <= 16'b0000_0000_0000_0000;
array[58274] <= 16'b0000_0000_0000_0000;
array[58275] <= 16'b0000_0000_0000_0000;
array[58276] <= 16'b0000_0000_0000_0000;
array[58277] <= 16'b0000_0000_0000_0000;
array[58278] <= 16'b0000_0000_0000_0000;
array[58279] <= 16'b0000_0000_0000_0000;
array[58280] <= 16'b0000_0000_0000_0000;
array[58281] <= 16'b0000_0000_0000_0000;
array[58282] <= 16'b0000_0000_0000_0000;
array[58283] <= 16'b0000_0000_0000_0000;
array[58284] <= 16'b0000_0000_0000_0000;
array[58285] <= 16'b0000_0000_0000_0000;
array[58286] <= 16'b0000_0000_0000_0000;
array[58287] <= 16'b0000_0000_0000_0000;
array[58288] <= 16'b0000_0000_0000_0000;
array[58289] <= 16'b0000_0000_0000_0000;
array[58290] <= 16'b0000_0000_0000_0000;
array[58291] <= 16'b0000_0000_0000_0000;
array[58292] <= 16'b0000_0000_0000_0000;
array[58293] <= 16'b0000_0000_0000_0000;
array[58294] <= 16'b0000_0000_0000_0000;
array[58295] <= 16'b0000_0000_0000_0000;
array[58296] <= 16'b0000_0000_0000_0000;
array[58297] <= 16'b0000_0000_0000_0000;
array[58298] <= 16'b0000_0000_0000_0000;
array[58299] <= 16'b0000_0000_0000_0000;
array[58300] <= 16'b0000_0000_0000_0000;
array[58301] <= 16'b0000_0000_0000_0000;
array[58302] <= 16'b0000_0000_0000_0000;
array[58303] <= 16'b0000_0000_0000_0000;
array[58304] <= 16'b0000_0000_0000_0000;
array[58305] <= 16'b0000_0000_0000_0000;
array[58306] <= 16'b0000_0000_0000_0000;
array[58307] <= 16'b0000_0000_0000_0000;
array[58308] <= 16'b0000_0000_0000_0000;
array[58309] <= 16'b0000_0000_0000_0000;
array[58310] <= 16'b0000_0000_0000_0000;
array[58311] <= 16'b0000_0000_0000_0000;
array[58312] <= 16'b0000_0000_0000_0000;
array[58313] <= 16'b0000_0000_0000_0000;
array[58314] <= 16'b0000_0000_0000_0000;
array[58315] <= 16'b0000_0000_0000_0000;
array[58316] <= 16'b0000_0000_0000_0000;
array[58317] <= 16'b0000_0000_0000_0000;
array[58318] <= 16'b0000_0000_0000_0000;
array[58319] <= 16'b0000_0000_0000_0000;
array[58320] <= 16'b0000_0000_0000_0000;
array[58321] <= 16'b0000_0000_0000_0000;
array[58322] <= 16'b0000_0000_0000_0000;
array[58323] <= 16'b0000_0000_0000_0000;
array[58324] <= 16'b0000_0000_0000_0000;
array[58325] <= 16'b0000_0000_0000_0000;
array[58326] <= 16'b0000_0000_0000_0000;
array[58327] <= 16'b0000_0000_0000_0000;
array[58328] <= 16'b0000_0000_0000_0000;
array[58329] <= 16'b0000_0000_0000_0000;
array[58330] <= 16'b0000_0000_0000_0000;
array[58331] <= 16'b0000_0000_0000_0000;
array[58332] <= 16'b0000_0000_0000_0000;
array[58333] <= 16'b0000_0000_0000_0000;
array[58334] <= 16'b0000_0000_0000_0000;
array[58335] <= 16'b0000_0000_0000_0000;
array[58336] <= 16'b0000_0000_0000_0000;
array[58337] <= 16'b0000_0000_0000_0000;
array[58338] <= 16'b0000_0000_0000_0000;
array[58339] <= 16'b0000_0000_0000_0000;
array[58340] <= 16'b0000_0000_0000_0000;
array[58341] <= 16'b0000_0000_0000_0000;
array[58342] <= 16'b0000_0000_0000_0000;
array[58343] <= 16'b0000_0000_0000_0000;
array[58344] <= 16'b0000_0000_0000_0000;
array[58345] <= 16'b0000_0000_0000_0000;
array[58346] <= 16'b0000_0000_0000_0000;
array[58347] <= 16'b0000_0000_0000_0000;
array[58348] <= 16'b0000_0000_0000_0000;
array[58349] <= 16'b0000_0000_0000_0000;
array[58350] <= 16'b0000_0000_0000_0000;
array[58351] <= 16'b0000_0000_0000_0000;
array[58352] <= 16'b0000_0000_0000_0000;
array[58353] <= 16'b0000_0000_0000_0000;
array[58354] <= 16'b0000_0000_0000_0000;
array[58355] <= 16'b0000_0000_0000_0000;
array[58356] <= 16'b0000_0000_0000_0000;
array[58357] <= 16'b0000_0000_0000_0000;
array[58358] <= 16'b0000_0000_0000_0000;
array[58359] <= 16'b0000_0000_0000_0000;
array[58360] <= 16'b0000_0000_0000_0000;
array[58361] <= 16'b0000_0000_0000_0000;
array[58362] <= 16'b0000_0000_0000_0000;
array[58363] <= 16'b0000_0000_0000_0000;
array[58364] <= 16'b0000_0000_0000_0000;
array[58365] <= 16'b0000_0000_0000_0000;
array[58366] <= 16'b0000_0000_0000_0000;
array[58367] <= 16'b0000_0000_0000_0000;
array[58368] <= 16'b0000_0000_0000_0000;
array[58369] <= 16'b0000_0000_0000_0000;
array[58370] <= 16'b0000_0000_0000_0000;
array[58371] <= 16'b0000_0000_0000_0000;
array[58372] <= 16'b0000_0000_0000_0000;
array[58373] <= 16'b0000_0000_0000_0000;
array[58374] <= 16'b0000_0000_0000_0000;
array[58375] <= 16'b0000_0000_0000_0000;
array[58376] <= 16'b0000_0000_0000_0000;
array[58377] <= 16'b0000_0000_0000_0000;
array[58378] <= 16'b0000_0000_0000_0000;
array[58379] <= 16'b0000_0000_0000_0000;
array[58380] <= 16'b0000_0000_0000_0000;
array[58381] <= 16'b0000_0000_0000_0000;
array[58382] <= 16'b0000_0000_0000_0000;
array[58383] <= 16'b0000_0000_0000_0000;
array[58384] <= 16'b0000_0000_0000_0000;
array[58385] <= 16'b0000_0000_0000_0000;
array[58386] <= 16'b0000_0000_0000_0000;
array[58387] <= 16'b0000_0000_0000_0000;
array[58388] <= 16'b0000_0000_0000_0000;
array[58389] <= 16'b0000_0000_0000_0000;
array[58390] <= 16'b0000_0000_0000_0000;
array[58391] <= 16'b0000_0000_0000_0000;
array[58392] <= 16'b0000_0000_0000_0000;
array[58393] <= 16'b0000_0000_0000_0000;
array[58394] <= 16'b0000_0000_0000_0000;
array[58395] <= 16'b0000_0000_0000_0000;
array[58396] <= 16'b0000_0000_0000_0000;
array[58397] <= 16'b0000_0000_0000_0000;
array[58398] <= 16'b0000_0000_0000_0000;
array[58399] <= 16'b0000_0000_0000_0000;
array[58400] <= 16'b0000_0000_0000_0000;
array[58401] <= 16'b0000_0000_0000_0000;
array[58402] <= 16'b0000_0000_0000_0000;
array[58403] <= 16'b0000_0000_0000_0000;
array[58404] <= 16'b0000_0000_0000_0000;
array[58405] <= 16'b0000_0000_0000_0000;
array[58406] <= 16'b0000_0000_0000_0000;
array[58407] <= 16'b0000_0000_0000_0000;
array[58408] <= 16'b0000_0000_0000_0000;
array[58409] <= 16'b0000_0000_0000_0000;
array[58410] <= 16'b0000_0000_0000_0000;
array[58411] <= 16'b0000_0000_0000_0000;
array[58412] <= 16'b0000_0000_0000_0000;
array[58413] <= 16'b0000_0000_0000_0000;
array[58414] <= 16'b0000_0000_0000_0000;
array[58415] <= 16'b0000_0000_0000_0000;
array[58416] <= 16'b0000_0000_0000_0000;
array[58417] <= 16'b0000_0000_0000_0000;
array[58418] <= 16'b0000_0000_0000_0000;
array[58419] <= 16'b0000_0000_0000_0000;
array[58420] <= 16'b0000_0000_0000_0000;
array[58421] <= 16'b0000_0000_0000_0000;
array[58422] <= 16'b0000_0000_0000_0000;
array[58423] <= 16'b0000_0000_0000_0000;
array[58424] <= 16'b0000_0000_0000_0000;
array[58425] <= 16'b0000_0000_0000_0000;
array[58426] <= 16'b0000_0000_0000_0000;
array[58427] <= 16'b0000_0000_0000_0000;
array[58428] <= 16'b0000_0000_0000_0000;
array[58429] <= 16'b0000_0000_0000_0000;
array[58430] <= 16'b0000_0000_0000_0000;
array[58431] <= 16'b0000_0000_0000_0000;
array[58432] <= 16'b0000_0000_0000_0000;
array[58433] <= 16'b0000_0000_0000_0000;
array[58434] <= 16'b0000_0000_0000_0000;
array[58435] <= 16'b0000_0000_0000_0000;
array[58436] <= 16'b0000_0000_0000_0000;
array[58437] <= 16'b0000_0000_0000_0000;
array[58438] <= 16'b0000_0000_0000_0000;
array[58439] <= 16'b0000_0000_0000_0000;
array[58440] <= 16'b0000_0000_0000_0000;
array[58441] <= 16'b0000_0000_0000_0000;
array[58442] <= 16'b0000_0000_0000_0000;
array[58443] <= 16'b0000_0000_0000_0000;
array[58444] <= 16'b0000_0000_0000_0000;
array[58445] <= 16'b0000_0000_0000_0000;
array[58446] <= 16'b0000_0000_0000_0000;
array[58447] <= 16'b0000_0000_0000_0000;
array[58448] <= 16'b0000_0000_0000_0000;
array[58449] <= 16'b0000_0000_0000_0000;
array[58450] <= 16'b0000_0000_0000_0000;
array[58451] <= 16'b0000_0000_0000_0000;
array[58452] <= 16'b0000_0000_0000_0000;
array[58453] <= 16'b0000_0000_0000_0000;
array[58454] <= 16'b0000_0000_0000_0000;
array[58455] <= 16'b0000_0000_0000_0000;
array[58456] <= 16'b0000_0000_0000_0000;
array[58457] <= 16'b0000_0000_0000_0000;
array[58458] <= 16'b0000_0000_0000_0000;
array[58459] <= 16'b0000_0000_0000_0000;
array[58460] <= 16'b0000_0000_0000_0000;
array[58461] <= 16'b0000_0000_0000_0000;
array[58462] <= 16'b0000_0000_0000_0000;
array[58463] <= 16'b0000_0000_0000_0000;
array[58464] <= 16'b0000_0000_0000_0000;
array[58465] <= 16'b0000_0000_0000_0000;
array[58466] <= 16'b0000_0000_0000_0000;
array[58467] <= 16'b0000_0000_0000_0000;
array[58468] <= 16'b0000_0000_0000_0000;
array[58469] <= 16'b0000_0000_0000_0000;
array[58470] <= 16'b0000_0000_0000_0000;
array[58471] <= 16'b0000_0000_0000_0000;
array[58472] <= 16'b0000_0000_0000_0000;
array[58473] <= 16'b0000_0000_0000_0000;
array[58474] <= 16'b0000_0000_0000_0000;
array[58475] <= 16'b0000_0000_0000_0000;
array[58476] <= 16'b0000_0000_0000_0000;
array[58477] <= 16'b0000_0000_0000_0000;
array[58478] <= 16'b0000_0000_0000_0000;
array[58479] <= 16'b0000_0000_0000_0000;
array[58480] <= 16'b0000_0000_0000_0000;
array[58481] <= 16'b0000_0000_0000_0000;
array[58482] <= 16'b0000_0000_0000_0000;
array[58483] <= 16'b0000_0000_0000_0000;
array[58484] <= 16'b0000_0000_0000_0000;
array[58485] <= 16'b0000_0000_0000_0000;
array[58486] <= 16'b0000_0000_0000_0000;
array[58487] <= 16'b0000_0000_0000_0000;
array[58488] <= 16'b0000_0000_0000_0000;
array[58489] <= 16'b0000_0000_0000_0000;
array[58490] <= 16'b0000_0000_0000_0000;
array[58491] <= 16'b0000_0000_0000_0000;
array[58492] <= 16'b0000_0000_0000_0000;
array[58493] <= 16'b0000_0000_0000_0000;
array[58494] <= 16'b0000_0000_0000_0000;
array[58495] <= 16'b0000_0000_0000_0000;
array[58496] <= 16'b0000_0000_0000_0000;
array[58497] <= 16'b0000_0000_0000_0000;
array[58498] <= 16'b0000_0000_0000_0000;
array[58499] <= 16'b0000_0000_0000_0000;
array[58500] <= 16'b0000_0000_0000_0000;
array[58501] <= 16'b0000_0000_0000_0000;
array[58502] <= 16'b0000_0000_0000_0000;
array[58503] <= 16'b0000_0000_0000_0000;
array[58504] <= 16'b0000_0000_0000_0000;
array[58505] <= 16'b0000_0000_0000_0000;
array[58506] <= 16'b0000_0000_0000_0000;
array[58507] <= 16'b0000_0000_0000_0000;
array[58508] <= 16'b0000_0000_0000_0000;
array[58509] <= 16'b0000_0000_0000_0000;
array[58510] <= 16'b0000_0000_0000_0000;
array[58511] <= 16'b0000_0000_0000_0000;
array[58512] <= 16'b0000_0000_0000_0000;
array[58513] <= 16'b0000_0000_0000_0000;
array[58514] <= 16'b0000_0000_0000_0000;
array[58515] <= 16'b0000_0000_0000_0000;
array[58516] <= 16'b0000_0000_0000_0000;
array[58517] <= 16'b0000_0000_0000_0000;
array[58518] <= 16'b0000_0000_0000_0000;
array[58519] <= 16'b0000_0000_0000_0000;
array[58520] <= 16'b0000_0000_0000_0000;
array[58521] <= 16'b0000_0000_0000_0000;
array[58522] <= 16'b0000_0000_0000_0000;
array[58523] <= 16'b0000_0000_0000_0000;
array[58524] <= 16'b0000_0000_0000_0000;
array[58525] <= 16'b0000_0000_0000_0000;
array[58526] <= 16'b0000_0000_0000_0000;
array[58527] <= 16'b0000_0000_0000_0000;
array[58528] <= 16'b0000_0000_0000_0000;
array[58529] <= 16'b0000_0000_0000_0000;
array[58530] <= 16'b0000_0000_0000_0000;
array[58531] <= 16'b0000_0000_0000_0000;
array[58532] <= 16'b0000_0000_0000_0000;
array[58533] <= 16'b0000_0000_0000_0000;
array[58534] <= 16'b0000_0000_0000_0000;
array[58535] <= 16'b0000_0000_0000_0000;
array[58536] <= 16'b0000_0000_0000_0000;
array[58537] <= 16'b0000_0000_0000_0000;
array[58538] <= 16'b0000_0000_0000_0000;
array[58539] <= 16'b0000_0000_0000_0000;
array[58540] <= 16'b0000_0000_0000_0000;
array[58541] <= 16'b0000_0000_0000_0000;
array[58542] <= 16'b0000_0000_0000_0000;
array[58543] <= 16'b0000_0000_0000_0000;
array[58544] <= 16'b0000_0000_0000_0000;
array[58545] <= 16'b0000_0000_0000_0000;
array[58546] <= 16'b0000_0000_0000_0000;
array[58547] <= 16'b0000_0000_0000_0000;
array[58548] <= 16'b0000_0000_0000_0000;
array[58549] <= 16'b0000_0000_0000_0000;
array[58550] <= 16'b0000_0000_0000_0000;
array[58551] <= 16'b0000_0000_0000_0000;
array[58552] <= 16'b0000_0000_0000_0000;
array[58553] <= 16'b0000_0000_0000_0000;
array[58554] <= 16'b0000_0000_0000_0000;
array[58555] <= 16'b0000_0000_0000_0000;
array[58556] <= 16'b0000_0000_0000_0000;
array[58557] <= 16'b0000_0000_0000_0000;
array[58558] <= 16'b0000_0000_0000_0000;
array[58559] <= 16'b0000_0000_0000_0000;
array[58560] <= 16'b0000_0000_0000_0000;
array[58561] <= 16'b0000_0000_0000_0000;
array[58562] <= 16'b0000_0000_0000_0000;
array[58563] <= 16'b0000_0000_0000_0000;
array[58564] <= 16'b0000_0000_0000_0000;
array[58565] <= 16'b0000_0000_0000_0000;
array[58566] <= 16'b0000_0000_0000_0000;
array[58567] <= 16'b0000_0000_0000_0000;
array[58568] <= 16'b0000_0000_0000_0000;
array[58569] <= 16'b0000_0000_0000_0000;
array[58570] <= 16'b0000_0000_0000_0000;
array[58571] <= 16'b0000_0000_0000_0000;
array[58572] <= 16'b0000_0000_0000_0000;
array[58573] <= 16'b0000_0000_0000_0000;
array[58574] <= 16'b0000_0000_0000_0000;
array[58575] <= 16'b0000_0000_0000_0000;
array[58576] <= 16'b0000_0000_0000_0000;
array[58577] <= 16'b0000_0000_0000_0000;
array[58578] <= 16'b0000_0000_0000_0000;
array[58579] <= 16'b0000_0000_0000_0000;
array[58580] <= 16'b0000_0000_0000_0000;
array[58581] <= 16'b0000_0000_0000_0000;
array[58582] <= 16'b0000_0000_0000_0000;
array[58583] <= 16'b0000_0000_0000_0000;
array[58584] <= 16'b0000_0000_0000_0000;
array[58585] <= 16'b0000_0000_0000_0000;
array[58586] <= 16'b0000_0000_0000_0000;
array[58587] <= 16'b0000_0000_0000_0000;
array[58588] <= 16'b0000_0000_0000_0000;
array[58589] <= 16'b0000_0000_0000_0000;
array[58590] <= 16'b0000_0000_0000_0000;
array[58591] <= 16'b0000_0000_0000_0000;
array[58592] <= 16'b0000_0000_0000_0000;
array[58593] <= 16'b0000_0000_0000_0000;
array[58594] <= 16'b0000_0000_0000_0000;
array[58595] <= 16'b0000_0000_0000_0000;
array[58596] <= 16'b0000_0000_0000_0000;
array[58597] <= 16'b0000_0000_0000_0000;
array[58598] <= 16'b0000_0000_0000_0000;
array[58599] <= 16'b0000_0000_0000_0000;
array[58600] <= 16'b0000_0000_0000_0000;
array[58601] <= 16'b0000_0000_0000_0000;
array[58602] <= 16'b0000_0000_0000_0000;
array[58603] <= 16'b0000_0000_0000_0000;
array[58604] <= 16'b0000_0000_0000_0000;
array[58605] <= 16'b0000_0000_0000_0000;
array[58606] <= 16'b0000_0000_0000_0000;
array[58607] <= 16'b0000_0000_0000_0000;
array[58608] <= 16'b0000_0000_0000_0000;
array[58609] <= 16'b0000_0000_0000_0000;
array[58610] <= 16'b0000_0000_0000_0000;
array[58611] <= 16'b0000_0000_0000_0000;
array[58612] <= 16'b0000_0000_0000_0000;
array[58613] <= 16'b0000_0000_0000_0000;
array[58614] <= 16'b0000_0000_0000_0000;
array[58615] <= 16'b0000_0000_0000_0000;
array[58616] <= 16'b0000_0000_0000_0000;
array[58617] <= 16'b0000_0000_0000_0000;
array[58618] <= 16'b0000_0000_0000_0000;
array[58619] <= 16'b0000_0000_0000_0000;
array[58620] <= 16'b0000_0000_0000_0000;
array[58621] <= 16'b0000_0000_0000_0000;
array[58622] <= 16'b0000_0000_0000_0000;
array[58623] <= 16'b0000_0000_0000_0000;
array[58624] <= 16'b0000_0000_0000_0000;
array[58625] <= 16'b0000_0000_0000_0000;
array[58626] <= 16'b0000_0000_0000_0000;
array[58627] <= 16'b0000_0000_0000_0000;
array[58628] <= 16'b0000_0000_0000_0000;
array[58629] <= 16'b0000_0000_0000_0000;
array[58630] <= 16'b0000_0000_0000_0000;
array[58631] <= 16'b0000_0000_0000_0000;
array[58632] <= 16'b0000_0000_0000_0000;
array[58633] <= 16'b0000_0000_0000_0000;
array[58634] <= 16'b0000_0000_0000_0000;
array[58635] <= 16'b0000_0000_0000_0000;
array[58636] <= 16'b0000_0000_0000_0000;
array[58637] <= 16'b0000_0000_0000_0000;
array[58638] <= 16'b0000_0000_0000_0000;
array[58639] <= 16'b0000_0000_0000_0000;
array[58640] <= 16'b0000_0000_0000_0000;
array[58641] <= 16'b0000_0000_0000_0000;
array[58642] <= 16'b0000_0000_0000_0000;
array[58643] <= 16'b0000_0000_0000_0000;
array[58644] <= 16'b0000_0000_0000_0000;
array[58645] <= 16'b0000_0000_0000_0000;
array[58646] <= 16'b0000_0000_0000_0000;
array[58647] <= 16'b0000_0000_0000_0000;
array[58648] <= 16'b0000_0000_0000_0000;
array[58649] <= 16'b0000_0000_0000_0000;
array[58650] <= 16'b0000_0000_0000_0000;
array[58651] <= 16'b0000_0000_0000_0000;
array[58652] <= 16'b0000_0000_0000_0000;
array[58653] <= 16'b0000_0000_0000_0000;
array[58654] <= 16'b0000_0000_0000_0000;
array[58655] <= 16'b0000_0000_0000_0000;
array[58656] <= 16'b0000_0000_0000_0000;
array[58657] <= 16'b0000_0000_0000_0000;
array[58658] <= 16'b0000_0000_0000_0000;
array[58659] <= 16'b0000_0000_0000_0000;
array[58660] <= 16'b0000_0000_0000_0000;
array[58661] <= 16'b0000_0000_0000_0000;
array[58662] <= 16'b0000_0000_0000_0000;
array[58663] <= 16'b0000_0000_0000_0000;
array[58664] <= 16'b0000_0000_0000_0000;
array[58665] <= 16'b0000_0000_0000_0000;
array[58666] <= 16'b0000_0000_0000_0000;
array[58667] <= 16'b0000_0000_0000_0000;
array[58668] <= 16'b0000_0000_0000_0000;
array[58669] <= 16'b0000_0000_0000_0000;
array[58670] <= 16'b0000_0000_0000_0000;
array[58671] <= 16'b0000_0000_0000_0000;
array[58672] <= 16'b0000_0000_0000_0000;
array[58673] <= 16'b0000_0000_0000_0000;
array[58674] <= 16'b0000_0000_0000_0000;
array[58675] <= 16'b0000_0000_0000_0000;
array[58676] <= 16'b0000_0000_0000_0000;
array[58677] <= 16'b0000_0000_0000_0000;
array[58678] <= 16'b0000_0000_0000_0000;
array[58679] <= 16'b0000_0000_0000_0000;
array[58680] <= 16'b0000_0000_0000_0000;
array[58681] <= 16'b0000_0000_0000_0000;
array[58682] <= 16'b0000_0000_0000_0000;
array[58683] <= 16'b0000_0000_0000_0000;
array[58684] <= 16'b0000_0000_0000_0000;
array[58685] <= 16'b0000_0000_0000_0000;
array[58686] <= 16'b0000_0000_0000_0000;
array[58687] <= 16'b0000_0000_0000_0000;
array[58688] <= 16'b0000_0000_0000_0000;
array[58689] <= 16'b0000_0000_0000_0000;
array[58690] <= 16'b0000_0000_0000_0000;
array[58691] <= 16'b0000_0000_0000_0000;
array[58692] <= 16'b0000_0000_0000_0000;
array[58693] <= 16'b0000_0000_0000_0000;
array[58694] <= 16'b0000_0000_0000_0000;
array[58695] <= 16'b0000_0000_0000_0000;
array[58696] <= 16'b0000_0000_0000_0000;
array[58697] <= 16'b0000_0000_0000_0000;
array[58698] <= 16'b0000_0000_0000_0000;
array[58699] <= 16'b0000_0000_0000_0000;
array[58700] <= 16'b0000_0000_0000_0000;
array[58701] <= 16'b0000_0000_0000_0000;
array[58702] <= 16'b0000_0000_0000_0000;
array[58703] <= 16'b0000_0000_0000_0000;
array[58704] <= 16'b0000_0000_0000_0000;
array[58705] <= 16'b0000_0000_0000_0000;
array[58706] <= 16'b0000_0000_0000_0000;
array[58707] <= 16'b0000_0000_0000_0000;
array[58708] <= 16'b0000_0000_0000_0000;
array[58709] <= 16'b0000_0000_0000_0000;
array[58710] <= 16'b0000_0000_0000_0000;
array[58711] <= 16'b0000_0000_0000_0000;
array[58712] <= 16'b0000_0000_0000_0000;
array[58713] <= 16'b0000_0000_0000_0000;
array[58714] <= 16'b0000_0000_0000_0000;
array[58715] <= 16'b0000_0000_0000_0000;
array[58716] <= 16'b0000_0000_0000_0000;
array[58717] <= 16'b0000_0000_0000_0000;
array[58718] <= 16'b0000_0000_0000_0000;
array[58719] <= 16'b0000_0000_0000_0000;
array[58720] <= 16'b0000_0000_0000_0000;
array[58721] <= 16'b0000_0000_0000_0000;
array[58722] <= 16'b0000_0000_0000_0000;
array[58723] <= 16'b0000_0000_0000_0000;
array[58724] <= 16'b0000_0000_0000_0000;
array[58725] <= 16'b0000_0000_0000_0000;
array[58726] <= 16'b0000_0000_0000_0000;
array[58727] <= 16'b0000_0000_0000_0000;
array[58728] <= 16'b0000_0000_0000_0000;
array[58729] <= 16'b0000_0000_0000_0000;
array[58730] <= 16'b0000_0000_0000_0000;
array[58731] <= 16'b0000_0000_0000_0000;
array[58732] <= 16'b0000_0000_0000_0000;
array[58733] <= 16'b0000_0000_0000_0000;
array[58734] <= 16'b0000_0000_0000_0000;
array[58735] <= 16'b0000_0000_0000_0000;
array[58736] <= 16'b0000_0000_0000_0000;
array[58737] <= 16'b0000_0000_0000_0000;
array[58738] <= 16'b0000_0000_0000_0000;
array[58739] <= 16'b0000_0000_0000_0000;
array[58740] <= 16'b0000_0000_0000_0000;
array[58741] <= 16'b0000_0000_0000_0000;
array[58742] <= 16'b0000_0000_0000_0000;
array[58743] <= 16'b0000_0000_0000_0000;
array[58744] <= 16'b0000_0000_0000_0000;
array[58745] <= 16'b0000_0000_0000_0000;
array[58746] <= 16'b0000_0000_0000_0000;
array[58747] <= 16'b0000_0000_0000_0000;
array[58748] <= 16'b0000_0000_0000_0000;
array[58749] <= 16'b0000_0000_0000_0000;
array[58750] <= 16'b0000_0000_0000_0000;
array[58751] <= 16'b0000_0000_0000_0000;
array[58752] <= 16'b0000_0000_0000_0000;
array[58753] <= 16'b0000_0000_0000_0000;
array[58754] <= 16'b0000_0000_0000_0000;
array[58755] <= 16'b0000_0000_0000_0000;
array[58756] <= 16'b0000_0000_0000_0000;
array[58757] <= 16'b0000_0000_0000_0000;
array[58758] <= 16'b0000_0000_0000_0000;
array[58759] <= 16'b0000_0000_0000_0000;
array[58760] <= 16'b0000_0000_0000_0000;
array[58761] <= 16'b0000_0000_0000_0000;
array[58762] <= 16'b0000_0000_0000_0000;
array[58763] <= 16'b0000_0000_0000_0000;
array[58764] <= 16'b0000_0000_0000_0000;
array[58765] <= 16'b0000_0000_0000_0000;
array[58766] <= 16'b0000_0000_0000_0000;
array[58767] <= 16'b0000_0000_0000_0000;
array[58768] <= 16'b0000_0000_0000_0000;
array[58769] <= 16'b0000_0000_0000_0000;
array[58770] <= 16'b0000_0000_0000_0000;
array[58771] <= 16'b0000_0000_0000_0000;
array[58772] <= 16'b0000_0000_0000_0000;
array[58773] <= 16'b0000_0000_0000_0000;
array[58774] <= 16'b0000_0000_0000_0000;
array[58775] <= 16'b0000_0000_0000_0000;
array[58776] <= 16'b0000_0000_0000_0000;
array[58777] <= 16'b0000_0000_0000_0000;
array[58778] <= 16'b0000_0000_0000_0000;
array[58779] <= 16'b0000_0000_0000_0000;
array[58780] <= 16'b0000_0000_0000_0000;
array[58781] <= 16'b0000_0000_0000_0000;
array[58782] <= 16'b0000_0000_0000_0000;
array[58783] <= 16'b0000_0000_0000_0000;
array[58784] <= 16'b0000_0000_0000_0000;
array[58785] <= 16'b0000_0000_0000_0000;
array[58786] <= 16'b0000_0000_0000_0000;
array[58787] <= 16'b0000_0000_0000_0000;
array[58788] <= 16'b0000_0000_0000_0000;
array[58789] <= 16'b0000_0000_0000_0000;
array[58790] <= 16'b0000_0000_0000_0000;
array[58791] <= 16'b0000_0000_0000_0000;
array[58792] <= 16'b0000_0000_0000_0000;
array[58793] <= 16'b0000_0000_0000_0000;
array[58794] <= 16'b0000_0000_0000_0000;
array[58795] <= 16'b0000_0000_0000_0000;
array[58796] <= 16'b0000_0000_0000_0000;
array[58797] <= 16'b0000_0000_0000_0000;
array[58798] <= 16'b0000_0000_0000_0000;
array[58799] <= 16'b0000_0000_0000_0000;
array[58800] <= 16'b0000_0000_0000_0000;
array[58801] <= 16'b0000_0000_0000_0000;
array[58802] <= 16'b0000_0000_0000_0000;
array[58803] <= 16'b0000_0000_0000_0000;
array[58804] <= 16'b0000_0000_0000_0000;
array[58805] <= 16'b0000_0000_0000_0000;
array[58806] <= 16'b0000_0000_0000_0000;
array[58807] <= 16'b0000_0000_0000_0000;
array[58808] <= 16'b0000_0000_0000_0000;
array[58809] <= 16'b0000_0000_0000_0000;
array[58810] <= 16'b0000_0000_0000_0000;
array[58811] <= 16'b0000_0000_0000_0000;
array[58812] <= 16'b0000_0000_0000_0000;
array[58813] <= 16'b0000_0000_0000_0000;
array[58814] <= 16'b0000_0000_0000_0000;
array[58815] <= 16'b0000_0000_0000_0000;
array[58816] <= 16'b0000_0000_0000_0000;
array[58817] <= 16'b0000_0000_0000_0000;
array[58818] <= 16'b0000_0000_0000_0000;
array[58819] <= 16'b0000_0000_0000_0000;
array[58820] <= 16'b0000_0000_0000_0000;
array[58821] <= 16'b0000_0000_0000_0000;
array[58822] <= 16'b0000_0000_0000_0000;
array[58823] <= 16'b0000_0000_0000_0000;
array[58824] <= 16'b0000_0000_0000_0000;
array[58825] <= 16'b0000_0000_0000_0000;
array[58826] <= 16'b0000_0000_0000_0000;
array[58827] <= 16'b0000_0000_0000_0000;
array[58828] <= 16'b0000_0000_0000_0000;
array[58829] <= 16'b0000_0000_0000_0000;
array[58830] <= 16'b0000_0000_0000_0000;
array[58831] <= 16'b0000_0000_0000_0000;
array[58832] <= 16'b0000_0000_0000_0000;
array[58833] <= 16'b0000_0000_0000_0000;
array[58834] <= 16'b0000_0000_0000_0000;
array[58835] <= 16'b0000_0000_0000_0000;
array[58836] <= 16'b0000_0000_0000_0000;
array[58837] <= 16'b0000_0000_0000_0000;
array[58838] <= 16'b0000_0000_0000_0000;
array[58839] <= 16'b0000_0000_0000_0000;
array[58840] <= 16'b0000_0000_0000_0000;
array[58841] <= 16'b0000_0000_0000_0000;
array[58842] <= 16'b0000_0000_0000_0000;
array[58843] <= 16'b0000_0000_0000_0000;
array[58844] <= 16'b0000_0000_0000_0000;
array[58845] <= 16'b0000_0000_0000_0000;
array[58846] <= 16'b0000_0000_0000_0000;
array[58847] <= 16'b0000_0000_0000_0000;
array[58848] <= 16'b0000_0000_0000_0000;
array[58849] <= 16'b0000_0000_0000_0000;
array[58850] <= 16'b0000_0000_0000_0000;
array[58851] <= 16'b0000_0000_0000_0000;
array[58852] <= 16'b0000_0000_0000_0000;
array[58853] <= 16'b0000_0000_0000_0000;
array[58854] <= 16'b0000_0000_0000_0000;
array[58855] <= 16'b0000_0000_0000_0000;
array[58856] <= 16'b0000_0000_0000_0000;
array[58857] <= 16'b0000_0000_0000_0000;
array[58858] <= 16'b0000_0000_0000_0000;
array[58859] <= 16'b0000_0000_0000_0000;
array[58860] <= 16'b0000_0000_0000_0000;
array[58861] <= 16'b0000_0000_0000_0000;
array[58862] <= 16'b0000_0000_0000_0000;
array[58863] <= 16'b0000_0000_0000_0000;
array[58864] <= 16'b0000_0000_0000_0000;
array[58865] <= 16'b0000_0000_0000_0000;
array[58866] <= 16'b0000_0000_0000_0000;
array[58867] <= 16'b0000_0000_0000_0000;
array[58868] <= 16'b0000_0000_0000_0000;
array[58869] <= 16'b0000_0000_0000_0000;
array[58870] <= 16'b0000_0000_0000_0000;
array[58871] <= 16'b0000_0000_0000_0000;
array[58872] <= 16'b0000_0000_0000_0000;
array[58873] <= 16'b0000_0000_0000_0000;
array[58874] <= 16'b0000_0000_0000_0000;
array[58875] <= 16'b0000_0000_0000_0000;
array[58876] <= 16'b0000_0000_0000_0000;
array[58877] <= 16'b0000_0000_0000_0000;
array[58878] <= 16'b0000_0000_0000_0000;
array[58879] <= 16'b0000_0000_0000_0000;
array[58880] <= 16'b0000_0000_0000_0000;
array[58881] <= 16'b0000_0000_0000_0000;
array[58882] <= 16'b0000_0000_0000_0000;
array[58883] <= 16'b0000_0000_0000_0000;
array[58884] <= 16'b0000_0000_0000_0000;
array[58885] <= 16'b0000_0000_0000_0000;
array[58886] <= 16'b0000_0000_0000_0000;
array[58887] <= 16'b0000_0000_0000_0000;
array[58888] <= 16'b0000_0000_0000_0000;
array[58889] <= 16'b0000_0000_0000_0000;
array[58890] <= 16'b0000_0000_0000_0000;
array[58891] <= 16'b0000_0000_0000_0000;
array[58892] <= 16'b0000_0000_0000_0000;
array[58893] <= 16'b0000_0000_0000_0000;
array[58894] <= 16'b0000_0000_0000_0000;
array[58895] <= 16'b0000_0000_0000_0000;
array[58896] <= 16'b0000_0000_0000_0000;
array[58897] <= 16'b0000_0000_0000_0000;
array[58898] <= 16'b0000_0000_0000_0000;
array[58899] <= 16'b0000_0000_0000_0000;
array[58900] <= 16'b0000_0000_0000_0000;
array[58901] <= 16'b0000_0000_0000_0000;
array[58902] <= 16'b0000_0000_0000_0000;
array[58903] <= 16'b0000_0000_0000_0000;
array[58904] <= 16'b0000_0000_0000_0000;
array[58905] <= 16'b0000_0000_0000_0000;
array[58906] <= 16'b0000_0000_0000_0000;
array[58907] <= 16'b0000_0000_0000_0000;
array[58908] <= 16'b0000_0000_0000_0000;
array[58909] <= 16'b0000_0000_0000_0000;
array[58910] <= 16'b0000_0000_0000_0000;
array[58911] <= 16'b0000_0000_0000_0000;
array[58912] <= 16'b0000_0000_0000_0000;
array[58913] <= 16'b0000_0000_0000_0000;
array[58914] <= 16'b0000_0000_0000_0000;
array[58915] <= 16'b0000_0000_0000_0000;
array[58916] <= 16'b0000_0000_0000_0000;
array[58917] <= 16'b0000_0000_0000_0000;
array[58918] <= 16'b0000_0000_0000_0000;
array[58919] <= 16'b0000_0000_0000_0000;
array[58920] <= 16'b0000_0000_0000_0000;
array[58921] <= 16'b0000_0000_0000_0000;
array[58922] <= 16'b0000_0000_0000_0000;
array[58923] <= 16'b0000_0000_0000_0000;
array[58924] <= 16'b0000_0000_0000_0000;
array[58925] <= 16'b0000_0000_0000_0000;
array[58926] <= 16'b0000_0000_0000_0000;
array[58927] <= 16'b0000_0000_0000_0000;
array[58928] <= 16'b0000_0000_0000_0000;
array[58929] <= 16'b0000_0000_0000_0000;
array[58930] <= 16'b0000_0000_0000_0000;
array[58931] <= 16'b0000_0000_0000_0000;
array[58932] <= 16'b0000_0000_0000_0000;
array[58933] <= 16'b0000_0000_0000_0000;
array[58934] <= 16'b0000_0000_0000_0000;
array[58935] <= 16'b0000_0000_0000_0000;
array[58936] <= 16'b0000_0000_0000_0000;
array[58937] <= 16'b0000_0000_0000_0000;
array[58938] <= 16'b0000_0000_0000_0000;
array[58939] <= 16'b0000_0000_0000_0000;
array[58940] <= 16'b0000_0000_0000_0000;
array[58941] <= 16'b0000_0000_0000_0000;
array[58942] <= 16'b0000_0000_0000_0000;
array[58943] <= 16'b0000_0000_0000_0000;
array[58944] <= 16'b0000_0000_0000_0000;
array[58945] <= 16'b0000_0000_0000_0000;
array[58946] <= 16'b0000_0000_0000_0000;
array[58947] <= 16'b0000_0000_0000_0000;
array[58948] <= 16'b0000_0000_0000_0000;
array[58949] <= 16'b0000_0000_0000_0000;
array[58950] <= 16'b0000_0000_0000_0000;
array[58951] <= 16'b0000_0000_0000_0000;
array[58952] <= 16'b0000_0000_0000_0000;
array[58953] <= 16'b0000_0000_0000_0000;
array[58954] <= 16'b0000_0000_0000_0000;
array[58955] <= 16'b0000_0000_0000_0000;
array[58956] <= 16'b0000_0000_0000_0000;
array[58957] <= 16'b0000_0000_0000_0000;
array[58958] <= 16'b0000_0000_0000_0000;
array[58959] <= 16'b0000_0000_0000_0000;
array[58960] <= 16'b0000_0000_0000_0000;
array[58961] <= 16'b0000_0000_0000_0000;
array[58962] <= 16'b0000_0000_0000_0000;
array[58963] <= 16'b0000_0000_0000_0000;
array[58964] <= 16'b0000_0000_0000_0000;
array[58965] <= 16'b0000_0000_0000_0000;
array[58966] <= 16'b0000_0000_0000_0000;
array[58967] <= 16'b0000_0000_0000_0000;
array[58968] <= 16'b0000_0000_0000_0000;
array[58969] <= 16'b0000_0000_0000_0000;
array[58970] <= 16'b0000_0000_0000_0000;
array[58971] <= 16'b0000_0000_0000_0000;
array[58972] <= 16'b0000_0000_0000_0000;
array[58973] <= 16'b0000_0000_0000_0000;
array[58974] <= 16'b0000_0000_0000_0000;
array[58975] <= 16'b0000_0000_0000_0000;
array[58976] <= 16'b0000_0000_0000_0000;
array[58977] <= 16'b0000_0000_0000_0000;
array[58978] <= 16'b0000_0000_0000_0000;
array[58979] <= 16'b0000_0000_0000_0000;
array[58980] <= 16'b0000_0000_0000_0000;
array[58981] <= 16'b0000_0000_0000_0000;
array[58982] <= 16'b0000_0000_0000_0000;
array[58983] <= 16'b0000_0000_0000_0000;
array[58984] <= 16'b0000_0000_0000_0000;
array[58985] <= 16'b0000_0000_0000_0000;
array[58986] <= 16'b0000_0000_0000_0000;
array[58987] <= 16'b0000_0000_0000_0000;
array[58988] <= 16'b0000_0000_0000_0000;
array[58989] <= 16'b0000_0000_0000_0000;
array[58990] <= 16'b0000_0000_0000_0000;
array[58991] <= 16'b0000_0000_0000_0000;
array[58992] <= 16'b0000_0000_0000_0000;
array[58993] <= 16'b0000_0000_0000_0000;
array[58994] <= 16'b0000_0000_0000_0000;
array[58995] <= 16'b0000_0000_0000_0000;
array[58996] <= 16'b0000_0000_0000_0000;
array[58997] <= 16'b0000_0000_0000_0000;
array[58998] <= 16'b0000_0000_0000_0000;
array[58999] <= 16'b0000_0000_0000_0000;
array[59000] <= 16'b0000_0000_0000_0000;
array[59001] <= 16'b0000_0000_0000_0000;
array[59002] <= 16'b0000_0000_0000_0000;
array[59003] <= 16'b0000_0000_0000_0000;
array[59004] <= 16'b0000_0000_0000_0000;
array[59005] <= 16'b0000_0000_0000_0000;
array[59006] <= 16'b0000_0000_0000_0000;
array[59007] <= 16'b0000_0000_0000_0000;
array[59008] <= 16'b0000_0000_0000_0000;
array[59009] <= 16'b0000_0000_0000_0000;
array[59010] <= 16'b0000_0000_0000_0000;
array[59011] <= 16'b0000_0000_0000_0000;
array[59012] <= 16'b0000_0000_0000_0000;
array[59013] <= 16'b0000_0000_0000_0000;
array[59014] <= 16'b0000_0000_0000_0000;
array[59015] <= 16'b0000_0000_0000_0000;
array[59016] <= 16'b0000_0000_0000_0000;
array[59017] <= 16'b0000_0000_0000_0000;
array[59018] <= 16'b0000_0000_0000_0000;
array[59019] <= 16'b0000_0000_0000_0000;
array[59020] <= 16'b0000_0000_0000_0000;
array[59021] <= 16'b0000_0000_0000_0000;
array[59022] <= 16'b0000_0000_0000_0000;
array[59023] <= 16'b0000_0000_0000_0000;
array[59024] <= 16'b0000_0000_0000_0000;
array[59025] <= 16'b0000_0000_0000_0000;
array[59026] <= 16'b0000_0000_0000_0000;
array[59027] <= 16'b0000_0000_0000_0000;
array[59028] <= 16'b0000_0000_0000_0000;
array[59029] <= 16'b0000_0000_0000_0000;
array[59030] <= 16'b0000_0000_0000_0000;
array[59031] <= 16'b0000_0000_0000_0000;
array[59032] <= 16'b0000_0000_0000_0000;
array[59033] <= 16'b0000_0000_0000_0000;
array[59034] <= 16'b0000_0000_0000_0000;
array[59035] <= 16'b0000_0000_0000_0000;
array[59036] <= 16'b0000_0000_0000_0000;
array[59037] <= 16'b0000_0000_0000_0000;
array[59038] <= 16'b0000_0000_0000_0000;
array[59039] <= 16'b0000_0000_0000_0000;
array[59040] <= 16'b0000_0000_0000_0000;
array[59041] <= 16'b0000_0000_0000_0000;
array[59042] <= 16'b0000_0000_0000_0000;
array[59043] <= 16'b0000_0000_0000_0000;
array[59044] <= 16'b0000_0000_0000_0000;
array[59045] <= 16'b0000_0000_0000_0000;
array[59046] <= 16'b0000_0000_0000_0000;
array[59047] <= 16'b0000_0000_0000_0000;
array[59048] <= 16'b0000_0000_0000_0000;
array[59049] <= 16'b0000_0000_0000_0000;
array[59050] <= 16'b0000_0000_0000_0000;
array[59051] <= 16'b0000_0000_0000_0000;
array[59052] <= 16'b0000_0000_0000_0000;
array[59053] <= 16'b0000_0000_0000_0000;
array[59054] <= 16'b0000_0000_0000_0000;
array[59055] <= 16'b0000_0000_0000_0000;
array[59056] <= 16'b0000_0000_0000_0000;
array[59057] <= 16'b0000_0000_0000_0000;
array[59058] <= 16'b0000_0000_0000_0000;
array[59059] <= 16'b0000_0000_0000_0000;
array[59060] <= 16'b0000_0000_0000_0000;
array[59061] <= 16'b0000_0000_0000_0000;
array[59062] <= 16'b0000_0000_0000_0000;
array[59063] <= 16'b0000_0000_0000_0000;
array[59064] <= 16'b0000_0000_0000_0000;
array[59065] <= 16'b0000_0000_0000_0000;
array[59066] <= 16'b0000_0000_0000_0000;
array[59067] <= 16'b0000_0000_0000_0000;
array[59068] <= 16'b0000_0000_0000_0000;
array[59069] <= 16'b0000_0000_0000_0000;
array[59070] <= 16'b0000_0000_0000_0000;
array[59071] <= 16'b0000_0000_0000_0000;
array[59072] <= 16'b0000_0000_0000_0000;
array[59073] <= 16'b0000_0000_0000_0000;
array[59074] <= 16'b0000_0000_0000_0000;
array[59075] <= 16'b0000_0000_0000_0000;
array[59076] <= 16'b0000_0000_0000_0000;
array[59077] <= 16'b0000_0000_0000_0000;
array[59078] <= 16'b0000_0000_0000_0000;
array[59079] <= 16'b0000_0000_0000_0000;
array[59080] <= 16'b0000_0000_0000_0000;
array[59081] <= 16'b0000_0000_0000_0000;
array[59082] <= 16'b0000_0000_0000_0000;
array[59083] <= 16'b0000_0000_0000_0000;
array[59084] <= 16'b0000_0000_0000_0000;
array[59085] <= 16'b0000_0000_0000_0000;
array[59086] <= 16'b0000_0000_0000_0000;
array[59087] <= 16'b0000_0000_0000_0000;
array[59088] <= 16'b0000_0000_0000_0000;
array[59089] <= 16'b0000_0000_0000_0000;
array[59090] <= 16'b0000_0000_0000_0000;
array[59091] <= 16'b0000_0000_0000_0000;
array[59092] <= 16'b0000_0000_0000_0000;
array[59093] <= 16'b0000_0000_0000_0000;
array[59094] <= 16'b0000_0000_0000_0000;
array[59095] <= 16'b0000_0000_0000_0000;
array[59096] <= 16'b0000_0000_0000_0000;
array[59097] <= 16'b0000_0000_0000_0000;
array[59098] <= 16'b0000_0000_0000_0000;
array[59099] <= 16'b0000_0000_0000_0000;
array[59100] <= 16'b0000_0000_0000_0000;
array[59101] <= 16'b0000_0000_0000_0000;
array[59102] <= 16'b0000_0000_0000_0000;
array[59103] <= 16'b0000_0000_0000_0000;
array[59104] <= 16'b0000_0000_0000_0000;
array[59105] <= 16'b0000_0000_0000_0000;
array[59106] <= 16'b0000_0000_0000_0000;
array[59107] <= 16'b0000_0000_0000_0000;
array[59108] <= 16'b0000_0000_0000_0000;
array[59109] <= 16'b0000_0000_0000_0000;
array[59110] <= 16'b0000_0000_0000_0000;
array[59111] <= 16'b0000_0000_0000_0000;
array[59112] <= 16'b0000_0000_0000_0000;
array[59113] <= 16'b0000_0000_0000_0000;
array[59114] <= 16'b0000_0000_0000_0000;
array[59115] <= 16'b0000_0000_0000_0000;
array[59116] <= 16'b0000_0000_0000_0000;
array[59117] <= 16'b0000_0000_0000_0000;
array[59118] <= 16'b0000_0000_0000_0000;
array[59119] <= 16'b0000_0000_0000_0000;
array[59120] <= 16'b0000_0000_0000_0000;
array[59121] <= 16'b0000_0000_0000_0000;
array[59122] <= 16'b0000_0000_0000_0000;
array[59123] <= 16'b0000_0000_0000_0000;
array[59124] <= 16'b0000_0000_0000_0000;
array[59125] <= 16'b0000_0000_0000_0000;
array[59126] <= 16'b0000_0000_0000_0000;
array[59127] <= 16'b0000_0000_0000_0000;
array[59128] <= 16'b0000_0000_0000_0000;
array[59129] <= 16'b0000_0000_0000_0000;
array[59130] <= 16'b0000_0000_0000_0000;
array[59131] <= 16'b0000_0000_0000_0000;
array[59132] <= 16'b0000_0000_0000_0000;
array[59133] <= 16'b0000_0000_0000_0000;
array[59134] <= 16'b0000_0000_0000_0000;
array[59135] <= 16'b0000_0000_0000_0000;
array[59136] <= 16'b0000_0000_0000_0000;
array[59137] <= 16'b0000_0000_0000_0000;
array[59138] <= 16'b0000_0000_0000_0000;
array[59139] <= 16'b0000_0000_0000_0000;
array[59140] <= 16'b0000_0000_0000_0000;
array[59141] <= 16'b0000_0000_0000_0000;
array[59142] <= 16'b0000_0000_0000_0000;
array[59143] <= 16'b0000_0000_0000_0000;
array[59144] <= 16'b0000_0000_0000_0000;
array[59145] <= 16'b0000_0000_0000_0000;
array[59146] <= 16'b0000_0000_0000_0000;
array[59147] <= 16'b0000_0000_0000_0000;
array[59148] <= 16'b0000_0000_0000_0000;
array[59149] <= 16'b0000_0000_0000_0000;
array[59150] <= 16'b0000_0000_0000_0000;
array[59151] <= 16'b0000_0000_0000_0000;
array[59152] <= 16'b0000_0000_0000_0000;
array[59153] <= 16'b0000_0000_0000_0000;
array[59154] <= 16'b0000_0000_0000_0000;
array[59155] <= 16'b0000_0000_0000_0000;
array[59156] <= 16'b0000_0000_0000_0000;
array[59157] <= 16'b0000_0000_0000_0000;
array[59158] <= 16'b0000_0000_0000_0000;
array[59159] <= 16'b0000_0000_0000_0000;
array[59160] <= 16'b0000_0000_0000_0000;
array[59161] <= 16'b0000_0000_0000_0000;
array[59162] <= 16'b0000_0000_0000_0000;
array[59163] <= 16'b0000_0000_0000_0000;
array[59164] <= 16'b0000_0000_0000_0000;
array[59165] <= 16'b0000_0000_0000_0000;
array[59166] <= 16'b0000_0000_0000_0000;
array[59167] <= 16'b0000_0000_0000_0000;
array[59168] <= 16'b0000_0000_0000_0000;
array[59169] <= 16'b0000_0000_0000_0000;
array[59170] <= 16'b0000_0000_0000_0000;
array[59171] <= 16'b0000_0000_0000_0000;
array[59172] <= 16'b0000_0000_0000_0000;
array[59173] <= 16'b0000_0000_0000_0000;
array[59174] <= 16'b0000_0000_0000_0000;
array[59175] <= 16'b0000_0000_0000_0000;
array[59176] <= 16'b0000_0000_0000_0000;
array[59177] <= 16'b0000_0000_0000_0000;
array[59178] <= 16'b0000_0000_0000_0000;
array[59179] <= 16'b0000_0000_0000_0000;
array[59180] <= 16'b0000_0000_0000_0000;
array[59181] <= 16'b0000_0000_0000_0000;
array[59182] <= 16'b0000_0000_0000_0000;
array[59183] <= 16'b0000_0000_0000_0000;
array[59184] <= 16'b0000_0000_0000_0000;
array[59185] <= 16'b0000_0000_0000_0000;
array[59186] <= 16'b0000_0000_0000_0000;
array[59187] <= 16'b0000_0000_0000_0000;
array[59188] <= 16'b0000_0000_0000_0000;
array[59189] <= 16'b0000_0000_0000_0000;
array[59190] <= 16'b0000_0000_0000_0000;
array[59191] <= 16'b0000_0000_0000_0000;
array[59192] <= 16'b0000_0000_0000_0000;
array[59193] <= 16'b0000_0000_0000_0000;
array[59194] <= 16'b0000_0000_0000_0000;
array[59195] <= 16'b0000_0000_0000_0000;
array[59196] <= 16'b0000_0000_0000_0000;
array[59197] <= 16'b0000_0000_0000_0000;
array[59198] <= 16'b0000_0000_0000_0000;
array[59199] <= 16'b0000_0000_0000_0000;
array[59200] <= 16'b0000_0000_0000_0000;
array[59201] <= 16'b0000_0000_0000_0000;
array[59202] <= 16'b0000_0000_0000_0000;
array[59203] <= 16'b0000_0000_0000_0000;
array[59204] <= 16'b0000_0000_0000_0000;
array[59205] <= 16'b0000_0000_0000_0000;
array[59206] <= 16'b0000_0000_0000_0000;
array[59207] <= 16'b0000_0000_0000_0000;
array[59208] <= 16'b0000_0000_0000_0000;
array[59209] <= 16'b0000_0000_0000_0000;
array[59210] <= 16'b0000_0000_0000_0000;
array[59211] <= 16'b0000_0000_0000_0000;
array[59212] <= 16'b0000_0000_0000_0000;
array[59213] <= 16'b0000_0000_0000_0000;
array[59214] <= 16'b0000_0000_0000_0000;
array[59215] <= 16'b0000_0000_0000_0000;
array[59216] <= 16'b0000_0000_0000_0000;
array[59217] <= 16'b0000_0000_0000_0000;
array[59218] <= 16'b0000_0000_0000_0000;
array[59219] <= 16'b0000_0000_0000_0000;
array[59220] <= 16'b0000_0000_0000_0000;
array[59221] <= 16'b0000_0000_0000_0000;
array[59222] <= 16'b0000_0000_0000_0000;
array[59223] <= 16'b0000_0000_0000_0000;
array[59224] <= 16'b0000_0000_0000_0000;
array[59225] <= 16'b0000_0000_0000_0000;
array[59226] <= 16'b0000_0000_0000_0000;
array[59227] <= 16'b0000_0000_0000_0000;
array[59228] <= 16'b0000_0000_0000_0000;
array[59229] <= 16'b0000_0000_0000_0000;
array[59230] <= 16'b0000_0000_0000_0000;
array[59231] <= 16'b0000_0000_0000_0000;
array[59232] <= 16'b0000_0000_0000_0000;
array[59233] <= 16'b0000_0000_0000_0000;
array[59234] <= 16'b0000_0000_0000_0000;
array[59235] <= 16'b0000_0000_0000_0000;
array[59236] <= 16'b0000_0000_0000_0000;
array[59237] <= 16'b0000_0000_0000_0000;
array[59238] <= 16'b0000_0000_0000_0000;
array[59239] <= 16'b0000_0000_0000_0000;
array[59240] <= 16'b0000_0000_0000_0000;
array[59241] <= 16'b0000_0000_0000_0000;
array[59242] <= 16'b0000_0000_0000_0000;
array[59243] <= 16'b0000_0000_0000_0000;
array[59244] <= 16'b0000_0000_0000_0000;
array[59245] <= 16'b0000_0000_0000_0000;
array[59246] <= 16'b0000_0000_0000_0000;
array[59247] <= 16'b0000_0000_0000_0000;
array[59248] <= 16'b0000_0000_0000_0000;
array[59249] <= 16'b0000_0000_0000_0000;
array[59250] <= 16'b0000_0000_0000_0000;
array[59251] <= 16'b0000_0000_0000_0000;
array[59252] <= 16'b0000_0000_0000_0000;
array[59253] <= 16'b0000_0000_0000_0000;
array[59254] <= 16'b0000_0000_0000_0000;
array[59255] <= 16'b0000_0000_0000_0000;
array[59256] <= 16'b0000_0000_0000_0000;
array[59257] <= 16'b0000_0000_0000_0000;
array[59258] <= 16'b0000_0000_0000_0000;
array[59259] <= 16'b0000_0000_0000_0000;
array[59260] <= 16'b0000_0000_0000_0000;
array[59261] <= 16'b0000_0000_0000_0000;
array[59262] <= 16'b0000_0000_0000_0000;
array[59263] <= 16'b0000_0000_0000_0000;
array[59264] <= 16'b0000_0000_0000_0000;
array[59265] <= 16'b0000_0000_0000_0000;
array[59266] <= 16'b0000_0000_0000_0000;
array[59267] <= 16'b0000_0000_0000_0000;
array[59268] <= 16'b0000_0000_0000_0000;
array[59269] <= 16'b0000_0000_0000_0000;
array[59270] <= 16'b0000_0000_0000_0000;
array[59271] <= 16'b0000_0000_0000_0000;
array[59272] <= 16'b0000_0000_0000_0000;
array[59273] <= 16'b0000_0000_0000_0000;
array[59274] <= 16'b0000_0000_0000_0000;
array[59275] <= 16'b0000_0000_0000_0000;
array[59276] <= 16'b0000_0000_0000_0000;
array[59277] <= 16'b0000_0000_0000_0000;
array[59278] <= 16'b0000_0000_0000_0000;
array[59279] <= 16'b0000_0000_0000_0000;
array[59280] <= 16'b0000_0000_0000_0000;
array[59281] <= 16'b0000_0000_0000_0000;
array[59282] <= 16'b0000_0000_0000_0000;
array[59283] <= 16'b0000_0000_0000_0000;
array[59284] <= 16'b0000_0000_0000_0000;
array[59285] <= 16'b0000_0000_0000_0000;
array[59286] <= 16'b0000_0000_0000_0000;
array[59287] <= 16'b0000_0000_0000_0000;
array[59288] <= 16'b0000_0000_0000_0000;
array[59289] <= 16'b0000_0000_0000_0000;
array[59290] <= 16'b0000_0000_0000_0000;
array[59291] <= 16'b0000_0000_0000_0000;
array[59292] <= 16'b0000_0000_0000_0000;
array[59293] <= 16'b0000_0000_0000_0000;
array[59294] <= 16'b0000_0000_0000_0000;
array[59295] <= 16'b0000_0000_0000_0000;
array[59296] <= 16'b0000_0000_0000_0000;
array[59297] <= 16'b0000_0000_0000_0000;
array[59298] <= 16'b0000_0000_0000_0000;
array[59299] <= 16'b0000_0000_0000_0000;
array[59300] <= 16'b0000_0000_0000_0000;
array[59301] <= 16'b0000_0000_0000_0000;
array[59302] <= 16'b0000_0000_0000_0000;
array[59303] <= 16'b0000_0000_0000_0000;
array[59304] <= 16'b0000_0000_0000_0000;
array[59305] <= 16'b0000_0000_0000_0000;
array[59306] <= 16'b0000_0000_0000_0000;
array[59307] <= 16'b0000_0000_0000_0000;
array[59308] <= 16'b0000_0000_0000_0000;
array[59309] <= 16'b0000_0000_0000_0000;
array[59310] <= 16'b0000_0000_0000_0000;
array[59311] <= 16'b0000_0000_0000_0000;
array[59312] <= 16'b0000_0000_0000_0000;
array[59313] <= 16'b0000_0000_0000_0000;
array[59314] <= 16'b0000_0000_0000_0000;
array[59315] <= 16'b0000_0000_0000_0000;
array[59316] <= 16'b0000_0000_0000_0000;
array[59317] <= 16'b0000_0000_0000_0000;
array[59318] <= 16'b0000_0000_0000_0000;
array[59319] <= 16'b0000_0000_0000_0000;
array[59320] <= 16'b0000_0000_0000_0000;
array[59321] <= 16'b0000_0000_0000_0000;
array[59322] <= 16'b0000_0000_0000_0000;
array[59323] <= 16'b0000_0000_0000_0000;
array[59324] <= 16'b0000_0000_0000_0000;
array[59325] <= 16'b0000_0000_0000_0000;
array[59326] <= 16'b0000_0000_0000_0000;
array[59327] <= 16'b0000_0000_0000_0000;
array[59328] <= 16'b0000_0000_0000_0000;
array[59329] <= 16'b0000_0000_0000_0000;
array[59330] <= 16'b0000_0000_0000_0000;
array[59331] <= 16'b0000_0000_0000_0000;
array[59332] <= 16'b0000_0000_0000_0000;
array[59333] <= 16'b0000_0000_0000_0000;
array[59334] <= 16'b0000_0000_0000_0000;
array[59335] <= 16'b0000_0000_0000_0000;
array[59336] <= 16'b0000_0000_0000_0000;
array[59337] <= 16'b0000_0000_0000_0000;
array[59338] <= 16'b0000_0000_0000_0000;
array[59339] <= 16'b0000_0000_0000_0000;
array[59340] <= 16'b0000_0000_0000_0000;
array[59341] <= 16'b0000_0000_0000_0000;
array[59342] <= 16'b0000_0000_0000_0000;
array[59343] <= 16'b0000_0000_0000_0000;
array[59344] <= 16'b0000_0000_0000_0000;
array[59345] <= 16'b0000_0000_0000_0000;
array[59346] <= 16'b0000_0000_0000_0000;
array[59347] <= 16'b0000_0000_0000_0000;
array[59348] <= 16'b0000_0000_0000_0000;
array[59349] <= 16'b0000_0000_0000_0000;
array[59350] <= 16'b0000_0000_0000_0000;
array[59351] <= 16'b0000_0000_0000_0000;
array[59352] <= 16'b0000_0000_0000_0000;
array[59353] <= 16'b0000_0000_0000_0000;
array[59354] <= 16'b0000_0000_0000_0000;
array[59355] <= 16'b0000_0000_0000_0000;
array[59356] <= 16'b0000_0000_0000_0000;
array[59357] <= 16'b0000_0000_0000_0000;
array[59358] <= 16'b0000_0000_0000_0000;
array[59359] <= 16'b0000_0000_0000_0000;
array[59360] <= 16'b0000_0000_0000_0000;
array[59361] <= 16'b0000_0000_0000_0000;
array[59362] <= 16'b0000_0000_0000_0000;
array[59363] <= 16'b0000_0000_0000_0000;
array[59364] <= 16'b0000_0000_0000_0000;
array[59365] <= 16'b0000_0000_0000_0000;
array[59366] <= 16'b0000_0000_0000_0000;
array[59367] <= 16'b0000_0000_0000_0000;
array[59368] <= 16'b0000_0000_0000_0000;
array[59369] <= 16'b0000_0000_0000_0000;
array[59370] <= 16'b0000_0000_0000_0000;
array[59371] <= 16'b0000_0000_0000_0000;
array[59372] <= 16'b0000_0000_0000_0000;
array[59373] <= 16'b0000_0000_0000_0000;
array[59374] <= 16'b0000_0000_0000_0000;
array[59375] <= 16'b0000_0000_0000_0000;
array[59376] <= 16'b0000_0000_0000_0000;
array[59377] <= 16'b0000_0000_0000_0000;
array[59378] <= 16'b0000_0000_0000_0000;
array[59379] <= 16'b0000_0000_0000_0000;
array[59380] <= 16'b0000_0000_0000_0000;
array[59381] <= 16'b0000_0000_0000_0000;
array[59382] <= 16'b0000_0000_0000_0000;
array[59383] <= 16'b0000_0000_0000_0000;
array[59384] <= 16'b0000_0000_0000_0000;
array[59385] <= 16'b0000_0000_0000_0000;
array[59386] <= 16'b0000_0000_0000_0000;
array[59387] <= 16'b0000_0000_0000_0000;
array[59388] <= 16'b0000_0000_0000_0000;
array[59389] <= 16'b0000_0000_0000_0000;
array[59390] <= 16'b0000_0000_0000_0000;
array[59391] <= 16'b0000_0000_0000_0000;
array[59392] <= 16'b0000_0000_0000_0000;
array[59393] <= 16'b0000_0000_0000_0000;
array[59394] <= 16'b0000_0000_0000_0000;
array[59395] <= 16'b0000_0000_0000_0000;
array[59396] <= 16'b0000_0000_0000_0000;
array[59397] <= 16'b0000_0000_0000_0000;
array[59398] <= 16'b0000_0000_0000_0000;
array[59399] <= 16'b0000_0000_0000_0000;
array[59400] <= 16'b0000_0000_0000_0000;
array[59401] <= 16'b0000_0000_0000_0000;
array[59402] <= 16'b0000_0000_0000_0000;
array[59403] <= 16'b0000_0000_0000_0000;
array[59404] <= 16'b0000_0000_0000_0000;
array[59405] <= 16'b0000_0000_0000_0000;
array[59406] <= 16'b0000_0000_0000_0000;
array[59407] <= 16'b0000_0000_0000_0000;
array[59408] <= 16'b0000_0000_0000_0000;
array[59409] <= 16'b0000_0000_0000_0000;
array[59410] <= 16'b0000_0000_0000_0000;
array[59411] <= 16'b0000_0000_0000_0000;
array[59412] <= 16'b0000_0000_0000_0000;
array[59413] <= 16'b0000_0000_0000_0000;
array[59414] <= 16'b0000_0000_0000_0000;
array[59415] <= 16'b0000_0000_0000_0000;
array[59416] <= 16'b0000_0000_0000_0000;
array[59417] <= 16'b0000_0000_0000_0000;
array[59418] <= 16'b0000_0000_0000_0000;
array[59419] <= 16'b0000_0000_0000_0000;
array[59420] <= 16'b0000_0000_0000_0000;
array[59421] <= 16'b0000_0000_0000_0000;
array[59422] <= 16'b0000_0000_0000_0000;
array[59423] <= 16'b0000_0000_0000_0000;
array[59424] <= 16'b0000_0000_0000_0000;
array[59425] <= 16'b0000_0000_0000_0000;
array[59426] <= 16'b0000_0000_0000_0000;
array[59427] <= 16'b0000_0000_0000_0000;
array[59428] <= 16'b0000_0000_0000_0000;
array[59429] <= 16'b0000_0000_0000_0000;
array[59430] <= 16'b0000_0000_0000_0000;
array[59431] <= 16'b0000_0000_0000_0000;
array[59432] <= 16'b0000_0000_0000_0000;
array[59433] <= 16'b0000_0000_0000_0000;
array[59434] <= 16'b0000_0000_0000_0000;
array[59435] <= 16'b0000_0000_0000_0000;
array[59436] <= 16'b0000_0000_0000_0000;
array[59437] <= 16'b0000_0000_0000_0000;
array[59438] <= 16'b0000_0000_0000_0000;
array[59439] <= 16'b0000_0000_0000_0000;
array[59440] <= 16'b0000_0000_0000_0000;
array[59441] <= 16'b0000_0000_0000_0000;
array[59442] <= 16'b0000_0000_0000_0000;
array[59443] <= 16'b0000_0000_0000_0000;
array[59444] <= 16'b0000_0000_0000_0000;
array[59445] <= 16'b0000_0000_0000_0000;
array[59446] <= 16'b0000_0000_0000_0000;
array[59447] <= 16'b0000_0000_0000_0000;
array[59448] <= 16'b0000_0000_0000_0000;
array[59449] <= 16'b0000_0000_0000_0000;
array[59450] <= 16'b0000_0000_0000_0000;
array[59451] <= 16'b0000_0000_0000_0000;
array[59452] <= 16'b0000_0000_0000_0000;
array[59453] <= 16'b0000_0000_0000_0000;
array[59454] <= 16'b0000_0000_0000_0000;
array[59455] <= 16'b0000_0000_0000_0000;
array[59456] <= 16'b0000_0000_0000_0000;
array[59457] <= 16'b0000_0000_0000_0000;
array[59458] <= 16'b0000_0000_0000_0000;
array[59459] <= 16'b0000_0000_0000_0000;
array[59460] <= 16'b0000_0000_0000_0000;
array[59461] <= 16'b0000_0000_0000_0000;
array[59462] <= 16'b0000_0000_0000_0000;
array[59463] <= 16'b0000_0000_0000_0000;
array[59464] <= 16'b0000_0000_0000_0000;
array[59465] <= 16'b0000_0000_0000_0000;
array[59466] <= 16'b0000_0000_0000_0000;
array[59467] <= 16'b0000_0000_0000_0000;
array[59468] <= 16'b0000_0000_0000_0000;
array[59469] <= 16'b0000_0000_0000_0000;
array[59470] <= 16'b0000_0000_0000_0000;
array[59471] <= 16'b0000_0000_0000_0000;
array[59472] <= 16'b0000_0000_0000_0000;
array[59473] <= 16'b0000_0000_0000_0000;
array[59474] <= 16'b0000_0000_0000_0000;
array[59475] <= 16'b0000_0000_0000_0000;
array[59476] <= 16'b0000_0000_0000_0000;
array[59477] <= 16'b0000_0000_0000_0000;
array[59478] <= 16'b0000_0000_0000_0000;
array[59479] <= 16'b0000_0000_0000_0000;
array[59480] <= 16'b0000_0000_0000_0000;
array[59481] <= 16'b0000_0000_0000_0000;
array[59482] <= 16'b0000_0000_0000_0000;
array[59483] <= 16'b0000_0000_0000_0000;
array[59484] <= 16'b0000_0000_0000_0000;
array[59485] <= 16'b0000_0000_0000_0000;
array[59486] <= 16'b0000_0000_0000_0000;
array[59487] <= 16'b0000_0000_0000_0000;
array[59488] <= 16'b0000_0000_0000_0000;
array[59489] <= 16'b0000_0000_0000_0000;
array[59490] <= 16'b0000_0000_0000_0000;
array[59491] <= 16'b0000_0000_0000_0000;
array[59492] <= 16'b0000_0000_0000_0000;
array[59493] <= 16'b0000_0000_0000_0000;
array[59494] <= 16'b0000_0000_0000_0000;
array[59495] <= 16'b0000_0000_0000_0000;
array[59496] <= 16'b0000_0000_0000_0000;
array[59497] <= 16'b0000_0000_0000_0000;
array[59498] <= 16'b0000_0000_0000_0000;
array[59499] <= 16'b0000_0000_0000_0000;
array[59500] <= 16'b0000_0000_0000_0000;
array[59501] <= 16'b0000_0000_0000_0000;
array[59502] <= 16'b0000_0000_0000_0000;
array[59503] <= 16'b0000_0000_0000_0000;
array[59504] <= 16'b0000_0000_0000_0000;
array[59505] <= 16'b0000_0000_0000_0000;
array[59506] <= 16'b0000_0000_0000_0000;
array[59507] <= 16'b0000_0000_0000_0000;
array[59508] <= 16'b0000_0000_0000_0000;
array[59509] <= 16'b0000_0000_0000_0000;
array[59510] <= 16'b0000_0000_0000_0000;
array[59511] <= 16'b0000_0000_0000_0000;
array[59512] <= 16'b0000_0000_0000_0000;
array[59513] <= 16'b0000_0000_0000_0000;
array[59514] <= 16'b0000_0000_0000_0000;
array[59515] <= 16'b0000_0000_0000_0000;
array[59516] <= 16'b0000_0000_0000_0000;
array[59517] <= 16'b0000_0000_0000_0000;
array[59518] <= 16'b0000_0000_0000_0000;
array[59519] <= 16'b0000_0000_0000_0000;
array[59520] <= 16'b0000_0000_0000_0000;
array[59521] <= 16'b0000_0000_0000_0000;
array[59522] <= 16'b0000_0000_0000_0000;
array[59523] <= 16'b0000_0000_0000_0000;
array[59524] <= 16'b0000_0000_0000_0000;
array[59525] <= 16'b0000_0000_0000_0000;
array[59526] <= 16'b0000_0000_0000_0000;
array[59527] <= 16'b0000_0000_0000_0000;
array[59528] <= 16'b0000_0000_0000_0000;
array[59529] <= 16'b0000_0000_0000_0000;
array[59530] <= 16'b0000_0000_0000_0000;
array[59531] <= 16'b0000_0000_0000_0000;
array[59532] <= 16'b0000_0000_0000_0000;
array[59533] <= 16'b0000_0000_0000_0000;
array[59534] <= 16'b0000_0000_0000_0000;
array[59535] <= 16'b0000_0000_0000_0000;
array[59536] <= 16'b0000_0000_0000_0000;
array[59537] <= 16'b0000_0000_0000_0000;
array[59538] <= 16'b0000_0000_0000_0000;
array[59539] <= 16'b0000_0000_0000_0000;
array[59540] <= 16'b0000_0000_0000_0000;
array[59541] <= 16'b0000_0000_0000_0000;
array[59542] <= 16'b0000_0000_0000_0000;
array[59543] <= 16'b0000_0000_0000_0000;
array[59544] <= 16'b0000_0000_0000_0000;
array[59545] <= 16'b0000_0000_0000_0000;
array[59546] <= 16'b0000_0000_0000_0000;
array[59547] <= 16'b0000_0000_0000_0000;
array[59548] <= 16'b0000_0000_0000_0000;
array[59549] <= 16'b0000_0000_0000_0000;
array[59550] <= 16'b0000_0000_0000_0000;
array[59551] <= 16'b0000_0000_0000_0000;
array[59552] <= 16'b0000_0000_0000_0000;
array[59553] <= 16'b0000_0000_0000_0000;
array[59554] <= 16'b0000_0000_0000_0000;
array[59555] <= 16'b0000_0000_0000_0000;
array[59556] <= 16'b0000_0000_0000_0000;
array[59557] <= 16'b0000_0000_0000_0000;
array[59558] <= 16'b0000_0000_0000_0000;
array[59559] <= 16'b0000_0000_0000_0000;
array[59560] <= 16'b0000_0000_0000_0000;
array[59561] <= 16'b0000_0000_0000_0000;
array[59562] <= 16'b0000_0000_0000_0000;
array[59563] <= 16'b0000_0000_0000_0000;
array[59564] <= 16'b0000_0000_0000_0000;
array[59565] <= 16'b0000_0000_0000_0000;
array[59566] <= 16'b0000_0000_0000_0000;
array[59567] <= 16'b0000_0000_0000_0000;
array[59568] <= 16'b0000_0000_0000_0000;
array[59569] <= 16'b0000_0000_0000_0000;
array[59570] <= 16'b0000_0000_0000_0000;
array[59571] <= 16'b0000_0000_0000_0000;
array[59572] <= 16'b0000_0000_0000_0000;
array[59573] <= 16'b0000_0000_0000_0000;
array[59574] <= 16'b0000_0000_0000_0000;
array[59575] <= 16'b0000_0000_0000_0000;
array[59576] <= 16'b0000_0000_0000_0000;
array[59577] <= 16'b0000_0000_0000_0000;
array[59578] <= 16'b0000_0000_0000_0000;
array[59579] <= 16'b0000_0000_0000_0000;
array[59580] <= 16'b0000_0000_0000_0000;
array[59581] <= 16'b0000_0000_0000_0000;
array[59582] <= 16'b0000_0000_0000_0000;
array[59583] <= 16'b0000_0000_0000_0000;
array[59584] <= 16'b0000_0000_0000_0000;
array[59585] <= 16'b0000_0000_0000_0000;
array[59586] <= 16'b0000_0000_0000_0000;
array[59587] <= 16'b0000_0000_0000_0000;
array[59588] <= 16'b0000_0000_0000_0000;
array[59589] <= 16'b0000_0000_0000_0000;
array[59590] <= 16'b0000_0000_0000_0000;
array[59591] <= 16'b0000_0000_0000_0000;
array[59592] <= 16'b0000_0000_0000_0000;
array[59593] <= 16'b0000_0000_0000_0000;
array[59594] <= 16'b0000_0000_0000_0000;
array[59595] <= 16'b0000_0000_0000_0000;
array[59596] <= 16'b0000_0000_0000_0000;
array[59597] <= 16'b0000_0000_0000_0000;
array[59598] <= 16'b0000_0000_0000_0000;
array[59599] <= 16'b0000_0000_0000_0000;
array[59600] <= 16'b0000_0000_0000_0000;
array[59601] <= 16'b0000_0000_0000_0000;
array[59602] <= 16'b0000_0000_0000_0000;
array[59603] <= 16'b0000_0000_0000_0000;
array[59604] <= 16'b0000_0000_0000_0000;
array[59605] <= 16'b0000_0000_0000_0000;
array[59606] <= 16'b0000_0000_0000_0000;
array[59607] <= 16'b0000_0000_0000_0000;
array[59608] <= 16'b0000_0000_0000_0000;
array[59609] <= 16'b0000_0000_0000_0000;
array[59610] <= 16'b0000_0000_0000_0000;
array[59611] <= 16'b0000_0000_0000_0000;
array[59612] <= 16'b0000_0000_0000_0000;
array[59613] <= 16'b0000_0000_0000_0000;
array[59614] <= 16'b0000_0000_0000_0000;
array[59615] <= 16'b0000_0000_0000_0000;
array[59616] <= 16'b0000_0000_0000_0000;
array[59617] <= 16'b0000_0000_0000_0000;
array[59618] <= 16'b0000_0000_0000_0000;
array[59619] <= 16'b0000_0000_0000_0000;
array[59620] <= 16'b0000_0000_0000_0000;
array[59621] <= 16'b0000_0000_0000_0000;
array[59622] <= 16'b0000_0000_0000_0000;
array[59623] <= 16'b0000_0000_0000_0000;
array[59624] <= 16'b0000_0000_0000_0000;
array[59625] <= 16'b0000_0000_0000_0000;
array[59626] <= 16'b0000_0000_0000_0000;
array[59627] <= 16'b0000_0000_0000_0000;
array[59628] <= 16'b0000_0000_0000_0000;
array[59629] <= 16'b0000_0000_0000_0000;
array[59630] <= 16'b0000_0000_0000_0000;
array[59631] <= 16'b0000_0000_0000_0000;
array[59632] <= 16'b0000_0000_0000_0000;
array[59633] <= 16'b0000_0000_0000_0000;
array[59634] <= 16'b0000_0000_0000_0000;
array[59635] <= 16'b0000_0000_0000_0000;
array[59636] <= 16'b0000_0000_0000_0000;
array[59637] <= 16'b0000_0000_0000_0000;
array[59638] <= 16'b0000_0000_0000_0000;
array[59639] <= 16'b0000_0000_0000_0000;
array[59640] <= 16'b0000_0000_0000_0000;
array[59641] <= 16'b0000_0000_0000_0000;
array[59642] <= 16'b0000_0000_0000_0000;
array[59643] <= 16'b0000_0000_0000_0000;
array[59644] <= 16'b0000_0000_0000_0000;
array[59645] <= 16'b0000_0000_0000_0000;
array[59646] <= 16'b0000_0000_0000_0000;
array[59647] <= 16'b0000_0000_0000_0000;
array[59648] <= 16'b0000_0000_0000_0000;
array[59649] <= 16'b0000_0000_0000_0000;
array[59650] <= 16'b0000_0000_0000_0000;
array[59651] <= 16'b0000_0000_0000_0000;
array[59652] <= 16'b0000_0000_0000_0000;
array[59653] <= 16'b0000_0000_0000_0000;
array[59654] <= 16'b0000_0000_0000_0000;
array[59655] <= 16'b0000_0000_0000_0000;
array[59656] <= 16'b0000_0000_0000_0000;
array[59657] <= 16'b0000_0000_0000_0000;
array[59658] <= 16'b0000_0000_0000_0000;
array[59659] <= 16'b0000_0000_0000_0000;
array[59660] <= 16'b0000_0000_0000_0000;
array[59661] <= 16'b0000_0000_0000_0000;
array[59662] <= 16'b0000_0000_0000_0000;
array[59663] <= 16'b0000_0000_0000_0000;
array[59664] <= 16'b0000_0000_0000_0000;
array[59665] <= 16'b0000_0000_0000_0000;
array[59666] <= 16'b0000_0000_0000_0000;
array[59667] <= 16'b0000_0000_0000_0000;
array[59668] <= 16'b0000_0000_0000_0000;
array[59669] <= 16'b0000_0000_0000_0000;
array[59670] <= 16'b0000_0000_0000_0000;
array[59671] <= 16'b0000_0000_0000_0000;
array[59672] <= 16'b0000_0000_0000_0000;
array[59673] <= 16'b0000_0000_0000_0000;
array[59674] <= 16'b0000_0000_0000_0000;
array[59675] <= 16'b0000_0000_0000_0000;
array[59676] <= 16'b0000_0000_0000_0000;
array[59677] <= 16'b0000_0000_0000_0000;
array[59678] <= 16'b0000_0000_0000_0000;
array[59679] <= 16'b0000_0000_0000_0000;
array[59680] <= 16'b0000_0000_0000_0000;
array[59681] <= 16'b0000_0000_0000_0000;
array[59682] <= 16'b0000_0000_0000_0000;
array[59683] <= 16'b0000_0000_0000_0000;
array[59684] <= 16'b0000_0000_0000_0000;
array[59685] <= 16'b0000_0000_0000_0000;
array[59686] <= 16'b0000_0000_0000_0000;
array[59687] <= 16'b0000_0000_0000_0000;
array[59688] <= 16'b0000_0000_0000_0000;
array[59689] <= 16'b0000_0000_0000_0000;
array[59690] <= 16'b0000_0000_0000_0000;
array[59691] <= 16'b0000_0000_0000_0000;
array[59692] <= 16'b0000_0000_0000_0000;
array[59693] <= 16'b0000_0000_0000_0000;
array[59694] <= 16'b0000_0000_0000_0000;
array[59695] <= 16'b0000_0000_0000_0000;
array[59696] <= 16'b0000_0000_0000_0000;
array[59697] <= 16'b0000_0000_0000_0000;
array[59698] <= 16'b0000_0000_0000_0000;
array[59699] <= 16'b0000_0000_0000_0000;
array[59700] <= 16'b0000_0000_0000_0000;
array[59701] <= 16'b0000_0000_0000_0000;
array[59702] <= 16'b0000_0000_0000_0000;
array[59703] <= 16'b0000_0000_0000_0000;
array[59704] <= 16'b0000_0000_0000_0000;
array[59705] <= 16'b0000_0000_0000_0000;
array[59706] <= 16'b0000_0000_0000_0000;
array[59707] <= 16'b0000_0000_0000_0000;
array[59708] <= 16'b0000_0000_0000_0000;
array[59709] <= 16'b0000_0000_0000_0000;
array[59710] <= 16'b0000_0000_0000_0000;
array[59711] <= 16'b0000_0000_0000_0000;
array[59712] <= 16'b0000_0000_0000_0000;
array[59713] <= 16'b0000_0000_0000_0000;
array[59714] <= 16'b0000_0000_0000_0000;
array[59715] <= 16'b0000_0000_0000_0000;
array[59716] <= 16'b0000_0000_0000_0000;
array[59717] <= 16'b0000_0000_0000_0000;
array[59718] <= 16'b0000_0000_0000_0000;
array[59719] <= 16'b0000_0000_0000_0000;
array[59720] <= 16'b0000_0000_0000_0000;
array[59721] <= 16'b0000_0000_0000_0000;
array[59722] <= 16'b0000_0000_0000_0000;
array[59723] <= 16'b0000_0000_0000_0000;
array[59724] <= 16'b0000_0000_0000_0000;
array[59725] <= 16'b0000_0000_0000_0000;
array[59726] <= 16'b0000_0000_0000_0000;
array[59727] <= 16'b0000_0000_0000_0000;
array[59728] <= 16'b0000_0000_0000_0000;
array[59729] <= 16'b0000_0000_0000_0000;
array[59730] <= 16'b0000_0000_0000_0000;
array[59731] <= 16'b0000_0000_0000_0000;
array[59732] <= 16'b0000_0000_0000_0000;
array[59733] <= 16'b0000_0000_0000_0000;
array[59734] <= 16'b0000_0000_0000_0000;
array[59735] <= 16'b0000_0000_0000_0000;
array[59736] <= 16'b0000_0000_0000_0000;
array[59737] <= 16'b0000_0000_0000_0000;
array[59738] <= 16'b0000_0000_0000_0000;
array[59739] <= 16'b0000_0000_0000_0000;
array[59740] <= 16'b0000_0000_0000_0000;
array[59741] <= 16'b0000_0000_0000_0000;
array[59742] <= 16'b0000_0000_0000_0000;
array[59743] <= 16'b0000_0000_0000_0000;
array[59744] <= 16'b0000_0000_0000_0000;
array[59745] <= 16'b0000_0000_0000_0000;
array[59746] <= 16'b0000_0000_0000_0000;
array[59747] <= 16'b0000_0000_0000_0000;
array[59748] <= 16'b0000_0000_0000_0000;
array[59749] <= 16'b0000_0000_0000_0000;
array[59750] <= 16'b0000_0000_0000_0000;
array[59751] <= 16'b0000_0000_0000_0000;
array[59752] <= 16'b0000_0000_0000_0000;
array[59753] <= 16'b0000_0000_0000_0000;
array[59754] <= 16'b0000_0000_0000_0000;
array[59755] <= 16'b0000_0000_0000_0000;
array[59756] <= 16'b0000_0000_0000_0000;
array[59757] <= 16'b0000_0000_0000_0000;
array[59758] <= 16'b0000_0000_0000_0000;
array[59759] <= 16'b0000_0000_0000_0000;
array[59760] <= 16'b0000_0000_0000_0000;
array[59761] <= 16'b0000_0000_0000_0000;
array[59762] <= 16'b0000_0000_0000_0000;
array[59763] <= 16'b0000_0000_0000_0000;
array[59764] <= 16'b0000_0000_0000_0000;
array[59765] <= 16'b0000_0000_0000_0000;
array[59766] <= 16'b0000_0000_0000_0000;
array[59767] <= 16'b0000_0000_0000_0000;
array[59768] <= 16'b0000_0000_0000_0000;
array[59769] <= 16'b0000_0000_0000_0000;
array[59770] <= 16'b0000_0000_0000_0000;
array[59771] <= 16'b0000_0000_0000_0000;
array[59772] <= 16'b0000_0000_0000_0000;
array[59773] <= 16'b0000_0000_0000_0000;
array[59774] <= 16'b0000_0000_0000_0000;
array[59775] <= 16'b0000_0000_0000_0000;
array[59776] <= 16'b0000_0000_0000_0000;
array[59777] <= 16'b0000_0000_0000_0000;
array[59778] <= 16'b0000_0000_0000_0000;
array[59779] <= 16'b0000_0000_0000_0000;
array[59780] <= 16'b0000_0000_0000_0000;
array[59781] <= 16'b0000_0000_0000_0000;
array[59782] <= 16'b0000_0000_0000_0000;
array[59783] <= 16'b0000_0000_0000_0000;
array[59784] <= 16'b0000_0000_0000_0000;
array[59785] <= 16'b0000_0000_0000_0000;
array[59786] <= 16'b0000_0000_0000_0000;
array[59787] <= 16'b0000_0000_0000_0000;
array[59788] <= 16'b0000_0000_0000_0000;
array[59789] <= 16'b0000_0000_0000_0000;
array[59790] <= 16'b0000_0000_0000_0000;
array[59791] <= 16'b0000_0000_0000_0000;
array[59792] <= 16'b0000_0000_0000_0000;
array[59793] <= 16'b0000_0000_0000_0000;
array[59794] <= 16'b0000_0000_0000_0000;
array[59795] <= 16'b0000_0000_0000_0000;
array[59796] <= 16'b0000_0000_0000_0000;
array[59797] <= 16'b0000_0000_0000_0000;
array[59798] <= 16'b0000_0000_0000_0000;
array[59799] <= 16'b0000_0000_0000_0000;
array[59800] <= 16'b0000_0000_0000_0000;
array[59801] <= 16'b0000_0000_0000_0000;
array[59802] <= 16'b0000_0000_0000_0000;
array[59803] <= 16'b0000_0000_0000_0000;
array[59804] <= 16'b0000_0000_0000_0000;
array[59805] <= 16'b0000_0000_0000_0000;
array[59806] <= 16'b0000_0000_0000_0000;
array[59807] <= 16'b0000_0000_0000_0000;
array[59808] <= 16'b0000_0000_0000_0000;
array[59809] <= 16'b0000_0000_0000_0000;
array[59810] <= 16'b0000_0000_0000_0000;
array[59811] <= 16'b0000_0000_0000_0000;
array[59812] <= 16'b0000_0000_0000_0000;
array[59813] <= 16'b0000_0000_0000_0000;
array[59814] <= 16'b0000_0000_0000_0000;
array[59815] <= 16'b0000_0000_0000_0000;
array[59816] <= 16'b0000_0000_0000_0000;
array[59817] <= 16'b0000_0000_0000_0000;
array[59818] <= 16'b0000_0000_0000_0000;
array[59819] <= 16'b0000_0000_0000_0000;
array[59820] <= 16'b0000_0000_0000_0000;
array[59821] <= 16'b0000_0000_0000_0000;
array[59822] <= 16'b0000_0000_0000_0000;
array[59823] <= 16'b0000_0000_0000_0000;
array[59824] <= 16'b0000_0000_0000_0000;
array[59825] <= 16'b0000_0000_0000_0000;
array[59826] <= 16'b0000_0000_0000_0000;
array[59827] <= 16'b0000_0000_0000_0000;
array[59828] <= 16'b0000_0000_0000_0000;
array[59829] <= 16'b0000_0000_0000_0000;
array[59830] <= 16'b0000_0000_0000_0000;
array[59831] <= 16'b0000_0000_0000_0000;
array[59832] <= 16'b0000_0000_0000_0000;
array[59833] <= 16'b0000_0000_0000_0000;
array[59834] <= 16'b0000_0000_0000_0000;
array[59835] <= 16'b0000_0000_0000_0000;
array[59836] <= 16'b0000_0000_0000_0000;
array[59837] <= 16'b0000_0000_0000_0000;
array[59838] <= 16'b0000_0000_0000_0000;
array[59839] <= 16'b0000_0000_0000_0000;
array[59840] <= 16'b0000_0000_0000_0000;
array[59841] <= 16'b0000_0000_0000_0000;
array[59842] <= 16'b0000_0000_0000_0000;
array[59843] <= 16'b0000_0000_0000_0000;
array[59844] <= 16'b0000_0000_0000_0000;
array[59845] <= 16'b0000_0000_0000_0000;
array[59846] <= 16'b0000_0000_0000_0000;
array[59847] <= 16'b0000_0000_0000_0000;
array[59848] <= 16'b0000_0000_0000_0000;
array[59849] <= 16'b0000_0000_0000_0000;
array[59850] <= 16'b0000_0000_0000_0000;
array[59851] <= 16'b0000_0000_0000_0000;
array[59852] <= 16'b0000_0000_0000_0000;
array[59853] <= 16'b0000_0000_0000_0000;
array[59854] <= 16'b0000_0000_0000_0000;
array[59855] <= 16'b0000_0000_0000_0000;
array[59856] <= 16'b0000_0000_0000_0000;
array[59857] <= 16'b0000_0000_0000_0000;
array[59858] <= 16'b0000_0000_0000_0000;
array[59859] <= 16'b0000_0000_0000_0000;
array[59860] <= 16'b0000_0000_0000_0000;
array[59861] <= 16'b0000_0000_0000_0000;
array[59862] <= 16'b0000_0000_0000_0000;
array[59863] <= 16'b0000_0000_0000_0000;
array[59864] <= 16'b0000_0000_0000_0000;
array[59865] <= 16'b0000_0000_0000_0000;
array[59866] <= 16'b0000_0000_0000_0000;
array[59867] <= 16'b0000_0000_0000_0000;
array[59868] <= 16'b0000_0000_0000_0000;
array[59869] <= 16'b0000_0000_0000_0000;
array[59870] <= 16'b0000_0000_0000_0000;
array[59871] <= 16'b0000_0000_0000_0000;
array[59872] <= 16'b0000_0000_0000_0000;
array[59873] <= 16'b0000_0000_0000_0000;
array[59874] <= 16'b0000_0000_0000_0000;
array[59875] <= 16'b0000_0000_0000_0000;
array[59876] <= 16'b0000_0000_0000_0000;
array[59877] <= 16'b0000_0000_0000_0000;
array[59878] <= 16'b0000_0000_0000_0000;
array[59879] <= 16'b0000_0000_0000_0000;
array[59880] <= 16'b0000_0000_0000_0000;
array[59881] <= 16'b0000_0000_0000_0000;
array[59882] <= 16'b0000_0000_0000_0000;
array[59883] <= 16'b0000_0000_0000_0000;
array[59884] <= 16'b0000_0000_0000_0000;
array[59885] <= 16'b0000_0000_0000_0000;
array[59886] <= 16'b0000_0000_0000_0000;
array[59887] <= 16'b0000_0000_0000_0000;
array[59888] <= 16'b0000_0000_0000_0000;
array[59889] <= 16'b0000_0000_0000_0000;
array[59890] <= 16'b0000_0000_0000_0000;
array[59891] <= 16'b0000_0000_0000_0000;
array[59892] <= 16'b0000_0000_0000_0000;
array[59893] <= 16'b0000_0000_0000_0000;
array[59894] <= 16'b0000_0000_0000_0000;
array[59895] <= 16'b0000_0000_0000_0000;
array[59896] <= 16'b0000_0000_0000_0000;
array[59897] <= 16'b0000_0000_0000_0000;
array[59898] <= 16'b0000_0000_0000_0000;
array[59899] <= 16'b0000_0000_0000_0000;
array[59900] <= 16'b0000_0000_0000_0000;
array[59901] <= 16'b0000_0000_0000_0000;
array[59902] <= 16'b0000_0000_0000_0000;
array[59903] <= 16'b0000_0000_0000_0000;
array[59904] <= 16'b0000_0000_0000_0000;
array[59905] <= 16'b0000_0000_0000_0000;
array[59906] <= 16'b0000_0000_0000_0000;
array[59907] <= 16'b0000_0000_0000_0000;
array[59908] <= 16'b0000_0000_0000_0000;
array[59909] <= 16'b0000_0000_0000_0000;
array[59910] <= 16'b0000_0000_0000_0000;
array[59911] <= 16'b0000_0000_0000_0000;
array[59912] <= 16'b0000_0000_0000_0000;
array[59913] <= 16'b0000_0000_0000_0000;
array[59914] <= 16'b0000_0000_0000_0000;
array[59915] <= 16'b0000_0000_0000_0000;
array[59916] <= 16'b0000_0000_0000_0000;
array[59917] <= 16'b0000_0000_0000_0000;
array[59918] <= 16'b0000_0000_0000_0000;
array[59919] <= 16'b0000_0000_0000_0000;
array[59920] <= 16'b0000_0000_0000_0000;
array[59921] <= 16'b0000_0000_0000_0000;
array[59922] <= 16'b0000_0000_0000_0000;
array[59923] <= 16'b0000_0000_0000_0000;
array[59924] <= 16'b0000_0000_0000_0000;
array[59925] <= 16'b0000_0000_0000_0000;
array[59926] <= 16'b0000_0000_0000_0000;
array[59927] <= 16'b0000_0000_0000_0000;
array[59928] <= 16'b0000_0000_0000_0000;
array[59929] <= 16'b0000_0000_0000_0000;
array[59930] <= 16'b0000_0000_0000_0000;
array[59931] <= 16'b0000_0000_0000_0000;
array[59932] <= 16'b0000_0000_0000_0000;
array[59933] <= 16'b0000_0000_0000_0000;
array[59934] <= 16'b0000_0000_0000_0000;
array[59935] <= 16'b0000_0000_0000_0000;
array[59936] <= 16'b0000_0000_0000_0000;
array[59937] <= 16'b0000_0000_0000_0000;
array[59938] <= 16'b0000_0000_0000_0000;
array[59939] <= 16'b0000_0000_0000_0000;
array[59940] <= 16'b0000_0000_0000_0000;
array[59941] <= 16'b0000_0000_0000_0000;
array[59942] <= 16'b0000_0000_0000_0000;
array[59943] <= 16'b0000_0000_0000_0000;
array[59944] <= 16'b0000_0000_0000_0000;
array[59945] <= 16'b0000_0000_0000_0000;
array[59946] <= 16'b0000_0000_0000_0000;
array[59947] <= 16'b0000_0000_0000_0000;
array[59948] <= 16'b0000_0000_0000_0000;
array[59949] <= 16'b0000_0000_0000_0000;
array[59950] <= 16'b0000_0000_0000_0000;
array[59951] <= 16'b0000_0000_0000_0000;
array[59952] <= 16'b0000_0000_0000_0000;
array[59953] <= 16'b0000_0000_0000_0000;
array[59954] <= 16'b0000_0000_0000_0000;
array[59955] <= 16'b0000_0000_0000_0000;
array[59956] <= 16'b0000_0000_0000_0000;
array[59957] <= 16'b0000_0000_0000_0000;
array[59958] <= 16'b0000_0000_0000_0000;
array[59959] <= 16'b0000_0000_0000_0000;
array[59960] <= 16'b0000_0000_0000_0000;
array[59961] <= 16'b0000_0000_0000_0000;
array[59962] <= 16'b0000_0000_0000_0000;
array[59963] <= 16'b0000_0000_0000_0000;
array[59964] <= 16'b0000_0000_0000_0000;
array[59965] <= 16'b0000_0000_0000_0000;
array[59966] <= 16'b0000_0000_0000_0000;
array[59967] <= 16'b0000_0000_0000_0000;
array[59968] <= 16'b0000_0000_0000_0000;
array[59969] <= 16'b0000_0000_0000_0000;
array[59970] <= 16'b0000_0000_0000_0000;
array[59971] <= 16'b0000_0000_0000_0000;
array[59972] <= 16'b0000_0000_0000_0000;
array[59973] <= 16'b0000_0000_0000_0000;
array[59974] <= 16'b0000_0000_0000_0000;
array[59975] <= 16'b0000_0000_0000_0000;
array[59976] <= 16'b0000_0000_0000_0000;
array[59977] <= 16'b0000_0000_0000_0000;
array[59978] <= 16'b0000_0000_0000_0000;
array[59979] <= 16'b0000_0000_0000_0000;
array[59980] <= 16'b0000_0000_0000_0000;
array[59981] <= 16'b0000_0000_0000_0000;
array[59982] <= 16'b0000_0000_0000_0000;
array[59983] <= 16'b0000_0000_0000_0000;
array[59984] <= 16'b0000_0000_0000_0000;
array[59985] <= 16'b0000_0000_0000_0000;
array[59986] <= 16'b0000_0000_0000_0000;
array[59987] <= 16'b0000_0000_0000_0000;
array[59988] <= 16'b0000_0000_0000_0000;
array[59989] <= 16'b0000_0000_0000_0000;
array[59990] <= 16'b0000_0000_0000_0000;
array[59991] <= 16'b0000_0000_0000_0000;
array[59992] <= 16'b0000_0000_0000_0000;
array[59993] <= 16'b0000_0000_0000_0000;
array[59994] <= 16'b0000_0000_0000_0000;
array[59995] <= 16'b0000_0000_0000_0000;
array[59996] <= 16'b0000_0000_0000_0000;
array[59997] <= 16'b0000_0000_0000_0000;
array[59998] <= 16'b0000_0000_0000_0000;
array[59999] <= 16'b0000_0000_0000_0000;
array[60000] <= 16'b0000_0000_0000_0000;
array[60001] <= 16'b0000_0000_0000_0000;
array[60002] <= 16'b0000_0000_0000_0000;
array[60003] <= 16'b0000_0000_0000_0000;
array[60004] <= 16'b0000_0000_0000_0000;
array[60005] <= 16'b0000_0000_0000_0000;
array[60006] <= 16'b0000_0000_0000_0000;
array[60007] <= 16'b0000_0000_0000_0000;
array[60008] <= 16'b0000_0000_0000_0000;
array[60009] <= 16'b0000_0000_0000_0000;
array[60010] <= 16'b0000_0000_0000_0000;
array[60011] <= 16'b0000_0000_0000_0000;
array[60012] <= 16'b0000_0000_0000_0000;
array[60013] <= 16'b0000_0000_0000_0000;
array[60014] <= 16'b0000_0000_0000_0000;
array[60015] <= 16'b0000_0000_0000_0000;
array[60016] <= 16'b0000_0000_0000_0000;
array[60017] <= 16'b0000_0000_0000_0000;
array[60018] <= 16'b0000_0000_0000_0000;
array[60019] <= 16'b0000_0000_0000_0000;
array[60020] <= 16'b0000_0000_0000_0000;
array[60021] <= 16'b0000_0000_0000_0000;
array[60022] <= 16'b0000_0000_0000_0000;
array[60023] <= 16'b0000_0000_0000_0000;
array[60024] <= 16'b0000_0000_0000_0000;
array[60025] <= 16'b0000_0000_0000_0000;
array[60026] <= 16'b0000_0000_0000_0000;
array[60027] <= 16'b0000_0000_0000_0000;
array[60028] <= 16'b0000_0000_0000_0000;
array[60029] <= 16'b0000_0000_0000_0000;
array[60030] <= 16'b0000_0000_0000_0000;
array[60031] <= 16'b0000_0000_0000_0000;
array[60032] <= 16'b0000_0000_0000_0000;
array[60033] <= 16'b0000_0000_0000_0000;
array[60034] <= 16'b0000_0000_0000_0000;
array[60035] <= 16'b0000_0000_0000_0000;
array[60036] <= 16'b0000_0000_0000_0000;
array[60037] <= 16'b0000_0000_0000_0000;
array[60038] <= 16'b0000_0000_0000_0000;
array[60039] <= 16'b0000_0000_0000_0000;
array[60040] <= 16'b0000_0000_0000_0000;
array[60041] <= 16'b0000_0000_0000_0000;
array[60042] <= 16'b0000_0000_0000_0000;
array[60043] <= 16'b0000_0000_0000_0000;
array[60044] <= 16'b0000_0000_0000_0000;
array[60045] <= 16'b0000_0000_0000_0000;
array[60046] <= 16'b0000_0000_0000_0000;
array[60047] <= 16'b0000_0000_0000_0000;
array[60048] <= 16'b0000_0000_0000_0000;
array[60049] <= 16'b0000_0000_0000_0000;
array[60050] <= 16'b0000_0000_0000_0000;
array[60051] <= 16'b0000_0000_0000_0000;
array[60052] <= 16'b0000_0000_0000_0000;
array[60053] <= 16'b0000_0000_0000_0000;
array[60054] <= 16'b0000_0000_0000_0000;
array[60055] <= 16'b0000_0000_0000_0000;
array[60056] <= 16'b0000_0000_0000_0000;
array[60057] <= 16'b0000_0000_0000_0000;
array[60058] <= 16'b0000_0000_0000_0000;
array[60059] <= 16'b0000_0000_0000_0000;
array[60060] <= 16'b0000_0000_0000_0000;
array[60061] <= 16'b0000_0000_0000_0000;
array[60062] <= 16'b0000_0000_0000_0000;
array[60063] <= 16'b0000_0000_0000_0000;
array[60064] <= 16'b0000_0000_0000_0000;
array[60065] <= 16'b0000_0000_0000_0000;
array[60066] <= 16'b0000_0000_0000_0000;
array[60067] <= 16'b0000_0000_0000_0000;
array[60068] <= 16'b0000_0000_0000_0000;
array[60069] <= 16'b0000_0000_0000_0000;
array[60070] <= 16'b0000_0000_0000_0000;
array[60071] <= 16'b0000_0000_0000_0000;
array[60072] <= 16'b0000_0000_0000_0000;
array[60073] <= 16'b0000_0000_0000_0000;
array[60074] <= 16'b0000_0000_0000_0000;
array[60075] <= 16'b0000_0000_0000_0000;
array[60076] <= 16'b0000_0000_0000_0000;
array[60077] <= 16'b0000_0000_0000_0000;
array[60078] <= 16'b0000_0000_0000_0000;
array[60079] <= 16'b0000_0000_0000_0000;
array[60080] <= 16'b0000_0000_0000_0000;
array[60081] <= 16'b0000_0000_0000_0000;
array[60082] <= 16'b0000_0000_0000_0000;
array[60083] <= 16'b0000_0000_0000_0000;
array[60084] <= 16'b0000_0000_0000_0000;
array[60085] <= 16'b0000_0000_0000_0000;
array[60086] <= 16'b0000_0000_0000_0000;
array[60087] <= 16'b0000_0000_0000_0000;
array[60088] <= 16'b0000_0000_0000_0000;
array[60089] <= 16'b0000_0000_0000_0000;
array[60090] <= 16'b0000_0000_0000_0000;
array[60091] <= 16'b0000_0000_0000_0000;
array[60092] <= 16'b0000_0000_0000_0000;
array[60093] <= 16'b0000_0000_0000_0000;
array[60094] <= 16'b0000_0000_0000_0000;
array[60095] <= 16'b0000_0000_0000_0000;
array[60096] <= 16'b0000_0000_0000_0000;
array[60097] <= 16'b0000_0000_0000_0000;
array[60098] <= 16'b0000_0000_0000_0000;
array[60099] <= 16'b0000_0000_0000_0000;
array[60100] <= 16'b0000_0000_0000_0000;
array[60101] <= 16'b0000_0000_0000_0000;
array[60102] <= 16'b0000_0000_0000_0000;
array[60103] <= 16'b0000_0000_0000_0000;
array[60104] <= 16'b0000_0000_0000_0000;
array[60105] <= 16'b0000_0000_0000_0000;
array[60106] <= 16'b0000_0000_0000_0000;
array[60107] <= 16'b0000_0000_0000_0000;
array[60108] <= 16'b0000_0000_0000_0000;
array[60109] <= 16'b0000_0000_0000_0000;
array[60110] <= 16'b0000_0000_0000_0000;
array[60111] <= 16'b0000_0000_0000_0000;
array[60112] <= 16'b0000_0000_0000_0000;
array[60113] <= 16'b0000_0000_0000_0000;
array[60114] <= 16'b0000_0000_0000_0000;
array[60115] <= 16'b0000_0000_0000_0000;
array[60116] <= 16'b0000_0000_0000_0000;
array[60117] <= 16'b0000_0000_0000_0000;
array[60118] <= 16'b0000_0000_0000_0000;
array[60119] <= 16'b0000_0000_0000_0000;
array[60120] <= 16'b0000_0000_0000_0000;
array[60121] <= 16'b0000_0000_0000_0000;
array[60122] <= 16'b0000_0000_0000_0000;
array[60123] <= 16'b0000_0000_0000_0000;
array[60124] <= 16'b0000_0000_0000_0000;
array[60125] <= 16'b0000_0000_0000_0000;
array[60126] <= 16'b0000_0000_0000_0000;
array[60127] <= 16'b0000_0000_0000_0000;
array[60128] <= 16'b0000_0000_0000_0000;
array[60129] <= 16'b0000_0000_0000_0000;
array[60130] <= 16'b0000_0000_0000_0000;
array[60131] <= 16'b0000_0000_0000_0000;
array[60132] <= 16'b0000_0000_0000_0000;
array[60133] <= 16'b0000_0000_0000_0000;
array[60134] <= 16'b0000_0000_0000_0000;
array[60135] <= 16'b0000_0000_0000_0000;
array[60136] <= 16'b0000_0000_0000_0000;
array[60137] <= 16'b0000_0000_0000_0000;
array[60138] <= 16'b0000_0000_0000_0000;
array[60139] <= 16'b0000_0000_0000_0000;
array[60140] <= 16'b0000_0000_0000_0000;
array[60141] <= 16'b0000_0000_0000_0000;
array[60142] <= 16'b0000_0000_0000_0000;
array[60143] <= 16'b0000_0000_0000_0000;
array[60144] <= 16'b0000_0000_0000_0000;
array[60145] <= 16'b0000_0000_0000_0000;
array[60146] <= 16'b0000_0000_0000_0000;
array[60147] <= 16'b0000_0000_0000_0000;
array[60148] <= 16'b0000_0000_0000_0000;
array[60149] <= 16'b0000_0000_0000_0000;
array[60150] <= 16'b0000_0000_0000_0000;
array[60151] <= 16'b0000_0000_0000_0000;
array[60152] <= 16'b0000_0000_0000_0000;
array[60153] <= 16'b0000_0000_0000_0000;
array[60154] <= 16'b0000_0000_0000_0000;
array[60155] <= 16'b0000_0000_0000_0000;
array[60156] <= 16'b0000_0000_0000_0000;
array[60157] <= 16'b0000_0000_0000_0000;
array[60158] <= 16'b0000_0000_0000_0000;
array[60159] <= 16'b0000_0000_0000_0000;
array[60160] <= 16'b0000_0000_0000_0000;
array[60161] <= 16'b0000_0000_0000_0000;
array[60162] <= 16'b0000_0000_0000_0000;
array[60163] <= 16'b0000_0000_0000_0000;
array[60164] <= 16'b0000_0000_0000_0000;
array[60165] <= 16'b0000_0000_0000_0000;
array[60166] <= 16'b0000_0000_0000_0000;
array[60167] <= 16'b0000_0000_0000_0000;
array[60168] <= 16'b0000_0000_0000_0000;
array[60169] <= 16'b0000_0000_0000_0000;
array[60170] <= 16'b0000_0000_0000_0000;
array[60171] <= 16'b0000_0000_0000_0000;
array[60172] <= 16'b0000_0000_0000_0000;
array[60173] <= 16'b0000_0000_0000_0000;
array[60174] <= 16'b0000_0000_0000_0000;
array[60175] <= 16'b0000_0000_0000_0000;
array[60176] <= 16'b0000_0000_0000_0000;
array[60177] <= 16'b0000_0000_0000_0000;
array[60178] <= 16'b0000_0000_0000_0000;
array[60179] <= 16'b0000_0000_0000_0000;
array[60180] <= 16'b0000_0000_0000_0000;
array[60181] <= 16'b0000_0000_0000_0000;
array[60182] <= 16'b0000_0000_0000_0000;
array[60183] <= 16'b0000_0000_0000_0000;
array[60184] <= 16'b0000_0000_0000_0000;
array[60185] <= 16'b0000_0000_0000_0000;
array[60186] <= 16'b0000_0000_0000_0000;
array[60187] <= 16'b0000_0000_0000_0000;
array[60188] <= 16'b0000_0000_0000_0000;
array[60189] <= 16'b0000_0000_0000_0000;
array[60190] <= 16'b0000_0000_0000_0000;
array[60191] <= 16'b0000_0000_0000_0000;
array[60192] <= 16'b0000_0000_0000_0000;
array[60193] <= 16'b0000_0000_0000_0000;
array[60194] <= 16'b0000_0000_0000_0000;
array[60195] <= 16'b0000_0000_0000_0000;
array[60196] <= 16'b0000_0000_0000_0000;
array[60197] <= 16'b0000_0000_0000_0000;
array[60198] <= 16'b0000_0000_0000_0000;
array[60199] <= 16'b0000_0000_0000_0000;
array[60200] <= 16'b0000_0000_0000_0000;
array[60201] <= 16'b0000_0000_0000_0000;
array[60202] <= 16'b0000_0000_0000_0000;
array[60203] <= 16'b0000_0000_0000_0000;
array[60204] <= 16'b0000_0000_0000_0000;
array[60205] <= 16'b0000_0000_0000_0000;
array[60206] <= 16'b0000_0000_0000_0000;
array[60207] <= 16'b0000_0000_0000_0000;
array[60208] <= 16'b0000_0000_0000_0000;
array[60209] <= 16'b0000_0000_0000_0000;
array[60210] <= 16'b0000_0000_0000_0000;
array[60211] <= 16'b0000_0000_0000_0000;
array[60212] <= 16'b0000_0000_0000_0000;
array[60213] <= 16'b0000_0000_0000_0000;
array[60214] <= 16'b0000_0000_0000_0000;
array[60215] <= 16'b0000_0000_0000_0000;
array[60216] <= 16'b0000_0000_0000_0000;
array[60217] <= 16'b0000_0000_0000_0000;
array[60218] <= 16'b0000_0000_0000_0000;
array[60219] <= 16'b0000_0000_0000_0000;
array[60220] <= 16'b0000_0000_0000_0000;
array[60221] <= 16'b0000_0000_0000_0000;
array[60222] <= 16'b0000_0000_0000_0000;
array[60223] <= 16'b0000_0000_0000_0000;
array[60224] <= 16'b0000_0000_0000_0000;
array[60225] <= 16'b0000_0000_0000_0000;
array[60226] <= 16'b0000_0000_0000_0000;
array[60227] <= 16'b0000_0000_0000_0000;
array[60228] <= 16'b0000_0000_0000_0000;
array[60229] <= 16'b0000_0000_0000_0000;
array[60230] <= 16'b0000_0000_0000_0000;
array[60231] <= 16'b0000_0000_0000_0000;
array[60232] <= 16'b0000_0000_0000_0000;
array[60233] <= 16'b0000_0000_0000_0000;
array[60234] <= 16'b0000_0000_0000_0000;
array[60235] <= 16'b0000_0000_0000_0000;
array[60236] <= 16'b0000_0000_0000_0000;
array[60237] <= 16'b0000_0000_0000_0000;
array[60238] <= 16'b0000_0000_0000_0000;
array[60239] <= 16'b0000_0000_0000_0000;
array[60240] <= 16'b0000_0000_0000_0000;
array[60241] <= 16'b0000_0000_0000_0000;
array[60242] <= 16'b0000_0000_0000_0000;
array[60243] <= 16'b0000_0000_0000_0000;
array[60244] <= 16'b0000_0000_0000_0000;
array[60245] <= 16'b0000_0000_0000_0000;
array[60246] <= 16'b0000_0000_0000_0000;
array[60247] <= 16'b0000_0000_0000_0000;
array[60248] <= 16'b0000_0000_0000_0000;
array[60249] <= 16'b0000_0000_0000_0000;
array[60250] <= 16'b0000_0000_0000_0000;
array[60251] <= 16'b0000_0000_0000_0000;
array[60252] <= 16'b0000_0000_0000_0000;
array[60253] <= 16'b0000_0000_0000_0000;
array[60254] <= 16'b0000_0000_0000_0000;
array[60255] <= 16'b0000_0000_0000_0000;
array[60256] <= 16'b0000_0000_0000_0000;
array[60257] <= 16'b0000_0000_0000_0000;
array[60258] <= 16'b0000_0000_0000_0000;
array[60259] <= 16'b0000_0000_0000_0000;
array[60260] <= 16'b0000_0000_0000_0000;
array[60261] <= 16'b0000_0000_0000_0000;
array[60262] <= 16'b0000_0000_0000_0000;
array[60263] <= 16'b0000_0000_0000_0000;
array[60264] <= 16'b0000_0000_0000_0000;
array[60265] <= 16'b0000_0000_0000_0000;
array[60266] <= 16'b0000_0000_0000_0000;
array[60267] <= 16'b0000_0000_0000_0000;
array[60268] <= 16'b0000_0000_0000_0000;
array[60269] <= 16'b0000_0000_0000_0000;
array[60270] <= 16'b0000_0000_0000_0000;
array[60271] <= 16'b0000_0000_0000_0000;
array[60272] <= 16'b0000_0000_0000_0000;
array[60273] <= 16'b0000_0000_0000_0000;
array[60274] <= 16'b0000_0000_0000_0000;
array[60275] <= 16'b0000_0000_0000_0000;
array[60276] <= 16'b0000_0000_0000_0000;
array[60277] <= 16'b0000_0000_0000_0000;
array[60278] <= 16'b0000_0000_0000_0000;
array[60279] <= 16'b0000_0000_0000_0000;
array[60280] <= 16'b0000_0000_0000_0000;
array[60281] <= 16'b0000_0000_0000_0000;
array[60282] <= 16'b0000_0000_0000_0000;
array[60283] <= 16'b0000_0000_0000_0000;
array[60284] <= 16'b0000_0000_0000_0000;
array[60285] <= 16'b0000_0000_0000_0000;
array[60286] <= 16'b0000_0000_0000_0000;
array[60287] <= 16'b0000_0000_0000_0000;
array[60288] <= 16'b0000_0000_0000_0000;
array[60289] <= 16'b0000_0000_0000_0000;
array[60290] <= 16'b0000_0000_0000_0000;
array[60291] <= 16'b0000_0000_0000_0000;
array[60292] <= 16'b0000_0000_0000_0000;
array[60293] <= 16'b0000_0000_0000_0000;
array[60294] <= 16'b0000_0000_0000_0000;
array[60295] <= 16'b0000_0000_0000_0000;
array[60296] <= 16'b0000_0000_0000_0000;
array[60297] <= 16'b0000_0000_0000_0000;
array[60298] <= 16'b0000_0000_0000_0000;
array[60299] <= 16'b0000_0000_0000_0000;
array[60300] <= 16'b0000_0000_0000_0000;
array[60301] <= 16'b0000_0000_0000_0000;
array[60302] <= 16'b0000_0000_0000_0000;
array[60303] <= 16'b0000_0000_0000_0000;
array[60304] <= 16'b0000_0000_0000_0000;
array[60305] <= 16'b0000_0000_0000_0000;
array[60306] <= 16'b0000_0000_0000_0000;
array[60307] <= 16'b0000_0000_0000_0000;
array[60308] <= 16'b0000_0000_0000_0000;
array[60309] <= 16'b0000_0000_0000_0000;
array[60310] <= 16'b0000_0000_0000_0000;
array[60311] <= 16'b0000_0000_0000_0000;
array[60312] <= 16'b0000_0000_0000_0000;
array[60313] <= 16'b0000_0000_0000_0000;
array[60314] <= 16'b0000_0000_0000_0000;
array[60315] <= 16'b0000_0000_0000_0000;
array[60316] <= 16'b0000_0000_0000_0000;
array[60317] <= 16'b0000_0000_0000_0000;
array[60318] <= 16'b0000_0000_0000_0000;
array[60319] <= 16'b0000_0000_0000_0000;
array[60320] <= 16'b0000_0000_0000_0000;
array[60321] <= 16'b0000_0000_0000_0000;
array[60322] <= 16'b0000_0000_0000_0000;
array[60323] <= 16'b0000_0000_0000_0000;
array[60324] <= 16'b0000_0000_0000_0000;
array[60325] <= 16'b0000_0000_0000_0000;
array[60326] <= 16'b0000_0000_0000_0000;
array[60327] <= 16'b0000_0000_0000_0000;
array[60328] <= 16'b0000_0000_0000_0000;
array[60329] <= 16'b0000_0000_0000_0000;
array[60330] <= 16'b0000_0000_0000_0000;
array[60331] <= 16'b0000_0000_0000_0000;
array[60332] <= 16'b0000_0000_0000_0000;
array[60333] <= 16'b0000_0000_0000_0000;
array[60334] <= 16'b0000_0000_0000_0000;
array[60335] <= 16'b0000_0000_0000_0000;
array[60336] <= 16'b0000_0000_0000_0000;
array[60337] <= 16'b0000_0000_0000_0000;
array[60338] <= 16'b0000_0000_0000_0000;
array[60339] <= 16'b0000_0000_0000_0000;
array[60340] <= 16'b0000_0000_0000_0000;
array[60341] <= 16'b0000_0000_0000_0000;
array[60342] <= 16'b0000_0000_0000_0000;
array[60343] <= 16'b0000_0000_0000_0000;
array[60344] <= 16'b0000_0000_0000_0000;
array[60345] <= 16'b0000_0000_0000_0000;
array[60346] <= 16'b0000_0000_0000_0000;
array[60347] <= 16'b0000_0000_0000_0000;
array[60348] <= 16'b0000_0000_0000_0000;
array[60349] <= 16'b0000_0000_0000_0000;
array[60350] <= 16'b0000_0000_0000_0000;
array[60351] <= 16'b0000_0000_0000_0000;
array[60352] <= 16'b0000_0000_0000_0000;
array[60353] <= 16'b0000_0000_0000_0000;
array[60354] <= 16'b0000_0000_0000_0000;
array[60355] <= 16'b0000_0000_0000_0000;
array[60356] <= 16'b0000_0000_0000_0000;
array[60357] <= 16'b0000_0000_0000_0000;
array[60358] <= 16'b0000_0000_0000_0000;
array[60359] <= 16'b0000_0000_0000_0000;
array[60360] <= 16'b0000_0000_0000_0000;
array[60361] <= 16'b0000_0000_0000_0000;
array[60362] <= 16'b0000_0000_0000_0000;
array[60363] <= 16'b0000_0000_0000_0000;
array[60364] <= 16'b0000_0000_0000_0000;
array[60365] <= 16'b0000_0000_0000_0000;
array[60366] <= 16'b0000_0000_0000_0000;
array[60367] <= 16'b0000_0000_0000_0000;
array[60368] <= 16'b0000_0000_0000_0000;
array[60369] <= 16'b0000_0000_0000_0000;
array[60370] <= 16'b0000_0000_0000_0000;
array[60371] <= 16'b0000_0000_0000_0000;
array[60372] <= 16'b0000_0000_0000_0000;
array[60373] <= 16'b0000_0000_0000_0000;
array[60374] <= 16'b0000_0000_0000_0000;
array[60375] <= 16'b0000_0000_0000_0000;
array[60376] <= 16'b0000_0000_0000_0000;
array[60377] <= 16'b0000_0000_0000_0000;
array[60378] <= 16'b0000_0000_0000_0000;
array[60379] <= 16'b0000_0000_0000_0000;
array[60380] <= 16'b0000_0000_0000_0000;
array[60381] <= 16'b0000_0000_0000_0000;
array[60382] <= 16'b0000_0000_0000_0000;
array[60383] <= 16'b0000_0000_0000_0000;
array[60384] <= 16'b0000_0000_0000_0000;
array[60385] <= 16'b0000_0000_0000_0000;
array[60386] <= 16'b0000_0000_0000_0000;
array[60387] <= 16'b0000_0000_0000_0000;
array[60388] <= 16'b0000_0000_0000_0000;
array[60389] <= 16'b0000_0000_0000_0000;
array[60390] <= 16'b0000_0000_0000_0000;
array[60391] <= 16'b0000_0000_0000_0000;
array[60392] <= 16'b0000_0000_0000_0000;
array[60393] <= 16'b0000_0000_0000_0000;
array[60394] <= 16'b0000_0000_0000_0000;
array[60395] <= 16'b0000_0000_0000_0000;
array[60396] <= 16'b0000_0000_0000_0000;
array[60397] <= 16'b0000_0000_0000_0000;
array[60398] <= 16'b0000_0000_0000_0000;
array[60399] <= 16'b0000_0000_0000_0000;
array[60400] <= 16'b0000_0000_0000_0000;
array[60401] <= 16'b0000_0000_0000_0000;
array[60402] <= 16'b0000_0000_0000_0000;
array[60403] <= 16'b0000_0000_0000_0000;
array[60404] <= 16'b0000_0000_0000_0000;
array[60405] <= 16'b0000_0000_0000_0000;
array[60406] <= 16'b0000_0000_0000_0000;
array[60407] <= 16'b0000_0000_0000_0000;
array[60408] <= 16'b0000_0000_0000_0000;
array[60409] <= 16'b0000_0000_0000_0000;
array[60410] <= 16'b0000_0000_0000_0000;
array[60411] <= 16'b0000_0000_0000_0000;
array[60412] <= 16'b0000_0000_0000_0000;
array[60413] <= 16'b0000_0000_0000_0000;
array[60414] <= 16'b0000_0000_0000_0000;
array[60415] <= 16'b0000_0000_0000_0000;
array[60416] <= 16'b0000_0000_0000_0000;
array[60417] <= 16'b0000_0000_0000_0000;
array[60418] <= 16'b0000_0000_0000_0000;
array[60419] <= 16'b0000_0000_0000_0000;
array[60420] <= 16'b0000_0000_0000_0000;
array[60421] <= 16'b0000_0000_0000_0000;
array[60422] <= 16'b0000_0000_0000_0000;
array[60423] <= 16'b0000_0000_0000_0000;
array[60424] <= 16'b0000_0000_0000_0000;
array[60425] <= 16'b0000_0000_0000_0000;
array[60426] <= 16'b0000_0000_0000_0000;
array[60427] <= 16'b0000_0000_0000_0000;
array[60428] <= 16'b0000_0000_0000_0000;
array[60429] <= 16'b0000_0000_0000_0000;
array[60430] <= 16'b0000_0000_0000_0000;
array[60431] <= 16'b0000_0000_0000_0000;
array[60432] <= 16'b0000_0000_0000_0000;
array[60433] <= 16'b0000_0000_0000_0000;
array[60434] <= 16'b0000_0000_0000_0000;
array[60435] <= 16'b0000_0000_0000_0000;
array[60436] <= 16'b0000_0000_0000_0000;
array[60437] <= 16'b0000_0000_0000_0000;
array[60438] <= 16'b0000_0000_0000_0000;
array[60439] <= 16'b0000_0000_0000_0000;
array[60440] <= 16'b0000_0000_0000_0000;
array[60441] <= 16'b0000_0000_0000_0000;
array[60442] <= 16'b0000_0000_0000_0000;
array[60443] <= 16'b0000_0000_0000_0000;
array[60444] <= 16'b0000_0000_0000_0000;
array[60445] <= 16'b0000_0000_0000_0000;
array[60446] <= 16'b0000_0000_0000_0000;
array[60447] <= 16'b0000_0000_0000_0000;
array[60448] <= 16'b0000_0000_0000_0000;
array[60449] <= 16'b0000_0000_0000_0000;
array[60450] <= 16'b0000_0000_0000_0000;
array[60451] <= 16'b0000_0000_0000_0000;
array[60452] <= 16'b0000_0000_0000_0000;
array[60453] <= 16'b0000_0000_0000_0000;
array[60454] <= 16'b0000_0000_0000_0000;
array[60455] <= 16'b0000_0000_0000_0000;
array[60456] <= 16'b0000_0000_0000_0000;
array[60457] <= 16'b0000_0000_0000_0000;
array[60458] <= 16'b0000_0000_0000_0000;
array[60459] <= 16'b0000_0000_0000_0000;
array[60460] <= 16'b0000_0000_0000_0000;
array[60461] <= 16'b0000_0000_0000_0000;
array[60462] <= 16'b0000_0000_0000_0000;
array[60463] <= 16'b0000_0000_0000_0000;
array[60464] <= 16'b0000_0000_0000_0000;
array[60465] <= 16'b0000_0000_0000_0000;
array[60466] <= 16'b0000_0000_0000_0000;
array[60467] <= 16'b0000_0000_0000_0000;
array[60468] <= 16'b0000_0000_0000_0000;
array[60469] <= 16'b0000_0000_0000_0000;
array[60470] <= 16'b0000_0000_0000_0000;
array[60471] <= 16'b0000_0000_0000_0000;
array[60472] <= 16'b0000_0000_0000_0000;
array[60473] <= 16'b0000_0000_0000_0000;
array[60474] <= 16'b0000_0000_0000_0000;
array[60475] <= 16'b0000_0000_0000_0000;
array[60476] <= 16'b0000_0000_0000_0000;
array[60477] <= 16'b0000_0000_0000_0000;
array[60478] <= 16'b0000_0000_0000_0000;
array[60479] <= 16'b0000_0000_0000_0000;
array[60480] <= 16'b0000_0000_0000_0000;
array[60481] <= 16'b0000_0000_0000_0000;
array[60482] <= 16'b0000_0000_0000_0000;
array[60483] <= 16'b0000_0000_0000_0000;
array[60484] <= 16'b0000_0000_0000_0000;
array[60485] <= 16'b0000_0000_0000_0000;
array[60486] <= 16'b0000_0000_0000_0000;
array[60487] <= 16'b0000_0000_0000_0000;
array[60488] <= 16'b0000_0000_0000_0000;
array[60489] <= 16'b0000_0000_0000_0000;
array[60490] <= 16'b0000_0000_0000_0000;
array[60491] <= 16'b0000_0000_0000_0000;
array[60492] <= 16'b0000_0000_0000_0000;
array[60493] <= 16'b0000_0000_0000_0000;
array[60494] <= 16'b0000_0000_0000_0000;
array[60495] <= 16'b0000_0000_0000_0000;
array[60496] <= 16'b0000_0000_0000_0000;
array[60497] <= 16'b0000_0000_0000_0000;
array[60498] <= 16'b0000_0000_0000_0000;
array[60499] <= 16'b0000_0000_0000_0000;
array[60500] <= 16'b0000_0000_0000_0000;
array[60501] <= 16'b0000_0000_0000_0000;
array[60502] <= 16'b0000_0000_0000_0000;
array[60503] <= 16'b0000_0000_0000_0000;
array[60504] <= 16'b0000_0000_0000_0000;
array[60505] <= 16'b0000_0000_0000_0000;
array[60506] <= 16'b0000_0000_0000_0000;
array[60507] <= 16'b0000_0000_0000_0000;
array[60508] <= 16'b0000_0000_0000_0000;
array[60509] <= 16'b0000_0000_0000_0000;
array[60510] <= 16'b0000_0000_0000_0000;
array[60511] <= 16'b0000_0000_0000_0000;
array[60512] <= 16'b0000_0000_0000_0000;
array[60513] <= 16'b0000_0000_0000_0000;
array[60514] <= 16'b0000_0000_0000_0000;
array[60515] <= 16'b0000_0000_0000_0000;
array[60516] <= 16'b0000_0000_0000_0000;
array[60517] <= 16'b0000_0000_0000_0000;
array[60518] <= 16'b0000_0000_0000_0000;
array[60519] <= 16'b0000_0000_0000_0000;
array[60520] <= 16'b0000_0000_0000_0000;
array[60521] <= 16'b0000_0000_0000_0000;
array[60522] <= 16'b0000_0000_0000_0000;
array[60523] <= 16'b0000_0000_0000_0000;
array[60524] <= 16'b0000_0000_0000_0000;
array[60525] <= 16'b0000_0000_0000_0000;
array[60526] <= 16'b0000_0000_0000_0000;
array[60527] <= 16'b0000_0000_0000_0000;
array[60528] <= 16'b0000_0000_0000_0000;
array[60529] <= 16'b0000_0000_0000_0000;
array[60530] <= 16'b0000_0000_0000_0000;
array[60531] <= 16'b0000_0000_0000_0000;
array[60532] <= 16'b0000_0000_0000_0000;
array[60533] <= 16'b0000_0000_0000_0000;
array[60534] <= 16'b0000_0000_0000_0000;
array[60535] <= 16'b0000_0000_0000_0000;
array[60536] <= 16'b0000_0000_0000_0000;
array[60537] <= 16'b0000_0000_0000_0000;
array[60538] <= 16'b0000_0000_0000_0000;
array[60539] <= 16'b0000_0000_0000_0000;
array[60540] <= 16'b0000_0000_0000_0000;
array[60541] <= 16'b0000_0000_0000_0000;
array[60542] <= 16'b0000_0000_0000_0000;
array[60543] <= 16'b0000_0000_0000_0000;
array[60544] <= 16'b0000_0000_0000_0000;
array[60545] <= 16'b0000_0000_0000_0000;
array[60546] <= 16'b0000_0000_0000_0000;
array[60547] <= 16'b0000_0000_0000_0000;
array[60548] <= 16'b0000_0000_0000_0000;
array[60549] <= 16'b0000_0000_0000_0000;
array[60550] <= 16'b0000_0000_0000_0000;
array[60551] <= 16'b0000_0000_0000_0000;
array[60552] <= 16'b0000_0000_0000_0000;
array[60553] <= 16'b0000_0000_0000_0000;
array[60554] <= 16'b0000_0000_0000_0000;
array[60555] <= 16'b0000_0000_0000_0000;
array[60556] <= 16'b0000_0000_0000_0000;
array[60557] <= 16'b0000_0000_0000_0000;
array[60558] <= 16'b0000_0000_0000_0000;
array[60559] <= 16'b0000_0000_0000_0000;
array[60560] <= 16'b0000_0000_0000_0000;
array[60561] <= 16'b0000_0000_0000_0000;
array[60562] <= 16'b0000_0000_0000_0000;
array[60563] <= 16'b0000_0000_0000_0000;
array[60564] <= 16'b0000_0000_0000_0000;
array[60565] <= 16'b0000_0000_0000_0000;
array[60566] <= 16'b0000_0000_0000_0000;
array[60567] <= 16'b0000_0000_0000_0000;
array[60568] <= 16'b0000_0000_0000_0000;
array[60569] <= 16'b0000_0000_0000_0000;
array[60570] <= 16'b0000_0000_0000_0000;
array[60571] <= 16'b0000_0000_0000_0000;
array[60572] <= 16'b0000_0000_0000_0000;
array[60573] <= 16'b0000_0000_0000_0000;
array[60574] <= 16'b0000_0000_0000_0000;
array[60575] <= 16'b0000_0000_0000_0000;
array[60576] <= 16'b0000_0000_0000_0000;
array[60577] <= 16'b0000_0000_0000_0000;
array[60578] <= 16'b0000_0000_0000_0000;
array[60579] <= 16'b0000_0000_0000_0000;
array[60580] <= 16'b0000_0000_0000_0000;
array[60581] <= 16'b0000_0000_0000_0000;
array[60582] <= 16'b0000_0000_0000_0000;
array[60583] <= 16'b0000_0000_0000_0000;
array[60584] <= 16'b0000_0000_0000_0000;
array[60585] <= 16'b0000_0000_0000_0000;
array[60586] <= 16'b0000_0000_0000_0000;
array[60587] <= 16'b0000_0000_0000_0000;
array[60588] <= 16'b0000_0000_0000_0000;
array[60589] <= 16'b0000_0000_0000_0000;
array[60590] <= 16'b0000_0000_0000_0000;
array[60591] <= 16'b0000_0000_0000_0000;
array[60592] <= 16'b0000_0000_0000_0000;
array[60593] <= 16'b0000_0000_0000_0000;
array[60594] <= 16'b0000_0000_0000_0000;
array[60595] <= 16'b0000_0000_0000_0000;
array[60596] <= 16'b0000_0000_0000_0000;
array[60597] <= 16'b0000_0000_0000_0000;
array[60598] <= 16'b0000_0000_0000_0000;
array[60599] <= 16'b0000_0000_0000_0000;
array[60600] <= 16'b0000_0000_0000_0000;
array[60601] <= 16'b0000_0000_0000_0000;
array[60602] <= 16'b0000_0000_0000_0000;
array[60603] <= 16'b0000_0000_0000_0000;
array[60604] <= 16'b0000_0000_0000_0000;
array[60605] <= 16'b0000_0000_0000_0000;
array[60606] <= 16'b0000_0000_0000_0000;
array[60607] <= 16'b0000_0000_0000_0000;
array[60608] <= 16'b0000_0000_0000_0000;
array[60609] <= 16'b0000_0000_0000_0000;
array[60610] <= 16'b0000_0000_0000_0000;
array[60611] <= 16'b0000_0000_0000_0000;
array[60612] <= 16'b0000_0000_0000_0000;
array[60613] <= 16'b0000_0000_0000_0000;
array[60614] <= 16'b0000_0000_0000_0000;
array[60615] <= 16'b0000_0000_0000_0000;
array[60616] <= 16'b0000_0000_0000_0000;
array[60617] <= 16'b0000_0000_0000_0000;
array[60618] <= 16'b0000_0000_0000_0000;
array[60619] <= 16'b0000_0000_0000_0000;
array[60620] <= 16'b0000_0000_0000_0000;
array[60621] <= 16'b0000_0000_0000_0000;
array[60622] <= 16'b0000_0000_0000_0000;
array[60623] <= 16'b0000_0000_0000_0000;
array[60624] <= 16'b0000_0000_0000_0000;
array[60625] <= 16'b0000_0000_0000_0000;
array[60626] <= 16'b0000_0000_0000_0000;
array[60627] <= 16'b0000_0000_0000_0000;
array[60628] <= 16'b0000_0000_0000_0000;
array[60629] <= 16'b0000_0000_0000_0000;
array[60630] <= 16'b0000_0000_0000_0000;
array[60631] <= 16'b0000_0000_0000_0000;
array[60632] <= 16'b0000_0000_0000_0000;
array[60633] <= 16'b0000_0000_0000_0000;
array[60634] <= 16'b0000_0000_0000_0000;
array[60635] <= 16'b0000_0000_0000_0000;
array[60636] <= 16'b0000_0000_0000_0000;
array[60637] <= 16'b0000_0000_0000_0000;
array[60638] <= 16'b0000_0000_0000_0000;
array[60639] <= 16'b0000_0000_0000_0000;
array[60640] <= 16'b0000_0000_0000_0000;
array[60641] <= 16'b0000_0000_0000_0000;
array[60642] <= 16'b0000_0000_0000_0000;
array[60643] <= 16'b0000_0000_0000_0000;
array[60644] <= 16'b0000_0000_0000_0000;
array[60645] <= 16'b0000_0000_0000_0000;
array[60646] <= 16'b0000_0000_0000_0000;
array[60647] <= 16'b0000_0000_0000_0000;
array[60648] <= 16'b0000_0000_0000_0000;
array[60649] <= 16'b0000_0000_0000_0000;
array[60650] <= 16'b0000_0000_0000_0000;
array[60651] <= 16'b0000_0000_0000_0000;
array[60652] <= 16'b0000_0000_0000_0000;
array[60653] <= 16'b0000_0000_0000_0000;
array[60654] <= 16'b0000_0000_0000_0000;
array[60655] <= 16'b0000_0000_0000_0000;
array[60656] <= 16'b0000_0000_0000_0000;
array[60657] <= 16'b0000_0000_0000_0000;
array[60658] <= 16'b0000_0000_0000_0000;
array[60659] <= 16'b0000_0000_0000_0000;
array[60660] <= 16'b0000_0000_0000_0000;
array[60661] <= 16'b0000_0000_0000_0000;
array[60662] <= 16'b0000_0000_0000_0000;
array[60663] <= 16'b0000_0000_0000_0000;
array[60664] <= 16'b0000_0000_0000_0000;
array[60665] <= 16'b0000_0000_0000_0000;
array[60666] <= 16'b0000_0000_0000_0000;
array[60667] <= 16'b0000_0000_0000_0000;
array[60668] <= 16'b0000_0000_0000_0000;
array[60669] <= 16'b0000_0000_0000_0000;
array[60670] <= 16'b0000_0000_0000_0000;
array[60671] <= 16'b0000_0000_0000_0000;
array[60672] <= 16'b0000_0000_0000_0000;
array[60673] <= 16'b0000_0000_0000_0000;
array[60674] <= 16'b0000_0000_0000_0000;
array[60675] <= 16'b0000_0000_0000_0000;
array[60676] <= 16'b0000_0000_0000_0000;
array[60677] <= 16'b0000_0000_0000_0000;
array[60678] <= 16'b0000_0000_0000_0000;
array[60679] <= 16'b0000_0000_0000_0000;
array[60680] <= 16'b0000_0000_0000_0000;
array[60681] <= 16'b0000_0000_0000_0000;
array[60682] <= 16'b0000_0000_0000_0000;
array[60683] <= 16'b0000_0000_0000_0000;
array[60684] <= 16'b0000_0000_0000_0000;
array[60685] <= 16'b0000_0000_0000_0000;
array[60686] <= 16'b0000_0000_0000_0000;
array[60687] <= 16'b0000_0000_0000_0000;
array[60688] <= 16'b0000_0000_0000_0000;
array[60689] <= 16'b0000_0000_0000_0000;
array[60690] <= 16'b0000_0000_0000_0000;
array[60691] <= 16'b0000_0000_0000_0000;
array[60692] <= 16'b0000_0000_0000_0000;
array[60693] <= 16'b0000_0000_0000_0000;
array[60694] <= 16'b0000_0000_0000_0000;
array[60695] <= 16'b0000_0000_0000_0000;
array[60696] <= 16'b0000_0000_0000_0000;
array[60697] <= 16'b0000_0000_0000_0000;
array[60698] <= 16'b0000_0000_0000_0000;
array[60699] <= 16'b0000_0000_0000_0000;
array[60700] <= 16'b0000_0000_0000_0000;
array[60701] <= 16'b0000_0000_0000_0000;
array[60702] <= 16'b0000_0000_0000_0000;
array[60703] <= 16'b0000_0000_0000_0000;
array[60704] <= 16'b0000_0000_0000_0000;
array[60705] <= 16'b0000_0000_0000_0000;
array[60706] <= 16'b0000_0000_0000_0000;
array[60707] <= 16'b0000_0000_0000_0000;
array[60708] <= 16'b0000_0000_0000_0000;
array[60709] <= 16'b0000_0000_0000_0000;
array[60710] <= 16'b0000_0000_0000_0000;
array[60711] <= 16'b0000_0000_0000_0000;
array[60712] <= 16'b0000_0000_0000_0000;
array[60713] <= 16'b0000_0000_0000_0000;
array[60714] <= 16'b0000_0000_0000_0000;
array[60715] <= 16'b0000_0000_0000_0000;
array[60716] <= 16'b0000_0000_0000_0000;
array[60717] <= 16'b0000_0000_0000_0000;
array[60718] <= 16'b0000_0000_0000_0000;
array[60719] <= 16'b0000_0000_0000_0000;
array[60720] <= 16'b0000_0000_0000_0000;
array[60721] <= 16'b0000_0000_0000_0000;
array[60722] <= 16'b0000_0000_0000_0000;
array[60723] <= 16'b0000_0000_0000_0000;
array[60724] <= 16'b0000_0000_0000_0000;
array[60725] <= 16'b0000_0000_0000_0000;
array[60726] <= 16'b0000_0000_0000_0000;
array[60727] <= 16'b0000_0000_0000_0000;
array[60728] <= 16'b0000_0000_0000_0000;
array[60729] <= 16'b0000_0000_0000_0000;
array[60730] <= 16'b0000_0000_0000_0000;
array[60731] <= 16'b0000_0000_0000_0000;
array[60732] <= 16'b0000_0000_0000_0000;
array[60733] <= 16'b0000_0000_0000_0000;
array[60734] <= 16'b0000_0000_0000_0000;
array[60735] <= 16'b0000_0000_0000_0000;
array[60736] <= 16'b0000_0000_0000_0000;
array[60737] <= 16'b0000_0000_0000_0000;
array[60738] <= 16'b0000_0000_0000_0000;
array[60739] <= 16'b0000_0000_0000_0000;
array[60740] <= 16'b0000_0000_0000_0000;
array[60741] <= 16'b0000_0000_0000_0000;
array[60742] <= 16'b0000_0000_0000_0000;
array[60743] <= 16'b0000_0000_0000_0000;
array[60744] <= 16'b0000_0000_0000_0000;
array[60745] <= 16'b0000_0000_0000_0000;
array[60746] <= 16'b0000_0000_0000_0000;
array[60747] <= 16'b0000_0000_0000_0000;
array[60748] <= 16'b0000_0000_0000_0000;
array[60749] <= 16'b0000_0000_0000_0000;
array[60750] <= 16'b0000_0000_0000_0000;
array[60751] <= 16'b0000_0000_0000_0000;
array[60752] <= 16'b0000_0000_0000_0000;
array[60753] <= 16'b0000_0000_0000_0000;
array[60754] <= 16'b0000_0000_0000_0000;
array[60755] <= 16'b0000_0000_0000_0000;
array[60756] <= 16'b0000_0000_0000_0000;
array[60757] <= 16'b0000_0000_0000_0000;
array[60758] <= 16'b0000_0000_0000_0000;
array[60759] <= 16'b0000_0000_0000_0000;
array[60760] <= 16'b0000_0000_0000_0000;
array[60761] <= 16'b0000_0000_0000_0000;
array[60762] <= 16'b0000_0000_0000_0000;
array[60763] <= 16'b0000_0000_0000_0000;
array[60764] <= 16'b0000_0000_0000_0000;
array[60765] <= 16'b0000_0000_0000_0000;
array[60766] <= 16'b0000_0000_0000_0000;
array[60767] <= 16'b0000_0000_0000_0000;
array[60768] <= 16'b0000_0000_0000_0000;
array[60769] <= 16'b0000_0000_0000_0000;
array[60770] <= 16'b0000_0000_0000_0000;
array[60771] <= 16'b0000_0000_0000_0000;
array[60772] <= 16'b0000_0000_0000_0000;
array[60773] <= 16'b0000_0000_0000_0000;
array[60774] <= 16'b0000_0000_0000_0000;
array[60775] <= 16'b0000_0000_0000_0000;
array[60776] <= 16'b0000_0000_0000_0000;
array[60777] <= 16'b0000_0000_0000_0000;
array[60778] <= 16'b0000_0000_0000_0000;
array[60779] <= 16'b0000_0000_0000_0000;
array[60780] <= 16'b0000_0000_0000_0000;
array[60781] <= 16'b0000_0000_0000_0000;
array[60782] <= 16'b0000_0000_0000_0000;
array[60783] <= 16'b0000_0000_0000_0000;
array[60784] <= 16'b0000_0000_0000_0000;
array[60785] <= 16'b0000_0000_0000_0000;
array[60786] <= 16'b0000_0000_0000_0000;
array[60787] <= 16'b0000_0000_0000_0000;
array[60788] <= 16'b0000_0000_0000_0000;
array[60789] <= 16'b0000_0000_0000_0000;
array[60790] <= 16'b0000_0000_0000_0000;
array[60791] <= 16'b0000_0000_0000_0000;
array[60792] <= 16'b0000_0000_0000_0000;
array[60793] <= 16'b0000_0000_0000_0000;
array[60794] <= 16'b0000_0000_0000_0000;
array[60795] <= 16'b0000_0000_0000_0000;
array[60796] <= 16'b0000_0000_0000_0000;
array[60797] <= 16'b0000_0000_0000_0000;
array[60798] <= 16'b0000_0000_0000_0000;
array[60799] <= 16'b0000_0000_0000_0000;
array[60800] <= 16'b0000_0000_0000_0000;
array[60801] <= 16'b0000_0000_0000_0000;
array[60802] <= 16'b0000_0000_0000_0000;
array[60803] <= 16'b0000_0000_0000_0000;
array[60804] <= 16'b0000_0000_0000_0000;
array[60805] <= 16'b0000_0000_0000_0000;
array[60806] <= 16'b0000_0000_0000_0000;
array[60807] <= 16'b0000_0000_0000_0000;
array[60808] <= 16'b0000_0000_0000_0000;
array[60809] <= 16'b0000_0000_0000_0000;
array[60810] <= 16'b0000_0000_0000_0000;
array[60811] <= 16'b0000_0000_0000_0000;
array[60812] <= 16'b0000_0000_0000_0000;
array[60813] <= 16'b0000_0000_0000_0000;
array[60814] <= 16'b0000_0000_0000_0000;
array[60815] <= 16'b0000_0000_0000_0000;
array[60816] <= 16'b0000_0000_0000_0000;
array[60817] <= 16'b0000_0000_0000_0000;
array[60818] <= 16'b0000_0000_0000_0000;
array[60819] <= 16'b0000_0000_0000_0000;
array[60820] <= 16'b0000_0000_0000_0000;
array[60821] <= 16'b0000_0000_0000_0000;
array[60822] <= 16'b0000_0000_0000_0000;
array[60823] <= 16'b0000_0000_0000_0000;
array[60824] <= 16'b0000_0000_0000_0000;
array[60825] <= 16'b0000_0000_0000_0000;
array[60826] <= 16'b0000_0000_0000_0000;
array[60827] <= 16'b0000_0000_0000_0000;
array[60828] <= 16'b0000_0000_0000_0000;
array[60829] <= 16'b0000_0000_0000_0000;
array[60830] <= 16'b0000_0000_0000_0000;
array[60831] <= 16'b0000_0000_0000_0000;
array[60832] <= 16'b0000_0000_0000_0000;
array[60833] <= 16'b0000_0000_0000_0000;
array[60834] <= 16'b0000_0000_0000_0000;
array[60835] <= 16'b0000_0000_0000_0000;
array[60836] <= 16'b0000_0000_0000_0000;
array[60837] <= 16'b0000_0000_0000_0000;
array[60838] <= 16'b0000_0000_0000_0000;
array[60839] <= 16'b0000_0000_0000_0000;
array[60840] <= 16'b0000_0000_0000_0000;
array[60841] <= 16'b0000_0000_0000_0000;
array[60842] <= 16'b0000_0000_0000_0000;
array[60843] <= 16'b0000_0000_0000_0000;
array[60844] <= 16'b0000_0000_0000_0000;
array[60845] <= 16'b0000_0000_0000_0000;
array[60846] <= 16'b0000_0000_0000_0000;
array[60847] <= 16'b0000_0000_0000_0000;
array[60848] <= 16'b0000_0000_0000_0000;
array[60849] <= 16'b0000_0000_0000_0000;
array[60850] <= 16'b0000_0000_0000_0000;
array[60851] <= 16'b0000_0000_0000_0000;
array[60852] <= 16'b0000_0000_0000_0000;
array[60853] <= 16'b0000_0000_0000_0000;
array[60854] <= 16'b0000_0000_0000_0000;
array[60855] <= 16'b0000_0000_0000_0000;
array[60856] <= 16'b0000_0000_0000_0000;
array[60857] <= 16'b0000_0000_0000_0000;
array[60858] <= 16'b0000_0000_0000_0000;
array[60859] <= 16'b0000_0000_0000_0000;
array[60860] <= 16'b0000_0000_0000_0000;
array[60861] <= 16'b0000_0000_0000_0000;
array[60862] <= 16'b0000_0000_0000_0000;
array[60863] <= 16'b0000_0000_0000_0000;
array[60864] <= 16'b0000_0000_0000_0000;
array[60865] <= 16'b0000_0000_0000_0000;
array[60866] <= 16'b0000_0000_0000_0000;
array[60867] <= 16'b0000_0000_0000_0000;
array[60868] <= 16'b0000_0000_0000_0000;
array[60869] <= 16'b0000_0000_0000_0000;
array[60870] <= 16'b0000_0000_0000_0000;
array[60871] <= 16'b0000_0000_0000_0000;
array[60872] <= 16'b0000_0000_0000_0000;
array[60873] <= 16'b0000_0000_0000_0000;
array[60874] <= 16'b0000_0000_0000_0000;
array[60875] <= 16'b0000_0000_0000_0000;
array[60876] <= 16'b0000_0000_0000_0000;
array[60877] <= 16'b0000_0000_0000_0000;
array[60878] <= 16'b0000_0000_0000_0000;
array[60879] <= 16'b0000_0000_0000_0000;
array[60880] <= 16'b0000_0000_0000_0000;
array[60881] <= 16'b0000_0000_0000_0000;
array[60882] <= 16'b0000_0000_0000_0000;
array[60883] <= 16'b0000_0000_0000_0000;
array[60884] <= 16'b0000_0000_0000_0000;
array[60885] <= 16'b0000_0000_0000_0000;
array[60886] <= 16'b0000_0000_0000_0000;
array[60887] <= 16'b0000_0000_0000_0000;
array[60888] <= 16'b0000_0000_0000_0000;
array[60889] <= 16'b0000_0000_0000_0000;
array[60890] <= 16'b0000_0000_0000_0000;
array[60891] <= 16'b0000_0000_0000_0000;
array[60892] <= 16'b0000_0000_0000_0000;
array[60893] <= 16'b0000_0000_0000_0000;
array[60894] <= 16'b0000_0000_0000_0000;
array[60895] <= 16'b0000_0000_0000_0000;
array[60896] <= 16'b0000_0000_0000_0000;
array[60897] <= 16'b0000_0000_0000_0000;
array[60898] <= 16'b0000_0000_0000_0000;
array[60899] <= 16'b0000_0000_0000_0000;
array[60900] <= 16'b0000_0000_0000_0000;
array[60901] <= 16'b0000_0000_0000_0000;
array[60902] <= 16'b0000_0000_0000_0000;
array[60903] <= 16'b0000_0000_0000_0000;
array[60904] <= 16'b0000_0000_0000_0000;
array[60905] <= 16'b0000_0000_0000_0000;
array[60906] <= 16'b0000_0000_0000_0000;
array[60907] <= 16'b0000_0000_0000_0000;
array[60908] <= 16'b0000_0000_0000_0000;
array[60909] <= 16'b0000_0000_0000_0000;
array[60910] <= 16'b0000_0000_0000_0000;
array[60911] <= 16'b0000_0000_0000_0000;
array[60912] <= 16'b0000_0000_0000_0000;
array[60913] <= 16'b0000_0000_0000_0000;
array[60914] <= 16'b0000_0000_0000_0000;
array[60915] <= 16'b0000_0000_0000_0000;
array[60916] <= 16'b0000_0000_0000_0000;
array[60917] <= 16'b0000_0000_0000_0000;
array[60918] <= 16'b0000_0000_0000_0000;
array[60919] <= 16'b0000_0000_0000_0000;
array[60920] <= 16'b0000_0000_0000_0000;
array[60921] <= 16'b0000_0000_0000_0000;
array[60922] <= 16'b0000_0000_0000_0000;
array[60923] <= 16'b0000_0000_0000_0000;
array[60924] <= 16'b0000_0000_0000_0000;
array[60925] <= 16'b0000_0000_0000_0000;
array[60926] <= 16'b0000_0000_0000_0000;
array[60927] <= 16'b0000_0000_0000_0000;
array[60928] <= 16'b0000_0000_0000_0000;
array[60929] <= 16'b0000_0000_0000_0000;
array[60930] <= 16'b0000_0000_0000_0000;
array[60931] <= 16'b0000_0000_0000_0000;
array[60932] <= 16'b0000_0000_0000_0000;
array[60933] <= 16'b0000_0000_0000_0000;
array[60934] <= 16'b0000_0000_0000_0000;
array[60935] <= 16'b0000_0000_0000_0000;
array[60936] <= 16'b0000_0000_0000_0000;
array[60937] <= 16'b0000_0000_0000_0000;
array[60938] <= 16'b0000_0000_0000_0000;
array[60939] <= 16'b0000_0000_0000_0000;
array[60940] <= 16'b0000_0000_0000_0000;
array[60941] <= 16'b0000_0000_0000_0000;
array[60942] <= 16'b0000_0000_0000_0000;
array[60943] <= 16'b0000_0000_0000_0000;
array[60944] <= 16'b0000_0000_0000_0000;
array[60945] <= 16'b0000_0000_0000_0000;
array[60946] <= 16'b0000_0000_0000_0000;
array[60947] <= 16'b0000_0000_0000_0000;
array[60948] <= 16'b0000_0000_0000_0000;
array[60949] <= 16'b0000_0000_0000_0000;
array[60950] <= 16'b0000_0000_0000_0000;
array[60951] <= 16'b0000_0000_0000_0000;
array[60952] <= 16'b0000_0000_0000_0000;
array[60953] <= 16'b0000_0000_0000_0000;
array[60954] <= 16'b0000_0000_0000_0000;
array[60955] <= 16'b0000_0000_0000_0000;
array[60956] <= 16'b0000_0000_0000_0000;
array[60957] <= 16'b0000_0000_0000_0000;
array[60958] <= 16'b0000_0000_0000_0000;
array[60959] <= 16'b0000_0000_0000_0000;
array[60960] <= 16'b0000_0000_0000_0000;
array[60961] <= 16'b0000_0000_0000_0000;
array[60962] <= 16'b0000_0000_0000_0000;
array[60963] <= 16'b0000_0000_0000_0000;
array[60964] <= 16'b0000_0000_0000_0000;
array[60965] <= 16'b0000_0000_0000_0000;
array[60966] <= 16'b0000_0000_0000_0000;
array[60967] <= 16'b0000_0000_0000_0000;
array[60968] <= 16'b0000_0000_0000_0000;
array[60969] <= 16'b0000_0000_0000_0000;
array[60970] <= 16'b0000_0000_0000_0000;
array[60971] <= 16'b0000_0000_0000_0000;
array[60972] <= 16'b0000_0000_0000_0000;
array[60973] <= 16'b0000_0000_0000_0000;
array[60974] <= 16'b0000_0000_0000_0000;
array[60975] <= 16'b0000_0000_0000_0000;
array[60976] <= 16'b0000_0000_0000_0000;
array[60977] <= 16'b0000_0000_0000_0000;
array[60978] <= 16'b0000_0000_0000_0000;
array[60979] <= 16'b0000_0000_0000_0000;
array[60980] <= 16'b0000_0000_0000_0000;
array[60981] <= 16'b0000_0000_0000_0000;
array[60982] <= 16'b0000_0000_0000_0000;
array[60983] <= 16'b0000_0000_0000_0000;
array[60984] <= 16'b0000_0000_0000_0000;
array[60985] <= 16'b0000_0000_0000_0000;
array[60986] <= 16'b0000_0000_0000_0000;
array[60987] <= 16'b0000_0000_0000_0000;
array[60988] <= 16'b0000_0000_0000_0000;
array[60989] <= 16'b0000_0000_0000_0000;
array[60990] <= 16'b0000_0000_0000_0000;
array[60991] <= 16'b0000_0000_0000_0000;
array[60992] <= 16'b0000_0000_0000_0000;
array[60993] <= 16'b0000_0000_0000_0000;
array[60994] <= 16'b0000_0000_0000_0000;
array[60995] <= 16'b0000_0000_0000_0000;
array[60996] <= 16'b0000_0000_0000_0000;
array[60997] <= 16'b0000_0000_0000_0000;
array[60998] <= 16'b0000_0000_0000_0000;
array[60999] <= 16'b0000_0000_0000_0000;
array[61000] <= 16'b0000_0000_0000_0000;
array[61001] <= 16'b0000_0000_0000_0000;
array[61002] <= 16'b0000_0000_0000_0000;
array[61003] <= 16'b0000_0000_0000_0000;
array[61004] <= 16'b0000_0000_0000_0000;
array[61005] <= 16'b0000_0000_0000_0000;
array[61006] <= 16'b0000_0000_0000_0000;
array[61007] <= 16'b0000_0000_0000_0000;
array[61008] <= 16'b0000_0000_0000_0000;
array[61009] <= 16'b0000_0000_0000_0000;
array[61010] <= 16'b0000_0000_0000_0000;
array[61011] <= 16'b0000_0000_0000_0000;
array[61012] <= 16'b0000_0000_0000_0000;
array[61013] <= 16'b0000_0000_0000_0000;
array[61014] <= 16'b0000_0000_0000_0000;
array[61015] <= 16'b0000_0000_0000_0000;
array[61016] <= 16'b0000_0000_0000_0000;
array[61017] <= 16'b0000_0000_0000_0000;
array[61018] <= 16'b0000_0000_0000_0000;
array[61019] <= 16'b0000_0000_0000_0000;
array[61020] <= 16'b0000_0000_0000_0000;
array[61021] <= 16'b0000_0000_0000_0000;
array[61022] <= 16'b0000_0000_0000_0000;
array[61023] <= 16'b0000_0000_0000_0000;
array[61024] <= 16'b0000_0000_0000_0000;
array[61025] <= 16'b0000_0000_0000_0000;
array[61026] <= 16'b0000_0000_0000_0000;
array[61027] <= 16'b0000_0000_0000_0000;
array[61028] <= 16'b0000_0000_0000_0000;
array[61029] <= 16'b0000_0000_0000_0000;
array[61030] <= 16'b0000_0000_0000_0000;
array[61031] <= 16'b0000_0000_0000_0000;
array[61032] <= 16'b0000_0000_0000_0000;
array[61033] <= 16'b0000_0000_0000_0000;
array[61034] <= 16'b0000_0000_0000_0000;
array[61035] <= 16'b0000_0000_0000_0000;
array[61036] <= 16'b0000_0000_0000_0000;
array[61037] <= 16'b0000_0000_0000_0000;
array[61038] <= 16'b0000_0000_0000_0000;
array[61039] <= 16'b0000_0000_0000_0000;
array[61040] <= 16'b0000_0000_0000_0000;
array[61041] <= 16'b0000_0000_0000_0000;
array[61042] <= 16'b0000_0000_0000_0000;
array[61043] <= 16'b0000_0000_0000_0000;
array[61044] <= 16'b0000_0000_0000_0000;
array[61045] <= 16'b0000_0000_0000_0000;
array[61046] <= 16'b0000_0000_0000_0000;
array[61047] <= 16'b0000_0000_0000_0000;
array[61048] <= 16'b0000_0000_0000_0000;
array[61049] <= 16'b0000_0000_0000_0000;
array[61050] <= 16'b0000_0000_0000_0000;
array[61051] <= 16'b0000_0000_0000_0000;
array[61052] <= 16'b0000_0000_0000_0000;
array[61053] <= 16'b0000_0000_0000_0000;
array[61054] <= 16'b0000_0000_0000_0000;
array[61055] <= 16'b0000_0000_0000_0000;
array[61056] <= 16'b0000_0000_0000_0000;
array[61057] <= 16'b0000_0000_0000_0000;
array[61058] <= 16'b0000_0000_0000_0000;
array[61059] <= 16'b0000_0000_0000_0000;
array[61060] <= 16'b0000_0000_0000_0000;
array[61061] <= 16'b0000_0000_0000_0000;
array[61062] <= 16'b0000_0000_0000_0000;
array[61063] <= 16'b0000_0000_0000_0000;
array[61064] <= 16'b0000_0000_0000_0000;
array[61065] <= 16'b0000_0000_0000_0000;
array[61066] <= 16'b0000_0000_0000_0000;
array[61067] <= 16'b0000_0000_0000_0000;
array[61068] <= 16'b0000_0000_0000_0000;
array[61069] <= 16'b0000_0000_0000_0000;
array[61070] <= 16'b0000_0000_0000_0000;
array[61071] <= 16'b0000_0000_0000_0000;
array[61072] <= 16'b0000_0000_0000_0000;
array[61073] <= 16'b0000_0000_0000_0000;
array[61074] <= 16'b0000_0000_0000_0000;
array[61075] <= 16'b0000_0000_0000_0000;
array[61076] <= 16'b0000_0000_0000_0000;
array[61077] <= 16'b0000_0000_0000_0000;
array[61078] <= 16'b0000_0000_0000_0000;
array[61079] <= 16'b0000_0000_0000_0000;
array[61080] <= 16'b0000_0000_0000_0000;
array[61081] <= 16'b0000_0000_0000_0000;
array[61082] <= 16'b0000_0000_0000_0000;
array[61083] <= 16'b0000_0000_0000_0000;
array[61084] <= 16'b0000_0000_0000_0000;
array[61085] <= 16'b0000_0000_0000_0000;
array[61086] <= 16'b0000_0000_0000_0000;
array[61087] <= 16'b0000_0000_0000_0000;
array[61088] <= 16'b0000_0000_0000_0000;
array[61089] <= 16'b0000_0000_0000_0000;
array[61090] <= 16'b0000_0000_0000_0000;
array[61091] <= 16'b0000_0000_0000_0000;
array[61092] <= 16'b0000_0000_0000_0000;
array[61093] <= 16'b0000_0000_0000_0000;
array[61094] <= 16'b0000_0000_0000_0000;
array[61095] <= 16'b0000_0000_0000_0000;
array[61096] <= 16'b0000_0000_0000_0000;
array[61097] <= 16'b0000_0000_0000_0000;
array[61098] <= 16'b0000_0000_0000_0000;
array[61099] <= 16'b0000_0000_0000_0000;
array[61100] <= 16'b0000_0000_0000_0000;
array[61101] <= 16'b0000_0000_0000_0000;
array[61102] <= 16'b0000_0000_0000_0000;
array[61103] <= 16'b0000_0000_0000_0000;
array[61104] <= 16'b0000_0000_0000_0000;
array[61105] <= 16'b0000_0000_0000_0000;
array[61106] <= 16'b0000_0000_0000_0000;
array[61107] <= 16'b0000_0000_0000_0000;
array[61108] <= 16'b0000_0000_0000_0000;
array[61109] <= 16'b0000_0000_0000_0000;
array[61110] <= 16'b0000_0000_0000_0000;
array[61111] <= 16'b0000_0000_0000_0000;
array[61112] <= 16'b0000_0000_0000_0000;
array[61113] <= 16'b0000_0000_0000_0000;
array[61114] <= 16'b0000_0000_0000_0000;
array[61115] <= 16'b0000_0000_0000_0000;
array[61116] <= 16'b0000_0000_0000_0000;
array[61117] <= 16'b0000_0000_0000_0000;
array[61118] <= 16'b0000_0000_0000_0000;
array[61119] <= 16'b0000_0000_0000_0000;
array[61120] <= 16'b0000_0000_0000_0000;
array[61121] <= 16'b0000_0000_0000_0000;
array[61122] <= 16'b0000_0000_0000_0000;
array[61123] <= 16'b0000_0000_0000_0000;
array[61124] <= 16'b0000_0000_0000_0000;
array[61125] <= 16'b0000_0000_0000_0000;
array[61126] <= 16'b0000_0000_0000_0000;
array[61127] <= 16'b0000_0000_0000_0000;
array[61128] <= 16'b0000_0000_0000_0000;
array[61129] <= 16'b0000_0000_0000_0000;
array[61130] <= 16'b0000_0000_0000_0000;
array[61131] <= 16'b0000_0000_0000_0000;
array[61132] <= 16'b0000_0000_0000_0000;
array[61133] <= 16'b0000_0000_0000_0000;
array[61134] <= 16'b0000_0000_0000_0000;
array[61135] <= 16'b0000_0000_0000_0000;
array[61136] <= 16'b0000_0000_0000_0000;
array[61137] <= 16'b0000_0000_0000_0000;
array[61138] <= 16'b0000_0000_0000_0000;
array[61139] <= 16'b0000_0000_0000_0000;
array[61140] <= 16'b0000_0000_0000_0000;
array[61141] <= 16'b0000_0000_0000_0000;
array[61142] <= 16'b0000_0000_0000_0000;
array[61143] <= 16'b0000_0000_0000_0000;
array[61144] <= 16'b0000_0000_0000_0000;
array[61145] <= 16'b0000_0000_0000_0000;
array[61146] <= 16'b0000_0000_0000_0000;
array[61147] <= 16'b0000_0000_0000_0000;
array[61148] <= 16'b0000_0000_0000_0000;
array[61149] <= 16'b0000_0000_0000_0000;
array[61150] <= 16'b0000_0000_0000_0000;
array[61151] <= 16'b0000_0000_0000_0000;
array[61152] <= 16'b0000_0000_0000_0000;
array[61153] <= 16'b0000_0000_0000_0000;
array[61154] <= 16'b0000_0000_0000_0000;
array[61155] <= 16'b0000_0000_0000_0000;
array[61156] <= 16'b0000_0000_0000_0000;
array[61157] <= 16'b0000_0000_0000_0000;
array[61158] <= 16'b0000_0000_0000_0000;
array[61159] <= 16'b0000_0000_0000_0000;
array[61160] <= 16'b0000_0000_0000_0000;
array[61161] <= 16'b0000_0000_0000_0000;
array[61162] <= 16'b0000_0000_0000_0000;
array[61163] <= 16'b0000_0000_0000_0000;
array[61164] <= 16'b0000_0000_0000_0000;
array[61165] <= 16'b0000_0000_0000_0000;
array[61166] <= 16'b0000_0000_0000_0000;
array[61167] <= 16'b0000_0000_0000_0000;
array[61168] <= 16'b0000_0000_0000_0000;
array[61169] <= 16'b0000_0000_0000_0000;
array[61170] <= 16'b0000_0000_0000_0000;
array[61171] <= 16'b0000_0000_0000_0000;
array[61172] <= 16'b0000_0000_0000_0000;
array[61173] <= 16'b0000_0000_0000_0000;
array[61174] <= 16'b0000_0000_0000_0000;
array[61175] <= 16'b0000_0000_0000_0000;
array[61176] <= 16'b0000_0000_0000_0000;
array[61177] <= 16'b0000_0000_0000_0000;
array[61178] <= 16'b0000_0000_0000_0000;
array[61179] <= 16'b0000_0000_0000_0000;
array[61180] <= 16'b0000_0000_0000_0000;
array[61181] <= 16'b0000_0000_0000_0000;
array[61182] <= 16'b0000_0000_0000_0000;
array[61183] <= 16'b0000_0000_0000_0000;
array[61184] <= 16'b0000_0000_0000_0000;
array[61185] <= 16'b0000_0000_0000_0000;
array[61186] <= 16'b0000_0000_0000_0000;
array[61187] <= 16'b0000_0000_0000_0000;
array[61188] <= 16'b0000_0000_0000_0000;
array[61189] <= 16'b0000_0000_0000_0000;
array[61190] <= 16'b0000_0000_0000_0000;
array[61191] <= 16'b0000_0000_0000_0000;
array[61192] <= 16'b0000_0000_0000_0000;
array[61193] <= 16'b0000_0000_0000_0000;
array[61194] <= 16'b0000_0000_0000_0000;
array[61195] <= 16'b0000_0000_0000_0000;
array[61196] <= 16'b0000_0000_0000_0000;
array[61197] <= 16'b0000_0000_0000_0000;
array[61198] <= 16'b0000_0000_0000_0000;
array[61199] <= 16'b0000_0000_0000_0000;
array[61200] <= 16'b0000_0000_0000_0000;
array[61201] <= 16'b0000_0000_0000_0000;
array[61202] <= 16'b0000_0000_0000_0000;
array[61203] <= 16'b0000_0000_0000_0000;
array[61204] <= 16'b0000_0000_0000_0000;
array[61205] <= 16'b0000_0000_0000_0000;
array[61206] <= 16'b0000_0000_0000_0000;
array[61207] <= 16'b0000_0000_0000_0000;
array[61208] <= 16'b0000_0000_0000_0000;
array[61209] <= 16'b0000_0000_0000_0000;
array[61210] <= 16'b0000_0000_0000_0000;
array[61211] <= 16'b0000_0000_0000_0000;
array[61212] <= 16'b0000_0000_0000_0000;
array[61213] <= 16'b0000_0000_0000_0000;
array[61214] <= 16'b0000_0000_0000_0000;
array[61215] <= 16'b0000_0000_0000_0000;
array[61216] <= 16'b0000_0000_0000_0000;
array[61217] <= 16'b0000_0000_0000_0000;
array[61218] <= 16'b0000_0000_0000_0000;
array[61219] <= 16'b0000_0000_0000_0000;
array[61220] <= 16'b0000_0000_0000_0000;
array[61221] <= 16'b0000_0000_0000_0000;
array[61222] <= 16'b0000_0000_0000_0000;
array[61223] <= 16'b0000_0000_0000_0000;
array[61224] <= 16'b0000_0000_0000_0000;
array[61225] <= 16'b0000_0000_0000_0000;
array[61226] <= 16'b0000_0000_0000_0000;
array[61227] <= 16'b0000_0000_0000_0000;
array[61228] <= 16'b0000_0000_0000_0000;
array[61229] <= 16'b0000_0000_0000_0000;
array[61230] <= 16'b0000_0000_0000_0000;
array[61231] <= 16'b0000_0000_0000_0000;
array[61232] <= 16'b0000_0000_0000_0000;
array[61233] <= 16'b0000_0000_0000_0000;
array[61234] <= 16'b0000_0000_0000_0000;
array[61235] <= 16'b0000_0000_0000_0000;
array[61236] <= 16'b0000_0000_0000_0000;
array[61237] <= 16'b0000_0000_0000_0000;
array[61238] <= 16'b0000_0000_0000_0000;
array[61239] <= 16'b0000_0000_0000_0000;
array[61240] <= 16'b0000_0000_0000_0000;
array[61241] <= 16'b0000_0000_0000_0000;
array[61242] <= 16'b0000_0000_0000_0000;
array[61243] <= 16'b0000_0000_0000_0000;
array[61244] <= 16'b0000_0000_0000_0000;
array[61245] <= 16'b0000_0000_0000_0000;
array[61246] <= 16'b0000_0000_0000_0000;
array[61247] <= 16'b0000_0000_0000_0000;
array[61248] <= 16'b0000_0000_0000_0000;
array[61249] <= 16'b0000_0000_0000_0000;
array[61250] <= 16'b0000_0000_0000_0000;
array[61251] <= 16'b0000_0000_0000_0000;
array[61252] <= 16'b0000_0000_0000_0000;
array[61253] <= 16'b0000_0000_0000_0000;
array[61254] <= 16'b0000_0000_0000_0000;
array[61255] <= 16'b0000_0000_0000_0000;
array[61256] <= 16'b0000_0000_0000_0000;
array[61257] <= 16'b0000_0000_0000_0000;
array[61258] <= 16'b0000_0000_0000_0000;
array[61259] <= 16'b0000_0000_0000_0000;
array[61260] <= 16'b0000_0000_0000_0000;
array[61261] <= 16'b0000_0000_0000_0000;
array[61262] <= 16'b0000_0000_0000_0000;
array[61263] <= 16'b0000_0000_0000_0000;
array[61264] <= 16'b0000_0000_0000_0000;
array[61265] <= 16'b0000_0000_0000_0000;
array[61266] <= 16'b0000_0000_0000_0000;
array[61267] <= 16'b0000_0000_0000_0000;
array[61268] <= 16'b0000_0000_0000_0000;
array[61269] <= 16'b0000_0000_0000_0000;
array[61270] <= 16'b0000_0000_0000_0000;
array[61271] <= 16'b0000_0000_0000_0000;
array[61272] <= 16'b0000_0000_0000_0000;
array[61273] <= 16'b0000_0000_0000_0000;
array[61274] <= 16'b0000_0000_0000_0000;
array[61275] <= 16'b0000_0000_0000_0000;
array[61276] <= 16'b0000_0000_0000_0000;
array[61277] <= 16'b0000_0000_0000_0000;
array[61278] <= 16'b0000_0000_0000_0000;
array[61279] <= 16'b0000_0000_0000_0000;
array[61280] <= 16'b0000_0000_0000_0000;
array[61281] <= 16'b0000_0000_0000_0000;
array[61282] <= 16'b0000_0000_0000_0000;
array[61283] <= 16'b0000_0000_0000_0000;
array[61284] <= 16'b0000_0000_0000_0000;
array[61285] <= 16'b0000_0000_0000_0000;
array[61286] <= 16'b0000_0000_0000_0000;
array[61287] <= 16'b0000_0000_0000_0000;
array[61288] <= 16'b0000_0000_0000_0000;
array[61289] <= 16'b0000_0000_0000_0000;
array[61290] <= 16'b0000_0000_0000_0000;
array[61291] <= 16'b0000_0000_0000_0000;
array[61292] <= 16'b0000_0000_0000_0000;
array[61293] <= 16'b0000_0000_0000_0000;
array[61294] <= 16'b0000_0000_0000_0000;
array[61295] <= 16'b0000_0000_0000_0000;
array[61296] <= 16'b0000_0000_0000_0000;
array[61297] <= 16'b0000_0000_0000_0000;
array[61298] <= 16'b0000_0000_0000_0000;
array[61299] <= 16'b0000_0000_0000_0000;
array[61300] <= 16'b0000_0000_0000_0000;
array[61301] <= 16'b0000_0000_0000_0000;
array[61302] <= 16'b0000_0000_0000_0000;
array[61303] <= 16'b0000_0000_0000_0000;
array[61304] <= 16'b0000_0000_0000_0000;
array[61305] <= 16'b0000_0000_0000_0000;
array[61306] <= 16'b0000_0000_0000_0000;
array[61307] <= 16'b0000_0000_0000_0000;
array[61308] <= 16'b0000_0000_0000_0000;
array[61309] <= 16'b0000_0000_0000_0000;
array[61310] <= 16'b0000_0000_0000_0000;
array[61311] <= 16'b0000_0000_0000_0000;
array[61312] <= 16'b0000_0000_0000_0000;
array[61313] <= 16'b0000_0000_0000_0000;
array[61314] <= 16'b0000_0000_0000_0000;
array[61315] <= 16'b0000_0000_0000_0000;
array[61316] <= 16'b0000_0000_0000_0000;
array[61317] <= 16'b0000_0000_0000_0000;
array[61318] <= 16'b0000_0000_0000_0000;
array[61319] <= 16'b0000_0000_0000_0000;
array[61320] <= 16'b0000_0000_0000_0000;
array[61321] <= 16'b0000_0000_0000_0000;
array[61322] <= 16'b0000_0000_0000_0000;
array[61323] <= 16'b0000_0000_0000_0000;
array[61324] <= 16'b0000_0000_0000_0000;
array[61325] <= 16'b0000_0000_0000_0000;
array[61326] <= 16'b0000_0000_0000_0000;
array[61327] <= 16'b0000_0000_0000_0000;
array[61328] <= 16'b0000_0000_0000_0000;
array[61329] <= 16'b0000_0000_0000_0000;
array[61330] <= 16'b0000_0000_0000_0000;
array[61331] <= 16'b0000_0000_0000_0000;
array[61332] <= 16'b0000_0000_0000_0000;
array[61333] <= 16'b0000_0000_0000_0000;
array[61334] <= 16'b0000_0000_0000_0000;
array[61335] <= 16'b0000_0000_0000_0000;
array[61336] <= 16'b0000_0000_0000_0000;
array[61337] <= 16'b0000_0000_0000_0000;
array[61338] <= 16'b0000_0000_0000_0000;
array[61339] <= 16'b0000_0000_0000_0000;
array[61340] <= 16'b0000_0000_0000_0000;
array[61341] <= 16'b0000_0000_0000_0000;
array[61342] <= 16'b0000_0000_0000_0000;
array[61343] <= 16'b0000_0000_0000_0000;
array[61344] <= 16'b0000_0000_0000_0000;
array[61345] <= 16'b0000_0000_0000_0000;
array[61346] <= 16'b0000_0000_0000_0000;
array[61347] <= 16'b0000_0000_0000_0000;
array[61348] <= 16'b0000_0000_0000_0000;
array[61349] <= 16'b0000_0000_0000_0000;
array[61350] <= 16'b0000_0000_0000_0000;
array[61351] <= 16'b0000_0000_0000_0000;
array[61352] <= 16'b0000_0000_0000_0000;
array[61353] <= 16'b0000_0000_0000_0000;
array[61354] <= 16'b0000_0000_0000_0000;
array[61355] <= 16'b0000_0000_0000_0000;
array[61356] <= 16'b0000_0000_0000_0000;
array[61357] <= 16'b0000_0000_0000_0000;
array[61358] <= 16'b0000_0000_0000_0000;
array[61359] <= 16'b0000_0000_0000_0000;
array[61360] <= 16'b0000_0000_0000_0000;
array[61361] <= 16'b0000_0000_0000_0000;
array[61362] <= 16'b0000_0000_0000_0000;
array[61363] <= 16'b0000_0000_0000_0000;
array[61364] <= 16'b0000_0000_0000_0000;
array[61365] <= 16'b0000_0000_0000_0000;
array[61366] <= 16'b0000_0000_0000_0000;
array[61367] <= 16'b0000_0000_0000_0000;
array[61368] <= 16'b0000_0000_0000_0000;
array[61369] <= 16'b0000_0000_0000_0000;
array[61370] <= 16'b0000_0000_0000_0000;
array[61371] <= 16'b0000_0000_0000_0000;
array[61372] <= 16'b0000_0000_0000_0000;
array[61373] <= 16'b0000_0000_0000_0000;
array[61374] <= 16'b0000_0000_0000_0000;
array[61375] <= 16'b0000_0000_0000_0000;
array[61376] <= 16'b0000_0000_0000_0000;
array[61377] <= 16'b0000_0000_0000_0000;
array[61378] <= 16'b0000_0000_0000_0000;
array[61379] <= 16'b0000_0000_0000_0000;
array[61380] <= 16'b0000_0000_0000_0000;
array[61381] <= 16'b0000_0000_0000_0000;
array[61382] <= 16'b0000_0000_0000_0000;
array[61383] <= 16'b0000_0000_0000_0000;
array[61384] <= 16'b0000_0000_0000_0000;
array[61385] <= 16'b0000_0000_0000_0000;
array[61386] <= 16'b0000_0000_0000_0000;
array[61387] <= 16'b0000_0000_0000_0000;
array[61388] <= 16'b0000_0000_0000_0000;
array[61389] <= 16'b0000_0000_0000_0000;
array[61390] <= 16'b0000_0000_0000_0000;
array[61391] <= 16'b0000_0000_0000_0000;
array[61392] <= 16'b0000_0000_0000_0000;
array[61393] <= 16'b0000_0000_0000_0000;
array[61394] <= 16'b0000_0000_0000_0000;
array[61395] <= 16'b0000_0000_0000_0000;
array[61396] <= 16'b0000_0000_0000_0000;
array[61397] <= 16'b0000_0000_0000_0000;
array[61398] <= 16'b0000_0000_0000_0000;
array[61399] <= 16'b0000_0000_0000_0000;
array[61400] <= 16'b0000_0000_0000_0000;
array[61401] <= 16'b0000_0000_0000_0000;
array[61402] <= 16'b0000_0000_0000_0000;
array[61403] <= 16'b0000_0000_0000_0000;
array[61404] <= 16'b0000_0000_0000_0000;
array[61405] <= 16'b0000_0000_0000_0000;
array[61406] <= 16'b0000_0000_0000_0000;
array[61407] <= 16'b0000_0000_0000_0000;
array[61408] <= 16'b0000_0000_0000_0000;
array[61409] <= 16'b0000_0000_0000_0000;
array[61410] <= 16'b0000_0000_0000_0000;
array[61411] <= 16'b0000_0000_0000_0000;
array[61412] <= 16'b0000_0000_0000_0000;
array[61413] <= 16'b0000_0000_0000_0000;
array[61414] <= 16'b0000_0000_0000_0000;
array[61415] <= 16'b0000_0000_0000_0000;
array[61416] <= 16'b0000_0000_0000_0000;
array[61417] <= 16'b0000_0000_0000_0000;
array[61418] <= 16'b0000_0000_0000_0000;
array[61419] <= 16'b0000_0000_0000_0000;
array[61420] <= 16'b0000_0000_0000_0000;
array[61421] <= 16'b0000_0000_0000_0000;
array[61422] <= 16'b0000_0000_0000_0000;
array[61423] <= 16'b0000_0000_0000_0000;
array[61424] <= 16'b0000_0000_0000_0000;
array[61425] <= 16'b0000_0000_0000_0000;
array[61426] <= 16'b0000_0000_0000_0000;
array[61427] <= 16'b0000_0000_0000_0000;
array[61428] <= 16'b0000_0000_0000_0000;
array[61429] <= 16'b0000_0000_0000_0000;
array[61430] <= 16'b0000_0000_0000_0000;
array[61431] <= 16'b0000_0000_0000_0000;
array[61432] <= 16'b0000_0000_0000_0000;
array[61433] <= 16'b0000_0000_0000_0000;
array[61434] <= 16'b0000_0000_0000_0000;
array[61435] <= 16'b0000_0000_0000_0000;
array[61436] <= 16'b0000_0000_0000_0000;
array[61437] <= 16'b0000_0000_0000_0000;
array[61438] <= 16'b0000_0000_0000_0000;
array[61439] <= 16'b0000_0000_0000_0000;
array[61440] <= 16'b0000_0000_0000_0000;
array[61441] <= 16'b0000_0000_0000_0000;
array[61442] <= 16'b0000_0000_0000_0000;
array[61443] <= 16'b0000_0000_0000_0000;
array[61444] <= 16'b0000_0000_0000_0000;
array[61445] <= 16'b0000_0000_0000_0000;
array[61446] <= 16'b0000_0000_0000_0000;
array[61447] <= 16'b0000_0000_0000_0000;
array[61448] <= 16'b0000_0000_0000_0000;
array[61449] <= 16'b0000_0000_0000_0000;
array[61450] <= 16'b0000_0000_0000_0000;
array[61451] <= 16'b0000_0000_0000_0000;
array[61452] <= 16'b0000_0000_0000_0000;
array[61453] <= 16'b0000_0000_0000_0000;
array[61454] <= 16'b0000_0000_0000_0000;
array[61455] <= 16'b0000_0000_0000_0000;
array[61456] <= 16'b0000_0000_0000_0000;
array[61457] <= 16'b0000_0000_0000_0000;
array[61458] <= 16'b0000_0000_0000_0000;
array[61459] <= 16'b0000_0000_0000_0000;
array[61460] <= 16'b0000_0000_0000_0000;
array[61461] <= 16'b0000_0000_0000_0000;
array[61462] <= 16'b0000_0000_0000_0000;
array[61463] <= 16'b0000_0000_0000_0000;
array[61464] <= 16'b0000_0000_0000_0000;
array[61465] <= 16'b0000_0000_0000_0000;
array[61466] <= 16'b0000_0000_0000_0000;
array[61467] <= 16'b0000_0000_0000_0000;
array[61468] <= 16'b0000_0000_0000_0000;
array[61469] <= 16'b0000_0000_0000_0000;
array[61470] <= 16'b0000_0000_0000_0000;
array[61471] <= 16'b0000_0000_0000_0000;
array[61472] <= 16'b0000_0000_0000_0000;
array[61473] <= 16'b0000_0000_0000_0000;
array[61474] <= 16'b0000_0000_0000_0000;
array[61475] <= 16'b0000_0000_0000_0000;
array[61476] <= 16'b0000_0000_0000_0000;
array[61477] <= 16'b0000_0000_0000_0000;
array[61478] <= 16'b0000_0000_0000_0000;
array[61479] <= 16'b0000_0000_0000_0000;
array[61480] <= 16'b0000_0000_0000_0000;
array[61481] <= 16'b0000_0000_0000_0000;
array[61482] <= 16'b0000_0000_0000_0000;
array[61483] <= 16'b0000_0000_0000_0000;
array[61484] <= 16'b0000_0000_0000_0000;
array[61485] <= 16'b0000_0000_0000_0000;
array[61486] <= 16'b0000_0000_0000_0000;
array[61487] <= 16'b0000_0000_0000_0000;
array[61488] <= 16'b0000_0000_0000_0000;
array[61489] <= 16'b0000_0000_0000_0000;
array[61490] <= 16'b0000_0000_0000_0000;
array[61491] <= 16'b0000_0000_0000_0000;
array[61492] <= 16'b0000_0000_0000_0000;
array[61493] <= 16'b0000_0000_0000_0000;
array[61494] <= 16'b0000_0000_0000_0000;
array[61495] <= 16'b0000_0000_0000_0000;
array[61496] <= 16'b0000_0000_0000_0000;
array[61497] <= 16'b0000_0000_0000_0000;
array[61498] <= 16'b0000_0000_0000_0000;
array[61499] <= 16'b0000_0000_0000_0000;
array[61500] <= 16'b0000_0000_0000_0000;
array[61501] <= 16'b0000_0000_0000_0000;
array[61502] <= 16'b0000_0000_0000_0000;
array[61503] <= 16'b0000_0000_0000_0000;
array[61504] <= 16'b0000_0000_0000_0000;
array[61505] <= 16'b0000_0000_0000_0000;
array[61506] <= 16'b0000_0000_0000_0000;
array[61507] <= 16'b0000_0000_0000_0000;
array[61508] <= 16'b0000_0000_0000_0000;
array[61509] <= 16'b0000_0000_0000_0000;
array[61510] <= 16'b0000_0000_0000_0000;
array[61511] <= 16'b0000_0000_0000_0000;
array[61512] <= 16'b0000_0000_0000_0000;
array[61513] <= 16'b0000_0000_0000_0000;
array[61514] <= 16'b0000_0000_0000_0000;
array[61515] <= 16'b0000_0000_0000_0000;
array[61516] <= 16'b0000_0000_0000_0000;
array[61517] <= 16'b0000_0000_0000_0000;
array[61518] <= 16'b0000_0000_0000_0000;
array[61519] <= 16'b0000_0000_0000_0000;
array[61520] <= 16'b0000_0000_0000_0000;
array[61521] <= 16'b0000_0000_0000_0000;
array[61522] <= 16'b0000_0000_0000_0000;
array[61523] <= 16'b0000_0000_0000_0000;
array[61524] <= 16'b0000_0000_0000_0000;
array[61525] <= 16'b0000_0000_0000_0000;
array[61526] <= 16'b0000_0000_0000_0000;
array[61527] <= 16'b0000_0000_0000_0000;
array[61528] <= 16'b0000_0000_0000_0000;
array[61529] <= 16'b0000_0000_0000_0000;
array[61530] <= 16'b0000_0000_0000_0000;
array[61531] <= 16'b0000_0000_0000_0000;
array[61532] <= 16'b0000_0000_0000_0000;
array[61533] <= 16'b0000_0000_0000_0000;
array[61534] <= 16'b0000_0000_0000_0000;
array[61535] <= 16'b0000_0000_0000_0000;
array[61536] <= 16'b0000_0000_0000_0000;
array[61537] <= 16'b0000_0000_0000_0000;
array[61538] <= 16'b0000_0000_0000_0000;
array[61539] <= 16'b0000_0000_0000_0000;
array[61540] <= 16'b0000_0000_0000_0000;
array[61541] <= 16'b0000_0000_0000_0000;
array[61542] <= 16'b0000_0000_0000_0000;
array[61543] <= 16'b0000_0000_0000_0000;
array[61544] <= 16'b0000_0000_0000_0000;
array[61545] <= 16'b0000_0000_0000_0000;
array[61546] <= 16'b0000_0000_0000_0000;
array[61547] <= 16'b0000_0000_0000_0000;
array[61548] <= 16'b0000_0000_0000_0000;
array[61549] <= 16'b0000_0000_0000_0000;
array[61550] <= 16'b0000_0000_0000_0000;
array[61551] <= 16'b0000_0000_0000_0000;
array[61552] <= 16'b0000_0000_0000_0000;
array[61553] <= 16'b0000_0000_0000_0000;
array[61554] <= 16'b0000_0000_0000_0000;
array[61555] <= 16'b0000_0000_0000_0000;
array[61556] <= 16'b0000_0000_0000_0000;
array[61557] <= 16'b0000_0000_0000_0000;
array[61558] <= 16'b0000_0000_0000_0000;
array[61559] <= 16'b0000_0000_0000_0000;
array[61560] <= 16'b0000_0000_0000_0000;
array[61561] <= 16'b0000_0000_0000_0000;
array[61562] <= 16'b0000_0000_0000_0000;
array[61563] <= 16'b0000_0000_0000_0000;
array[61564] <= 16'b0000_0000_0000_0000;
array[61565] <= 16'b0000_0000_0000_0000;
array[61566] <= 16'b0000_0000_0000_0000;
array[61567] <= 16'b0000_0000_0000_0000;
array[61568] <= 16'b0000_0000_0000_0000;
array[61569] <= 16'b0000_0000_0000_0000;
array[61570] <= 16'b0000_0000_0000_0000;
array[61571] <= 16'b0000_0000_0000_0000;
array[61572] <= 16'b0000_0000_0000_0000;
array[61573] <= 16'b0000_0000_0000_0000;
array[61574] <= 16'b0000_0000_0000_0000;
array[61575] <= 16'b0000_0000_0000_0000;
array[61576] <= 16'b0000_0000_0000_0000;
array[61577] <= 16'b0000_0000_0000_0000;
array[61578] <= 16'b0000_0000_0000_0000;
array[61579] <= 16'b0000_0000_0000_0000;
array[61580] <= 16'b0000_0000_0000_0000;
array[61581] <= 16'b0000_0000_0000_0000;
array[61582] <= 16'b0000_0000_0000_0000;
array[61583] <= 16'b0000_0000_0000_0000;
array[61584] <= 16'b0000_0000_0000_0000;
array[61585] <= 16'b0000_0000_0000_0000;
array[61586] <= 16'b0000_0000_0000_0000;
array[61587] <= 16'b0000_0000_0000_0000;
array[61588] <= 16'b0000_0000_0000_0000;
array[61589] <= 16'b0000_0000_0000_0000;
array[61590] <= 16'b0000_0000_0000_0000;
array[61591] <= 16'b0000_0000_0000_0000;
array[61592] <= 16'b0000_0000_0000_0000;
array[61593] <= 16'b0000_0000_0000_0000;
array[61594] <= 16'b0000_0000_0000_0000;
array[61595] <= 16'b0000_0000_0000_0000;
array[61596] <= 16'b0000_0000_0000_0000;
array[61597] <= 16'b0000_0000_0000_0000;
array[61598] <= 16'b0000_0000_0000_0000;
array[61599] <= 16'b0000_0000_0000_0000;
array[61600] <= 16'b0000_0000_0000_0000;
array[61601] <= 16'b0000_0000_0000_0000;
array[61602] <= 16'b0000_0000_0000_0000;
array[61603] <= 16'b0000_0000_0000_0000;
array[61604] <= 16'b0000_0000_0000_0000;
array[61605] <= 16'b0000_0000_0000_0000;
array[61606] <= 16'b0000_0000_0000_0000;
array[61607] <= 16'b0000_0000_0000_0000;
array[61608] <= 16'b0000_0000_0000_0000;
array[61609] <= 16'b0000_0000_0000_0000;
array[61610] <= 16'b0000_0000_0000_0000;
array[61611] <= 16'b0000_0000_0000_0000;
array[61612] <= 16'b0000_0000_0000_0000;
array[61613] <= 16'b0000_0000_0000_0000;
array[61614] <= 16'b0000_0000_0000_0000;
array[61615] <= 16'b0000_0000_0000_0000;
array[61616] <= 16'b0000_0000_0000_0000;
array[61617] <= 16'b0000_0000_0000_0000;
array[61618] <= 16'b0000_0000_0000_0000;
array[61619] <= 16'b0000_0000_0000_0000;
array[61620] <= 16'b0000_0000_0000_0000;
array[61621] <= 16'b0000_0000_0000_0000;
array[61622] <= 16'b0000_0000_0000_0000;
array[61623] <= 16'b0000_0000_0000_0000;
array[61624] <= 16'b0000_0000_0000_0000;
array[61625] <= 16'b0000_0000_0000_0000;
array[61626] <= 16'b0000_0000_0000_0000;
array[61627] <= 16'b0000_0000_0000_0000;
array[61628] <= 16'b0000_0000_0000_0000;
array[61629] <= 16'b0000_0000_0000_0000;
array[61630] <= 16'b0000_0000_0000_0000;
array[61631] <= 16'b0000_0000_0000_0000;
array[61632] <= 16'b0000_0000_0000_0000;
array[61633] <= 16'b0000_0000_0000_0000;
array[61634] <= 16'b0000_0000_0000_0000;
array[61635] <= 16'b0000_0000_0000_0000;
array[61636] <= 16'b0000_0000_0000_0000;
array[61637] <= 16'b0000_0000_0000_0000;
array[61638] <= 16'b0000_0000_0000_0000;
array[61639] <= 16'b0000_0000_0000_0000;
array[61640] <= 16'b0000_0000_0000_0000;
array[61641] <= 16'b0000_0000_0000_0000;
array[61642] <= 16'b0000_0000_0000_0000;
array[61643] <= 16'b0000_0000_0000_0000;
array[61644] <= 16'b0000_0000_0000_0000;
array[61645] <= 16'b0000_0000_0000_0000;
array[61646] <= 16'b0000_0000_0000_0000;
array[61647] <= 16'b0000_0000_0000_0000;
array[61648] <= 16'b0000_0000_0000_0000;
array[61649] <= 16'b0000_0000_0000_0000;
array[61650] <= 16'b0000_0000_0000_0000;
array[61651] <= 16'b0000_0000_0000_0000;
array[61652] <= 16'b0000_0000_0000_0000;
array[61653] <= 16'b0000_0000_0000_0000;
array[61654] <= 16'b0000_0000_0000_0000;
array[61655] <= 16'b0000_0000_0000_0000;
array[61656] <= 16'b0000_0000_0000_0000;
array[61657] <= 16'b0000_0000_0000_0000;
array[61658] <= 16'b0000_0000_0000_0000;
array[61659] <= 16'b0000_0000_0000_0000;
array[61660] <= 16'b0000_0000_0000_0000;
array[61661] <= 16'b0000_0000_0000_0000;
array[61662] <= 16'b0000_0000_0000_0000;
array[61663] <= 16'b0000_0000_0000_0000;
array[61664] <= 16'b0000_0000_0000_0000;
array[61665] <= 16'b0000_0000_0000_0000;
array[61666] <= 16'b0000_0000_0000_0000;
array[61667] <= 16'b0000_0000_0000_0000;
array[61668] <= 16'b0000_0000_0000_0000;
array[61669] <= 16'b0000_0000_0000_0000;
array[61670] <= 16'b0000_0000_0000_0000;
array[61671] <= 16'b0000_0000_0000_0000;
array[61672] <= 16'b0000_0000_0000_0000;
array[61673] <= 16'b0000_0000_0000_0000;
array[61674] <= 16'b0000_0000_0000_0000;
array[61675] <= 16'b0000_0000_0000_0000;
array[61676] <= 16'b0000_0000_0000_0000;
array[61677] <= 16'b0000_0000_0000_0000;
array[61678] <= 16'b0000_0000_0000_0000;
array[61679] <= 16'b0000_0000_0000_0000;
array[61680] <= 16'b0000_0000_0000_0000;
array[61681] <= 16'b0000_0000_0000_0000;
array[61682] <= 16'b0000_0000_0000_0000;
array[61683] <= 16'b0000_0000_0000_0000;
array[61684] <= 16'b0000_0000_0000_0000;
array[61685] <= 16'b0000_0000_0000_0000;
array[61686] <= 16'b0000_0000_0000_0000;
array[61687] <= 16'b0000_0000_0000_0000;
array[61688] <= 16'b0000_0000_0000_0000;
array[61689] <= 16'b0000_0000_0000_0000;
array[61690] <= 16'b0000_0000_0000_0000;
array[61691] <= 16'b0000_0000_0000_0000;
array[61692] <= 16'b0000_0000_0000_0000;
array[61693] <= 16'b0000_0000_0000_0000;
array[61694] <= 16'b0000_0000_0000_0000;
array[61695] <= 16'b0000_0000_0000_0000;
array[61696] <= 16'b0000_0000_0000_0000;
array[61697] <= 16'b0000_0000_0000_0000;
array[61698] <= 16'b0000_0000_0000_0000;
array[61699] <= 16'b0000_0000_0000_0000;
array[61700] <= 16'b0000_0000_0000_0000;
array[61701] <= 16'b0000_0000_0000_0000;
array[61702] <= 16'b0000_0000_0000_0000;
array[61703] <= 16'b0000_0000_0000_0000;
array[61704] <= 16'b0000_0000_0000_0000;
array[61705] <= 16'b0000_0000_0000_0000;
array[61706] <= 16'b0000_0000_0000_0000;
array[61707] <= 16'b0000_0000_0000_0000;
array[61708] <= 16'b0000_0000_0000_0000;
array[61709] <= 16'b0000_0000_0000_0000;
array[61710] <= 16'b0000_0000_0000_0000;
array[61711] <= 16'b0000_0000_0000_0000;
array[61712] <= 16'b0000_0000_0000_0000;
array[61713] <= 16'b0000_0000_0000_0000;
array[61714] <= 16'b0000_0000_0000_0000;
array[61715] <= 16'b0000_0000_0000_0000;
array[61716] <= 16'b0000_0000_0000_0000;
array[61717] <= 16'b0000_0000_0000_0000;
array[61718] <= 16'b0000_0000_0000_0000;
array[61719] <= 16'b0000_0000_0000_0000;
array[61720] <= 16'b0000_0000_0000_0000;
array[61721] <= 16'b0000_0000_0000_0000;
array[61722] <= 16'b0000_0000_0000_0000;
array[61723] <= 16'b0000_0000_0000_0000;
array[61724] <= 16'b0000_0000_0000_0000;
array[61725] <= 16'b0000_0000_0000_0000;
array[61726] <= 16'b0000_0000_0000_0000;
array[61727] <= 16'b0000_0000_0000_0000;
array[61728] <= 16'b0000_0000_0000_0000;
array[61729] <= 16'b0000_0000_0000_0000;
array[61730] <= 16'b0000_0000_0000_0000;
array[61731] <= 16'b0000_0000_0000_0000;
array[61732] <= 16'b0000_0000_0000_0000;
array[61733] <= 16'b0000_0000_0000_0000;
array[61734] <= 16'b0000_0000_0000_0000;
array[61735] <= 16'b0000_0000_0000_0000;
array[61736] <= 16'b0000_0000_0000_0000;
array[61737] <= 16'b0000_0000_0000_0000;
array[61738] <= 16'b0000_0000_0000_0000;
array[61739] <= 16'b0000_0000_0000_0000;
array[61740] <= 16'b0000_0000_0000_0000;
array[61741] <= 16'b0000_0000_0000_0000;
array[61742] <= 16'b0000_0000_0000_0000;
array[61743] <= 16'b0000_0000_0000_0000;
array[61744] <= 16'b0000_0000_0000_0000;
array[61745] <= 16'b0000_0000_0000_0000;
array[61746] <= 16'b0000_0000_0000_0000;
array[61747] <= 16'b0000_0000_0000_0000;
array[61748] <= 16'b0000_0000_0000_0000;
array[61749] <= 16'b0000_0000_0000_0000;
array[61750] <= 16'b0000_0000_0000_0000;
array[61751] <= 16'b0000_0000_0000_0000;
array[61752] <= 16'b0000_0000_0000_0000;
array[61753] <= 16'b0000_0000_0000_0000;
array[61754] <= 16'b0000_0000_0000_0000;
array[61755] <= 16'b0000_0000_0000_0000;
array[61756] <= 16'b0000_0000_0000_0000;
array[61757] <= 16'b0000_0000_0000_0000;
array[61758] <= 16'b0000_0000_0000_0000;
array[61759] <= 16'b0000_0000_0000_0000;
array[61760] <= 16'b0000_0000_0000_0000;
array[61761] <= 16'b0000_0000_0000_0000;
array[61762] <= 16'b0000_0000_0000_0000;
array[61763] <= 16'b0000_0000_0000_0000;
array[61764] <= 16'b0000_0000_0000_0000;
array[61765] <= 16'b0000_0000_0000_0000;
array[61766] <= 16'b0000_0000_0000_0000;
array[61767] <= 16'b0000_0000_0000_0000;
array[61768] <= 16'b0000_0000_0000_0000;
array[61769] <= 16'b0000_0000_0000_0000;
array[61770] <= 16'b0000_0000_0000_0000;
array[61771] <= 16'b0000_0000_0000_0000;
array[61772] <= 16'b0000_0000_0000_0000;
array[61773] <= 16'b0000_0000_0000_0000;
array[61774] <= 16'b0000_0000_0000_0000;
array[61775] <= 16'b0000_0000_0000_0000;
array[61776] <= 16'b0000_0000_0000_0000;
array[61777] <= 16'b0000_0000_0000_0000;
array[61778] <= 16'b0000_0000_0000_0000;
array[61779] <= 16'b0000_0000_0000_0000;
array[61780] <= 16'b0000_0000_0000_0000;
array[61781] <= 16'b0000_0000_0000_0000;
array[61782] <= 16'b0000_0000_0000_0000;
array[61783] <= 16'b0000_0000_0000_0000;
array[61784] <= 16'b0000_0000_0000_0000;
array[61785] <= 16'b0000_0000_0000_0000;
array[61786] <= 16'b0000_0000_0000_0000;
array[61787] <= 16'b0000_0000_0000_0000;
array[61788] <= 16'b0000_0000_0000_0000;
array[61789] <= 16'b0000_0000_0000_0000;
array[61790] <= 16'b0000_0000_0000_0000;
array[61791] <= 16'b0000_0000_0000_0000;
array[61792] <= 16'b0000_0000_0000_0000;
array[61793] <= 16'b0000_0000_0000_0000;
array[61794] <= 16'b0000_0000_0000_0000;
array[61795] <= 16'b0000_0000_0000_0000;
array[61796] <= 16'b0000_0000_0000_0000;
array[61797] <= 16'b0000_0000_0000_0000;
array[61798] <= 16'b0000_0000_0000_0000;
array[61799] <= 16'b0000_0000_0000_0000;
array[61800] <= 16'b0000_0000_0000_0000;
array[61801] <= 16'b0000_0000_0000_0000;
array[61802] <= 16'b0000_0000_0000_0000;
array[61803] <= 16'b0000_0000_0000_0000;
array[61804] <= 16'b0000_0000_0000_0000;
array[61805] <= 16'b0000_0000_0000_0000;
array[61806] <= 16'b0000_0000_0000_0000;
array[61807] <= 16'b0000_0000_0000_0000;
array[61808] <= 16'b0000_0000_0000_0000;
array[61809] <= 16'b0000_0000_0000_0000;
array[61810] <= 16'b0000_0000_0000_0000;
array[61811] <= 16'b0000_0000_0000_0000;
array[61812] <= 16'b0000_0000_0000_0000;
array[61813] <= 16'b0000_0000_0000_0000;
array[61814] <= 16'b0000_0000_0000_0000;
array[61815] <= 16'b0000_0000_0000_0000;
array[61816] <= 16'b0000_0000_0000_0000;
array[61817] <= 16'b0000_0000_0000_0000;
array[61818] <= 16'b0000_0000_0000_0000;
array[61819] <= 16'b0000_0000_0000_0000;
array[61820] <= 16'b0000_0000_0000_0000;
array[61821] <= 16'b0000_0000_0000_0000;
array[61822] <= 16'b0000_0000_0000_0000;
array[61823] <= 16'b0000_0000_0000_0000;
array[61824] <= 16'b0000_0000_0000_0000;
array[61825] <= 16'b0000_0000_0000_0000;
array[61826] <= 16'b0000_0000_0000_0000;
array[61827] <= 16'b0000_0000_0000_0000;
array[61828] <= 16'b0000_0000_0000_0000;
array[61829] <= 16'b0000_0000_0000_0000;
array[61830] <= 16'b0000_0000_0000_0000;
array[61831] <= 16'b0000_0000_0000_0000;
array[61832] <= 16'b0000_0000_0000_0000;
array[61833] <= 16'b0000_0000_0000_0000;
array[61834] <= 16'b0000_0000_0000_0000;
array[61835] <= 16'b0000_0000_0000_0000;
array[61836] <= 16'b0000_0000_0000_0000;
array[61837] <= 16'b0000_0000_0000_0000;
array[61838] <= 16'b0000_0000_0000_0000;
array[61839] <= 16'b0000_0000_0000_0000;
array[61840] <= 16'b0000_0000_0000_0000;
array[61841] <= 16'b0000_0000_0000_0000;
array[61842] <= 16'b0000_0000_0000_0000;
array[61843] <= 16'b0000_0000_0000_0000;
array[61844] <= 16'b0000_0000_0000_0000;
array[61845] <= 16'b0000_0000_0000_0000;
array[61846] <= 16'b0000_0000_0000_0000;
array[61847] <= 16'b0000_0000_0000_0000;
array[61848] <= 16'b0000_0000_0000_0000;
array[61849] <= 16'b0000_0000_0000_0000;
array[61850] <= 16'b0000_0000_0000_0000;
array[61851] <= 16'b0000_0000_0000_0000;
array[61852] <= 16'b0000_0000_0000_0000;
array[61853] <= 16'b0000_0000_0000_0000;
array[61854] <= 16'b0000_0000_0000_0000;
array[61855] <= 16'b0000_0000_0000_0000;
array[61856] <= 16'b0000_0000_0000_0000;
array[61857] <= 16'b0000_0000_0000_0000;
array[61858] <= 16'b0000_0000_0000_0000;
array[61859] <= 16'b0000_0000_0000_0000;
array[61860] <= 16'b0000_0000_0000_0000;
array[61861] <= 16'b0000_0000_0000_0000;
array[61862] <= 16'b0000_0000_0000_0000;
array[61863] <= 16'b0000_0000_0000_0000;
array[61864] <= 16'b0000_0000_0000_0000;
array[61865] <= 16'b0000_0000_0000_0000;
array[61866] <= 16'b0000_0000_0000_0000;
array[61867] <= 16'b0000_0000_0000_0000;
array[61868] <= 16'b0000_0000_0000_0000;
array[61869] <= 16'b0000_0000_0000_0000;
array[61870] <= 16'b0000_0000_0000_0000;
array[61871] <= 16'b0000_0000_0000_0000;
array[61872] <= 16'b0000_0000_0000_0000;
array[61873] <= 16'b0000_0000_0000_0000;
array[61874] <= 16'b0000_0000_0000_0000;
array[61875] <= 16'b0000_0000_0000_0000;
array[61876] <= 16'b0000_0000_0000_0000;
array[61877] <= 16'b0000_0000_0000_0000;
array[61878] <= 16'b0000_0000_0000_0000;
array[61879] <= 16'b0000_0000_0000_0000;
array[61880] <= 16'b0000_0000_0000_0000;
array[61881] <= 16'b0000_0000_0000_0000;
array[61882] <= 16'b0000_0000_0000_0000;
array[61883] <= 16'b0000_0000_0000_0000;
array[61884] <= 16'b0000_0000_0000_0000;
array[61885] <= 16'b0000_0000_0000_0000;
array[61886] <= 16'b0000_0000_0000_0000;
array[61887] <= 16'b0000_0000_0000_0000;
array[61888] <= 16'b0000_0000_0000_0000;
array[61889] <= 16'b0000_0000_0000_0000;
array[61890] <= 16'b0000_0000_0000_0000;
array[61891] <= 16'b0000_0000_0000_0000;
array[61892] <= 16'b0000_0000_0000_0000;
array[61893] <= 16'b0000_0000_0000_0000;
array[61894] <= 16'b0000_0000_0000_0000;
array[61895] <= 16'b0000_0000_0000_0000;
array[61896] <= 16'b0000_0000_0000_0000;
array[61897] <= 16'b0000_0000_0000_0000;
array[61898] <= 16'b0000_0000_0000_0000;
array[61899] <= 16'b0000_0000_0000_0000;
array[61900] <= 16'b0000_0000_0000_0000;
array[61901] <= 16'b0000_0000_0000_0000;
array[61902] <= 16'b0000_0000_0000_0000;
array[61903] <= 16'b0000_0000_0000_0000;
array[61904] <= 16'b0000_0000_0000_0000;
array[61905] <= 16'b0000_0000_0000_0000;
array[61906] <= 16'b0000_0000_0000_0000;
array[61907] <= 16'b0000_0000_0000_0000;
array[61908] <= 16'b0000_0000_0000_0000;
array[61909] <= 16'b0000_0000_0000_0000;
array[61910] <= 16'b0000_0000_0000_0000;
array[61911] <= 16'b0000_0000_0000_0000;
array[61912] <= 16'b0000_0000_0000_0000;
array[61913] <= 16'b0000_0000_0000_0000;
array[61914] <= 16'b0000_0000_0000_0000;
array[61915] <= 16'b0000_0000_0000_0000;
array[61916] <= 16'b0000_0000_0000_0000;
array[61917] <= 16'b0000_0000_0000_0000;
array[61918] <= 16'b0000_0000_0000_0000;
array[61919] <= 16'b0000_0000_0000_0000;
array[61920] <= 16'b0000_0000_0000_0000;
array[61921] <= 16'b0000_0000_0000_0000;
array[61922] <= 16'b0000_0000_0000_0000;
array[61923] <= 16'b0000_0000_0000_0000;
array[61924] <= 16'b0000_0000_0000_0000;
array[61925] <= 16'b0000_0000_0000_0000;
array[61926] <= 16'b0000_0000_0000_0000;
array[61927] <= 16'b0000_0000_0000_0000;
array[61928] <= 16'b0000_0000_0000_0000;
array[61929] <= 16'b0000_0000_0000_0000;
array[61930] <= 16'b0000_0000_0000_0000;
array[61931] <= 16'b0000_0000_0000_0000;
array[61932] <= 16'b0000_0000_0000_0000;
array[61933] <= 16'b0000_0000_0000_0000;
array[61934] <= 16'b0000_0000_0000_0000;
array[61935] <= 16'b0000_0000_0000_0000;
array[61936] <= 16'b0000_0000_0000_0000;
array[61937] <= 16'b0000_0000_0000_0000;
array[61938] <= 16'b0000_0000_0000_0000;
array[61939] <= 16'b0000_0000_0000_0000;
array[61940] <= 16'b0000_0000_0000_0000;
array[61941] <= 16'b0000_0000_0000_0000;
array[61942] <= 16'b0000_0000_0000_0000;
array[61943] <= 16'b0000_0000_0000_0000;
array[61944] <= 16'b0000_0000_0000_0000;
array[61945] <= 16'b0000_0000_0000_0000;
array[61946] <= 16'b0000_0000_0000_0000;
array[61947] <= 16'b0000_0000_0000_0000;
array[61948] <= 16'b0000_0000_0000_0000;
array[61949] <= 16'b0000_0000_0000_0000;
array[61950] <= 16'b0000_0000_0000_0000;
array[61951] <= 16'b0000_0000_0000_0000;
array[61952] <= 16'b0000_0000_0000_0000;
array[61953] <= 16'b0000_0000_0000_0000;
array[61954] <= 16'b0000_0000_0000_0000;
array[61955] <= 16'b0000_0000_0000_0000;
array[61956] <= 16'b0000_0000_0000_0000;
array[61957] <= 16'b0000_0000_0000_0000;
array[61958] <= 16'b0000_0000_0000_0000;
array[61959] <= 16'b0000_0000_0000_0000;
array[61960] <= 16'b0000_0000_0000_0000;
array[61961] <= 16'b0000_0000_0000_0000;
array[61962] <= 16'b0000_0000_0000_0000;
array[61963] <= 16'b0000_0000_0000_0000;
array[61964] <= 16'b0000_0000_0000_0000;
array[61965] <= 16'b0000_0000_0000_0000;
array[61966] <= 16'b0000_0000_0000_0000;
array[61967] <= 16'b0000_0000_0000_0000;
array[61968] <= 16'b0000_0000_0000_0000;
array[61969] <= 16'b0000_0000_0000_0000;
array[61970] <= 16'b0000_0000_0000_0000;
array[61971] <= 16'b0000_0000_0000_0000;
array[61972] <= 16'b0000_0000_0000_0000;
array[61973] <= 16'b0000_0000_0000_0000;
array[61974] <= 16'b0000_0000_0000_0000;
array[61975] <= 16'b0000_0000_0000_0000;
array[61976] <= 16'b0000_0000_0000_0000;
array[61977] <= 16'b0000_0000_0000_0000;
array[61978] <= 16'b0000_0000_0000_0000;
array[61979] <= 16'b0000_0000_0000_0000;
array[61980] <= 16'b0000_0000_0000_0000;
array[61981] <= 16'b0000_0000_0000_0000;
array[61982] <= 16'b0000_0000_0000_0000;
array[61983] <= 16'b0000_0000_0000_0000;
array[61984] <= 16'b0000_0000_0000_0000;
array[61985] <= 16'b0000_0000_0000_0000;
array[61986] <= 16'b0000_0000_0000_0000;
array[61987] <= 16'b0000_0000_0000_0000;
array[61988] <= 16'b0000_0000_0000_0000;
array[61989] <= 16'b0000_0000_0000_0000;
array[61990] <= 16'b0000_0000_0000_0000;
array[61991] <= 16'b0000_0000_0000_0000;
array[61992] <= 16'b0000_0000_0000_0000;
array[61993] <= 16'b0000_0000_0000_0000;
array[61994] <= 16'b0000_0000_0000_0000;
array[61995] <= 16'b0000_0000_0000_0000;
array[61996] <= 16'b0000_0000_0000_0000;
array[61997] <= 16'b0000_0000_0000_0000;
array[61998] <= 16'b0000_0000_0000_0000;
array[61999] <= 16'b0000_0000_0000_0000;
array[62000] <= 16'b0000_0000_0000_0000;
array[62001] <= 16'b0000_0000_0000_0000;
array[62002] <= 16'b0000_0000_0000_0000;
array[62003] <= 16'b0000_0000_0000_0000;
array[62004] <= 16'b0000_0000_0000_0000;
array[62005] <= 16'b0000_0000_0000_0000;
array[62006] <= 16'b0000_0000_0000_0000;
array[62007] <= 16'b0000_0000_0000_0000;
array[62008] <= 16'b0000_0000_0000_0000;
array[62009] <= 16'b0000_0000_0000_0000;
array[62010] <= 16'b0000_0000_0000_0000;
array[62011] <= 16'b0000_0000_0000_0000;
array[62012] <= 16'b0000_0000_0000_0000;
array[62013] <= 16'b0000_0000_0000_0000;
array[62014] <= 16'b0000_0000_0000_0000;
array[62015] <= 16'b0000_0000_0000_0000;
array[62016] <= 16'b0000_0000_0000_0000;
array[62017] <= 16'b0000_0000_0000_0000;
array[62018] <= 16'b0000_0000_0000_0000;
array[62019] <= 16'b0000_0000_0000_0000;
array[62020] <= 16'b0000_0000_0000_0000;
array[62021] <= 16'b0000_0000_0000_0000;
array[62022] <= 16'b0000_0000_0000_0000;
array[62023] <= 16'b0000_0000_0000_0000;
array[62024] <= 16'b0000_0000_0000_0000;
array[62025] <= 16'b0000_0000_0000_0000;
array[62026] <= 16'b0000_0000_0000_0000;
array[62027] <= 16'b0000_0000_0000_0000;
array[62028] <= 16'b0000_0000_0000_0000;
array[62029] <= 16'b0000_0000_0000_0000;
array[62030] <= 16'b0000_0000_0000_0000;
array[62031] <= 16'b0000_0000_0000_0000;
array[62032] <= 16'b0000_0000_0000_0000;
array[62033] <= 16'b0000_0000_0000_0000;
array[62034] <= 16'b0000_0000_0000_0000;
array[62035] <= 16'b0000_0000_0000_0000;
array[62036] <= 16'b0000_0000_0000_0000;
array[62037] <= 16'b0000_0000_0000_0000;
array[62038] <= 16'b0000_0000_0000_0000;
array[62039] <= 16'b0000_0000_0000_0000;
array[62040] <= 16'b0000_0000_0000_0000;
array[62041] <= 16'b0000_0000_0000_0000;
array[62042] <= 16'b0000_0000_0000_0000;
array[62043] <= 16'b0000_0000_0000_0000;
array[62044] <= 16'b0000_0000_0000_0000;
array[62045] <= 16'b0000_0000_0000_0000;
array[62046] <= 16'b0000_0000_0000_0000;
array[62047] <= 16'b0000_0000_0000_0000;
array[62048] <= 16'b0000_0000_0000_0000;
array[62049] <= 16'b0000_0000_0000_0000;
array[62050] <= 16'b0000_0000_0000_0000;
array[62051] <= 16'b0000_0000_0000_0000;
array[62052] <= 16'b0000_0000_0000_0000;
array[62053] <= 16'b0000_0000_0000_0000;
array[62054] <= 16'b0000_0000_0000_0000;
array[62055] <= 16'b0000_0000_0000_0000;
array[62056] <= 16'b0000_0000_0000_0000;
array[62057] <= 16'b0000_0000_0000_0000;
array[62058] <= 16'b0000_0000_0000_0000;
array[62059] <= 16'b0000_0000_0000_0000;
array[62060] <= 16'b0000_0000_0000_0000;
array[62061] <= 16'b0000_0000_0000_0000;
array[62062] <= 16'b0000_0000_0000_0000;
array[62063] <= 16'b0000_0000_0000_0000;
array[62064] <= 16'b0000_0000_0000_0000;
array[62065] <= 16'b0000_0000_0000_0000;
array[62066] <= 16'b0000_0000_0000_0000;
array[62067] <= 16'b0000_0000_0000_0000;
array[62068] <= 16'b0000_0000_0000_0000;
array[62069] <= 16'b0000_0000_0000_0000;
array[62070] <= 16'b0000_0000_0000_0000;
array[62071] <= 16'b0000_0000_0000_0000;
array[62072] <= 16'b0000_0000_0000_0000;
array[62073] <= 16'b0000_0000_0000_0000;
array[62074] <= 16'b0000_0000_0000_0000;
array[62075] <= 16'b0000_0000_0000_0000;
array[62076] <= 16'b0000_0000_0000_0000;
array[62077] <= 16'b0000_0000_0000_0000;
array[62078] <= 16'b0000_0000_0000_0000;
array[62079] <= 16'b0000_0000_0000_0000;
array[62080] <= 16'b0000_0000_0000_0000;
array[62081] <= 16'b0000_0000_0000_0000;
array[62082] <= 16'b0000_0000_0000_0000;
array[62083] <= 16'b0000_0000_0000_0000;
array[62084] <= 16'b0000_0000_0000_0000;
array[62085] <= 16'b0000_0000_0000_0000;
array[62086] <= 16'b0000_0000_0000_0000;
array[62087] <= 16'b0000_0000_0000_0000;
array[62088] <= 16'b0000_0000_0000_0000;
array[62089] <= 16'b0000_0000_0000_0000;
array[62090] <= 16'b0000_0000_0000_0000;
array[62091] <= 16'b0000_0000_0000_0000;
array[62092] <= 16'b0000_0000_0000_0000;
array[62093] <= 16'b0000_0000_0000_0000;
array[62094] <= 16'b0000_0000_0000_0000;
array[62095] <= 16'b0000_0000_0000_0000;
array[62096] <= 16'b0000_0000_0000_0000;
array[62097] <= 16'b0000_0000_0000_0000;
array[62098] <= 16'b0000_0000_0000_0000;
array[62099] <= 16'b0000_0000_0000_0000;
array[62100] <= 16'b0000_0000_0000_0000;
array[62101] <= 16'b0000_0000_0000_0000;
array[62102] <= 16'b0000_0000_0000_0000;
array[62103] <= 16'b0000_0000_0000_0000;
array[62104] <= 16'b0000_0000_0000_0000;
array[62105] <= 16'b0000_0000_0000_0000;
array[62106] <= 16'b0000_0000_0000_0000;
array[62107] <= 16'b0000_0000_0000_0000;
array[62108] <= 16'b0000_0000_0000_0000;
array[62109] <= 16'b0000_0000_0000_0000;
array[62110] <= 16'b0000_0000_0000_0000;
array[62111] <= 16'b0000_0000_0000_0000;
array[62112] <= 16'b0000_0000_0000_0000;
array[62113] <= 16'b0000_0000_0000_0000;
array[62114] <= 16'b0000_0000_0000_0000;
array[62115] <= 16'b0000_0000_0000_0000;
array[62116] <= 16'b0000_0000_0000_0000;
array[62117] <= 16'b0000_0000_0000_0000;
array[62118] <= 16'b0000_0000_0000_0000;
array[62119] <= 16'b0000_0000_0000_0000;
array[62120] <= 16'b0000_0000_0000_0000;
array[62121] <= 16'b0000_0000_0000_0000;
array[62122] <= 16'b0000_0000_0000_0000;
array[62123] <= 16'b0000_0000_0000_0000;
array[62124] <= 16'b0000_0000_0000_0000;
array[62125] <= 16'b0000_0000_0000_0000;
array[62126] <= 16'b0000_0000_0000_0000;
array[62127] <= 16'b0000_0000_0000_0000;
array[62128] <= 16'b0000_0000_0000_0000;
array[62129] <= 16'b0000_0000_0000_0000;
array[62130] <= 16'b0000_0000_0000_0000;
array[62131] <= 16'b0000_0000_0000_0000;
array[62132] <= 16'b0000_0000_0000_0000;
array[62133] <= 16'b0000_0000_0000_0000;
array[62134] <= 16'b0000_0000_0000_0000;
array[62135] <= 16'b0000_0000_0000_0000;
array[62136] <= 16'b0000_0000_0000_0000;
array[62137] <= 16'b0000_0000_0000_0000;
array[62138] <= 16'b0000_0000_0000_0000;
array[62139] <= 16'b0000_0000_0000_0000;
array[62140] <= 16'b0000_0000_0000_0000;
array[62141] <= 16'b0000_0000_0000_0000;
array[62142] <= 16'b0000_0000_0000_0000;
array[62143] <= 16'b0000_0000_0000_0000;
array[62144] <= 16'b0000_0000_0000_0000;
array[62145] <= 16'b0000_0000_0000_0000;
array[62146] <= 16'b0000_0000_0000_0000;
array[62147] <= 16'b0000_0000_0000_0000;
array[62148] <= 16'b0000_0000_0000_0000;
array[62149] <= 16'b0000_0000_0000_0000;
array[62150] <= 16'b0000_0000_0000_0000;
array[62151] <= 16'b0000_0000_0000_0000;
array[62152] <= 16'b0000_0000_0000_0000;
array[62153] <= 16'b0000_0000_0000_0000;
array[62154] <= 16'b0000_0000_0000_0000;
array[62155] <= 16'b0000_0000_0000_0000;
array[62156] <= 16'b0000_0000_0000_0000;
array[62157] <= 16'b0000_0000_0000_0000;
array[62158] <= 16'b0000_0000_0000_0000;
array[62159] <= 16'b0000_0000_0000_0000;
array[62160] <= 16'b0000_0000_0000_0000;
array[62161] <= 16'b0000_0000_0000_0000;
array[62162] <= 16'b0000_0000_0000_0000;
array[62163] <= 16'b0000_0000_0000_0000;
array[62164] <= 16'b0000_0000_0000_0000;
array[62165] <= 16'b0000_0000_0000_0000;
array[62166] <= 16'b0000_0000_0000_0000;
array[62167] <= 16'b0000_0000_0000_0000;
array[62168] <= 16'b0000_0000_0000_0000;
array[62169] <= 16'b0000_0000_0000_0000;
array[62170] <= 16'b0000_0000_0000_0000;
array[62171] <= 16'b0000_0000_0000_0000;
array[62172] <= 16'b0000_0000_0000_0000;
array[62173] <= 16'b0000_0000_0000_0000;
array[62174] <= 16'b0000_0000_0000_0000;
array[62175] <= 16'b0000_0000_0000_0000;
array[62176] <= 16'b0000_0000_0000_0000;
array[62177] <= 16'b0000_0000_0000_0000;
array[62178] <= 16'b0000_0000_0000_0000;
array[62179] <= 16'b0000_0000_0000_0000;
array[62180] <= 16'b0000_0000_0000_0000;
array[62181] <= 16'b0000_0000_0000_0000;
array[62182] <= 16'b0000_0000_0000_0000;
array[62183] <= 16'b0000_0000_0000_0000;
array[62184] <= 16'b0000_0000_0000_0000;
array[62185] <= 16'b0000_0000_0000_0000;
array[62186] <= 16'b0000_0000_0000_0000;
array[62187] <= 16'b0000_0000_0000_0000;
array[62188] <= 16'b0000_0000_0000_0000;
array[62189] <= 16'b0000_0000_0000_0000;
array[62190] <= 16'b0000_0000_0000_0000;
array[62191] <= 16'b0000_0000_0000_0000;
array[62192] <= 16'b0000_0000_0000_0000;
array[62193] <= 16'b0000_0000_0000_0000;
array[62194] <= 16'b0000_0000_0000_0000;
array[62195] <= 16'b0000_0000_0000_0000;
array[62196] <= 16'b0000_0000_0000_0000;
array[62197] <= 16'b0000_0000_0000_0000;
array[62198] <= 16'b0000_0000_0000_0000;
array[62199] <= 16'b0000_0000_0000_0000;
array[62200] <= 16'b0000_0000_0000_0000;
array[62201] <= 16'b0000_0000_0000_0000;
array[62202] <= 16'b0000_0000_0000_0000;
array[62203] <= 16'b0000_0000_0000_0000;
array[62204] <= 16'b0000_0000_0000_0000;
array[62205] <= 16'b0000_0000_0000_0000;
array[62206] <= 16'b0000_0000_0000_0000;
array[62207] <= 16'b0000_0000_0000_0000;
array[62208] <= 16'b0000_0000_0000_0000;
array[62209] <= 16'b0000_0000_0000_0000;
array[62210] <= 16'b0000_0000_0000_0000;
array[62211] <= 16'b0000_0000_0000_0000;
array[62212] <= 16'b0000_0000_0000_0000;
array[62213] <= 16'b0000_0000_0000_0000;
array[62214] <= 16'b0000_0000_0000_0000;
array[62215] <= 16'b0000_0000_0000_0000;
array[62216] <= 16'b0000_0000_0000_0000;
array[62217] <= 16'b0000_0000_0000_0000;
array[62218] <= 16'b0000_0000_0000_0000;
array[62219] <= 16'b0000_0000_0000_0000;
array[62220] <= 16'b0000_0000_0000_0000;
array[62221] <= 16'b0000_0000_0000_0000;
array[62222] <= 16'b0000_0000_0000_0000;
array[62223] <= 16'b0000_0000_0000_0000;
array[62224] <= 16'b0000_0000_0000_0000;
array[62225] <= 16'b0000_0000_0000_0000;
array[62226] <= 16'b0000_0000_0000_0000;
array[62227] <= 16'b0000_0000_0000_0000;
array[62228] <= 16'b0000_0000_0000_0000;
array[62229] <= 16'b0000_0000_0000_0000;
array[62230] <= 16'b0000_0000_0000_0000;
array[62231] <= 16'b0000_0000_0000_0000;
array[62232] <= 16'b0000_0000_0000_0000;
array[62233] <= 16'b0000_0000_0000_0000;
array[62234] <= 16'b0000_0000_0000_0000;
array[62235] <= 16'b0000_0000_0000_0000;
array[62236] <= 16'b0000_0000_0000_0000;
array[62237] <= 16'b0000_0000_0000_0000;
array[62238] <= 16'b0000_0000_0000_0000;
array[62239] <= 16'b0000_0000_0000_0000;
array[62240] <= 16'b0000_0000_0000_0000;
array[62241] <= 16'b0000_0000_0000_0000;
array[62242] <= 16'b0000_0000_0000_0000;
array[62243] <= 16'b0000_0000_0000_0000;
array[62244] <= 16'b0000_0000_0000_0000;
array[62245] <= 16'b0000_0000_0000_0000;
array[62246] <= 16'b0000_0000_0000_0000;
array[62247] <= 16'b0000_0000_0000_0000;
array[62248] <= 16'b0000_0000_0000_0000;
array[62249] <= 16'b0000_0000_0000_0000;
array[62250] <= 16'b0000_0000_0000_0000;
array[62251] <= 16'b0000_0000_0000_0000;
array[62252] <= 16'b0000_0000_0000_0000;
array[62253] <= 16'b0000_0000_0000_0000;
array[62254] <= 16'b0000_0000_0000_0000;
array[62255] <= 16'b0000_0000_0000_0000;
array[62256] <= 16'b0000_0000_0000_0000;
array[62257] <= 16'b0000_0000_0000_0000;
array[62258] <= 16'b0000_0000_0000_0000;
array[62259] <= 16'b0000_0000_0000_0000;
array[62260] <= 16'b0000_0000_0000_0000;
array[62261] <= 16'b0000_0000_0000_0000;
array[62262] <= 16'b0000_0000_0000_0000;
array[62263] <= 16'b0000_0000_0000_0000;
array[62264] <= 16'b0000_0000_0000_0000;
array[62265] <= 16'b0000_0000_0000_0000;
array[62266] <= 16'b0000_0000_0000_0000;
array[62267] <= 16'b0000_0000_0000_0000;
array[62268] <= 16'b0000_0000_0000_0000;
array[62269] <= 16'b0000_0000_0000_0000;
array[62270] <= 16'b0000_0000_0000_0000;
array[62271] <= 16'b0000_0000_0000_0000;
array[62272] <= 16'b0000_0000_0000_0000;
array[62273] <= 16'b0000_0000_0000_0000;
array[62274] <= 16'b0000_0000_0000_0000;
array[62275] <= 16'b0000_0000_0000_0000;
array[62276] <= 16'b0000_0000_0000_0000;
array[62277] <= 16'b0000_0000_0000_0000;
array[62278] <= 16'b0000_0000_0000_0000;
array[62279] <= 16'b0000_0000_0000_0000;
array[62280] <= 16'b0000_0000_0000_0000;
array[62281] <= 16'b0000_0000_0000_0000;
array[62282] <= 16'b0000_0000_0000_0000;
array[62283] <= 16'b0000_0000_0000_0000;
array[62284] <= 16'b0000_0000_0000_0000;
array[62285] <= 16'b0000_0000_0000_0000;
array[62286] <= 16'b0000_0000_0000_0000;
array[62287] <= 16'b0000_0000_0000_0000;
array[62288] <= 16'b0000_0000_0000_0000;
array[62289] <= 16'b0000_0000_0000_0000;
array[62290] <= 16'b0000_0000_0000_0000;
array[62291] <= 16'b0000_0000_0000_0000;
array[62292] <= 16'b0000_0000_0000_0000;
array[62293] <= 16'b0000_0000_0000_0000;
array[62294] <= 16'b0000_0000_0000_0000;
array[62295] <= 16'b0000_0000_0000_0000;
array[62296] <= 16'b0000_0000_0000_0000;
array[62297] <= 16'b0000_0000_0000_0000;
array[62298] <= 16'b0000_0000_0000_0000;
array[62299] <= 16'b0000_0000_0000_0000;
array[62300] <= 16'b0000_0000_0000_0000;
array[62301] <= 16'b0000_0000_0000_0000;
array[62302] <= 16'b0000_0000_0000_0000;
array[62303] <= 16'b0000_0000_0000_0000;
array[62304] <= 16'b0000_0000_0000_0000;
array[62305] <= 16'b0000_0000_0000_0000;
array[62306] <= 16'b0000_0000_0000_0000;
array[62307] <= 16'b0000_0000_0000_0000;
array[62308] <= 16'b0000_0000_0000_0000;
array[62309] <= 16'b0000_0000_0000_0000;
array[62310] <= 16'b0000_0000_0000_0000;
array[62311] <= 16'b0000_0000_0000_0000;
array[62312] <= 16'b0000_0000_0000_0000;
array[62313] <= 16'b0000_0000_0000_0000;
array[62314] <= 16'b0000_0000_0000_0000;
array[62315] <= 16'b0000_0000_0000_0000;
array[62316] <= 16'b0000_0000_0000_0000;
array[62317] <= 16'b0000_0000_0000_0000;
array[62318] <= 16'b0000_0000_0000_0000;
array[62319] <= 16'b0000_0000_0000_0000;
array[62320] <= 16'b0000_0000_0000_0000;
array[62321] <= 16'b0000_0000_0000_0000;
array[62322] <= 16'b0000_0000_0000_0000;
array[62323] <= 16'b0000_0000_0000_0000;
array[62324] <= 16'b0000_0000_0000_0000;
array[62325] <= 16'b0000_0000_0000_0000;
array[62326] <= 16'b0000_0000_0000_0000;
array[62327] <= 16'b0000_0000_0000_0000;
array[62328] <= 16'b0000_0000_0000_0000;
array[62329] <= 16'b0000_0000_0000_0000;
array[62330] <= 16'b0000_0000_0000_0000;
array[62331] <= 16'b0000_0000_0000_0000;
array[62332] <= 16'b0000_0000_0000_0000;
array[62333] <= 16'b0000_0000_0000_0000;
array[62334] <= 16'b0000_0000_0000_0000;
array[62335] <= 16'b0000_0000_0000_0000;
array[62336] <= 16'b0000_0000_0000_0000;
array[62337] <= 16'b0000_0000_0000_0000;
array[62338] <= 16'b0000_0000_0000_0000;
array[62339] <= 16'b0000_0000_0000_0000;
array[62340] <= 16'b0000_0000_0000_0000;
array[62341] <= 16'b0000_0000_0000_0000;
array[62342] <= 16'b0000_0000_0000_0000;
array[62343] <= 16'b0000_0000_0000_0000;
array[62344] <= 16'b0000_0000_0000_0000;
array[62345] <= 16'b0000_0000_0000_0000;
array[62346] <= 16'b0000_0000_0000_0000;
array[62347] <= 16'b0000_0000_0000_0000;
array[62348] <= 16'b0000_0000_0000_0000;
array[62349] <= 16'b0000_0000_0000_0000;
array[62350] <= 16'b0000_0000_0000_0000;
array[62351] <= 16'b0000_0000_0000_0000;
array[62352] <= 16'b0000_0000_0000_0000;
array[62353] <= 16'b0000_0000_0000_0000;
array[62354] <= 16'b0000_0000_0000_0000;
array[62355] <= 16'b0000_0000_0000_0000;
array[62356] <= 16'b0000_0000_0000_0000;
array[62357] <= 16'b0000_0000_0000_0000;
array[62358] <= 16'b0000_0000_0000_0000;
array[62359] <= 16'b0000_0000_0000_0000;
array[62360] <= 16'b0000_0000_0000_0000;
array[62361] <= 16'b0000_0000_0000_0000;
array[62362] <= 16'b0000_0000_0000_0000;
array[62363] <= 16'b0000_0000_0000_0000;
array[62364] <= 16'b0000_0000_0000_0000;
array[62365] <= 16'b0000_0000_0000_0000;
array[62366] <= 16'b0000_0000_0000_0000;
array[62367] <= 16'b0000_0000_0000_0000;
array[62368] <= 16'b0000_0000_0000_0000;
array[62369] <= 16'b0000_0000_0000_0000;
array[62370] <= 16'b0000_0000_0000_0000;
array[62371] <= 16'b0000_0000_0000_0000;
array[62372] <= 16'b0000_0000_0000_0000;
array[62373] <= 16'b0000_0000_0000_0000;
array[62374] <= 16'b0000_0000_0000_0000;
array[62375] <= 16'b0000_0000_0000_0000;
array[62376] <= 16'b0000_0000_0000_0000;
array[62377] <= 16'b0000_0000_0000_0000;
array[62378] <= 16'b0000_0000_0000_0000;
array[62379] <= 16'b0000_0000_0000_0000;
array[62380] <= 16'b0000_0000_0000_0000;
array[62381] <= 16'b0000_0000_0000_0000;
array[62382] <= 16'b0000_0000_0000_0000;
array[62383] <= 16'b0000_0000_0000_0000;
array[62384] <= 16'b0000_0000_0000_0000;
array[62385] <= 16'b0000_0000_0000_0000;
array[62386] <= 16'b0000_0000_0000_0000;
array[62387] <= 16'b0000_0000_0000_0000;
array[62388] <= 16'b0000_0000_0000_0000;
array[62389] <= 16'b0000_0000_0000_0000;
array[62390] <= 16'b0000_0000_0000_0000;
array[62391] <= 16'b0000_0000_0000_0000;
array[62392] <= 16'b0000_0000_0000_0000;
array[62393] <= 16'b0000_0000_0000_0000;
array[62394] <= 16'b0000_0000_0000_0000;
array[62395] <= 16'b0000_0000_0000_0000;
array[62396] <= 16'b0000_0000_0000_0000;
array[62397] <= 16'b0000_0000_0000_0000;
array[62398] <= 16'b0000_0000_0000_0000;
array[62399] <= 16'b0000_0000_0000_0000;
array[62400] <= 16'b0000_0000_0000_0000;
array[62401] <= 16'b0000_0000_0000_0000;
array[62402] <= 16'b0000_0000_0000_0000;
array[62403] <= 16'b0000_0000_0000_0000;
array[62404] <= 16'b0000_0000_0000_0000;
array[62405] <= 16'b0000_0000_0000_0000;
array[62406] <= 16'b0000_0000_0000_0000;
array[62407] <= 16'b0000_0000_0000_0000;
array[62408] <= 16'b0000_0000_0000_0000;
array[62409] <= 16'b0000_0000_0000_0000;
array[62410] <= 16'b0000_0000_0000_0000;
array[62411] <= 16'b0000_0000_0000_0000;
array[62412] <= 16'b0000_0000_0000_0000;
array[62413] <= 16'b0000_0000_0000_0000;
array[62414] <= 16'b0000_0000_0000_0000;
array[62415] <= 16'b0000_0000_0000_0000;
array[62416] <= 16'b0000_0000_0000_0000;
array[62417] <= 16'b0000_0000_0000_0000;
array[62418] <= 16'b0000_0000_0000_0000;
array[62419] <= 16'b0000_0000_0000_0000;
array[62420] <= 16'b0000_0000_0000_0000;
array[62421] <= 16'b0000_0000_0000_0000;
array[62422] <= 16'b0000_0000_0000_0000;
array[62423] <= 16'b0000_0000_0000_0000;
array[62424] <= 16'b0000_0000_0000_0000;
array[62425] <= 16'b0000_0000_0000_0000;
array[62426] <= 16'b0000_0000_0000_0000;
array[62427] <= 16'b0000_0000_0000_0000;
array[62428] <= 16'b0000_0000_0000_0000;
array[62429] <= 16'b0000_0000_0000_0000;
array[62430] <= 16'b0000_0000_0000_0000;
array[62431] <= 16'b0000_0000_0000_0000;
array[62432] <= 16'b0000_0000_0000_0000;
array[62433] <= 16'b0000_0000_0000_0000;
array[62434] <= 16'b0000_0000_0000_0000;
array[62435] <= 16'b0000_0000_0000_0000;
array[62436] <= 16'b0000_0000_0000_0000;
array[62437] <= 16'b0000_0000_0000_0000;
array[62438] <= 16'b0000_0000_0000_0000;
array[62439] <= 16'b0000_0000_0000_0000;
array[62440] <= 16'b0000_0000_0000_0000;
array[62441] <= 16'b0000_0000_0000_0000;
array[62442] <= 16'b0000_0000_0000_0000;
array[62443] <= 16'b0000_0000_0000_0000;
array[62444] <= 16'b0000_0000_0000_0000;
array[62445] <= 16'b0000_0000_0000_0000;
array[62446] <= 16'b0000_0000_0000_0000;
array[62447] <= 16'b0000_0000_0000_0000;
array[62448] <= 16'b0000_0000_0000_0000;
array[62449] <= 16'b0000_0000_0000_0000;
array[62450] <= 16'b0000_0000_0000_0000;
array[62451] <= 16'b0000_0000_0000_0000;
array[62452] <= 16'b0000_0000_0000_0000;
array[62453] <= 16'b0000_0000_0000_0000;
array[62454] <= 16'b0000_0000_0000_0000;
array[62455] <= 16'b0000_0000_0000_0000;
array[62456] <= 16'b0000_0000_0000_0000;
array[62457] <= 16'b0000_0000_0000_0000;
array[62458] <= 16'b0000_0000_0000_0000;
array[62459] <= 16'b0000_0000_0000_0000;
array[62460] <= 16'b0000_0000_0000_0000;
array[62461] <= 16'b0000_0000_0000_0000;
array[62462] <= 16'b0000_0000_0000_0000;
array[62463] <= 16'b0000_0000_0000_0000;
array[62464] <= 16'b0000_0000_0000_0000;
array[62465] <= 16'b0000_0000_0000_0000;
array[62466] <= 16'b0000_0000_0000_0000;
array[62467] <= 16'b0000_0000_0000_0000;
array[62468] <= 16'b0000_0000_0000_0000;
array[62469] <= 16'b0000_0000_0000_0000;
array[62470] <= 16'b0000_0000_0000_0000;
array[62471] <= 16'b0000_0000_0000_0000;
array[62472] <= 16'b0000_0000_0000_0000;
array[62473] <= 16'b0000_0000_0000_0000;
array[62474] <= 16'b0000_0000_0000_0000;
array[62475] <= 16'b0000_0000_0000_0000;
array[62476] <= 16'b0000_0000_0000_0000;
array[62477] <= 16'b0000_0000_0000_0000;
array[62478] <= 16'b0000_0000_0000_0000;
array[62479] <= 16'b0000_0000_0000_0000;
array[62480] <= 16'b0000_0000_0000_0000;
array[62481] <= 16'b0000_0000_0000_0000;
array[62482] <= 16'b0000_0000_0000_0000;
array[62483] <= 16'b0000_0000_0000_0000;
array[62484] <= 16'b0000_0000_0000_0000;
array[62485] <= 16'b0000_0000_0000_0000;
array[62486] <= 16'b0000_0000_0000_0000;
array[62487] <= 16'b0000_0000_0000_0000;
array[62488] <= 16'b0000_0000_0000_0000;
array[62489] <= 16'b0000_0000_0000_0000;
array[62490] <= 16'b0000_0000_0000_0000;
array[62491] <= 16'b0000_0000_0000_0000;
array[62492] <= 16'b0000_0000_0000_0000;
array[62493] <= 16'b0000_0000_0000_0000;
array[62494] <= 16'b0000_0000_0000_0000;
array[62495] <= 16'b0000_0000_0000_0000;
array[62496] <= 16'b0000_0000_0000_0000;
array[62497] <= 16'b0000_0000_0000_0000;
array[62498] <= 16'b0000_0000_0000_0000;
array[62499] <= 16'b0000_0000_0000_0000;
array[62500] <= 16'b0000_0000_0000_0000;
array[62501] <= 16'b0000_0000_0000_0000;
array[62502] <= 16'b0000_0000_0000_0000;
array[62503] <= 16'b0000_0000_0000_0000;
array[62504] <= 16'b0000_0000_0000_0000;
array[62505] <= 16'b0000_0000_0000_0000;
array[62506] <= 16'b0000_0000_0000_0000;
array[62507] <= 16'b0000_0000_0000_0000;
array[62508] <= 16'b0000_0000_0000_0000;
array[62509] <= 16'b0000_0000_0000_0000;
array[62510] <= 16'b0000_0000_0000_0000;
array[62511] <= 16'b0000_0000_0000_0000;
array[62512] <= 16'b0000_0000_0000_0000;
array[62513] <= 16'b0000_0000_0000_0000;
array[62514] <= 16'b0000_0000_0000_0000;
array[62515] <= 16'b0000_0000_0000_0000;
array[62516] <= 16'b0000_0000_0000_0000;
array[62517] <= 16'b0000_0000_0000_0000;
array[62518] <= 16'b0000_0000_0000_0000;
array[62519] <= 16'b0000_0000_0000_0000;
array[62520] <= 16'b0000_0000_0000_0000;
array[62521] <= 16'b0000_0000_0000_0000;
array[62522] <= 16'b0000_0000_0000_0000;
array[62523] <= 16'b0000_0000_0000_0000;
array[62524] <= 16'b0000_0000_0000_0000;
array[62525] <= 16'b0000_0000_0000_0000;
array[62526] <= 16'b0000_0000_0000_0000;
array[62527] <= 16'b0000_0000_0000_0000;
array[62528] <= 16'b0000_0000_0000_0000;
array[62529] <= 16'b0000_0000_0000_0000;
array[62530] <= 16'b0000_0000_0000_0000;
array[62531] <= 16'b0000_0000_0000_0000;
array[62532] <= 16'b0000_0000_0000_0000;
array[62533] <= 16'b0000_0000_0000_0000;
array[62534] <= 16'b0000_0000_0000_0000;
array[62535] <= 16'b0000_0000_0000_0000;
array[62536] <= 16'b0000_0000_0000_0000;
array[62537] <= 16'b0000_0000_0000_0000;
array[62538] <= 16'b0000_0000_0000_0000;
array[62539] <= 16'b0000_0000_0000_0000;
array[62540] <= 16'b0000_0000_0000_0000;
array[62541] <= 16'b0000_0000_0000_0000;
array[62542] <= 16'b0000_0000_0000_0000;
array[62543] <= 16'b0000_0000_0000_0000;
array[62544] <= 16'b0000_0000_0000_0000;
array[62545] <= 16'b0000_0000_0000_0000;
array[62546] <= 16'b0000_0000_0000_0000;
array[62547] <= 16'b0000_0000_0000_0000;
array[62548] <= 16'b0000_0000_0000_0000;
array[62549] <= 16'b0000_0000_0000_0000;
array[62550] <= 16'b0000_0000_0000_0000;
array[62551] <= 16'b0000_0000_0000_0000;
array[62552] <= 16'b0000_0000_0000_0000;
array[62553] <= 16'b0000_0000_0000_0000;
array[62554] <= 16'b0000_0000_0000_0000;
array[62555] <= 16'b0000_0000_0000_0000;
array[62556] <= 16'b0000_0000_0000_0000;
array[62557] <= 16'b0000_0000_0000_0000;
array[62558] <= 16'b0000_0000_0000_0000;
array[62559] <= 16'b0000_0000_0000_0000;
array[62560] <= 16'b0000_0000_0000_0000;
array[62561] <= 16'b0000_0000_0000_0000;
array[62562] <= 16'b0000_0000_0000_0000;
array[62563] <= 16'b0000_0000_0000_0000;
array[62564] <= 16'b0000_0000_0000_0000;
array[62565] <= 16'b0000_0000_0000_0000;
array[62566] <= 16'b0000_0000_0000_0000;
array[62567] <= 16'b0000_0000_0000_0000;
array[62568] <= 16'b0000_0000_0000_0000;
array[62569] <= 16'b0000_0000_0000_0000;
array[62570] <= 16'b0000_0000_0000_0000;
array[62571] <= 16'b0000_0000_0000_0000;
array[62572] <= 16'b0000_0000_0000_0000;
array[62573] <= 16'b0000_0000_0000_0000;
array[62574] <= 16'b0000_0000_0000_0000;
array[62575] <= 16'b0000_0000_0000_0000;
array[62576] <= 16'b0000_0000_0000_0000;
array[62577] <= 16'b0000_0000_0000_0000;
array[62578] <= 16'b0000_0000_0000_0000;
array[62579] <= 16'b0000_0000_0000_0000;
array[62580] <= 16'b0000_0000_0000_0000;
array[62581] <= 16'b0000_0000_0000_0000;
array[62582] <= 16'b0000_0000_0000_0000;
array[62583] <= 16'b0000_0000_0000_0000;
array[62584] <= 16'b0000_0000_0000_0000;
array[62585] <= 16'b0000_0000_0000_0000;
array[62586] <= 16'b0000_0000_0000_0000;
array[62587] <= 16'b0000_0000_0000_0000;
array[62588] <= 16'b0000_0000_0000_0000;
array[62589] <= 16'b0000_0000_0000_0000;
array[62590] <= 16'b0000_0000_0000_0000;
array[62591] <= 16'b0000_0000_0000_0000;
array[62592] <= 16'b0000_0000_0000_0000;
array[62593] <= 16'b0000_0000_0000_0000;
array[62594] <= 16'b0000_0000_0000_0000;
array[62595] <= 16'b0000_0000_0000_0000;
array[62596] <= 16'b0000_0000_0000_0000;
array[62597] <= 16'b0000_0000_0000_0000;
array[62598] <= 16'b0000_0000_0000_0000;
array[62599] <= 16'b0000_0000_0000_0000;
array[62600] <= 16'b0000_0000_0000_0000;
array[62601] <= 16'b0000_0000_0000_0000;
array[62602] <= 16'b0000_0000_0000_0000;
array[62603] <= 16'b0000_0000_0000_0000;
array[62604] <= 16'b0000_0000_0000_0000;
array[62605] <= 16'b0000_0000_0000_0000;
array[62606] <= 16'b0000_0000_0000_0000;
array[62607] <= 16'b0000_0000_0000_0000;
array[62608] <= 16'b0000_0000_0000_0000;
array[62609] <= 16'b0000_0000_0000_0000;
array[62610] <= 16'b0000_0000_0000_0000;
array[62611] <= 16'b0000_0000_0000_0000;
array[62612] <= 16'b0000_0000_0000_0000;
array[62613] <= 16'b0000_0000_0000_0000;
array[62614] <= 16'b0000_0000_0000_0000;
array[62615] <= 16'b0000_0000_0000_0000;
array[62616] <= 16'b0000_0000_0000_0000;
array[62617] <= 16'b0000_0000_0000_0000;
array[62618] <= 16'b0000_0000_0000_0000;
array[62619] <= 16'b0000_0000_0000_0000;
array[62620] <= 16'b0000_0000_0000_0000;
array[62621] <= 16'b0000_0000_0000_0000;
array[62622] <= 16'b0000_0000_0000_0000;
array[62623] <= 16'b0000_0000_0000_0000;
array[62624] <= 16'b0000_0000_0000_0000;
array[62625] <= 16'b0000_0000_0000_0000;
array[62626] <= 16'b0000_0000_0000_0000;
array[62627] <= 16'b0000_0000_0000_0000;
array[62628] <= 16'b0000_0000_0000_0000;
array[62629] <= 16'b0000_0000_0000_0000;
array[62630] <= 16'b0000_0000_0000_0000;
array[62631] <= 16'b0000_0000_0000_0000;
array[62632] <= 16'b0000_0000_0000_0000;
array[62633] <= 16'b0000_0000_0000_0000;
array[62634] <= 16'b0000_0000_0000_0000;
array[62635] <= 16'b0000_0000_0000_0000;
array[62636] <= 16'b0000_0000_0000_0000;
array[62637] <= 16'b0000_0000_0000_0000;
array[62638] <= 16'b0000_0000_0000_0000;
array[62639] <= 16'b0000_0000_0000_0000;
array[62640] <= 16'b0000_0000_0000_0000;
array[62641] <= 16'b0000_0000_0000_0000;
array[62642] <= 16'b0000_0000_0000_0000;
array[62643] <= 16'b0000_0000_0000_0000;
array[62644] <= 16'b0000_0000_0000_0000;
array[62645] <= 16'b0000_0000_0000_0000;
array[62646] <= 16'b0000_0000_0000_0000;
array[62647] <= 16'b0000_0000_0000_0000;
array[62648] <= 16'b0000_0000_0000_0000;
array[62649] <= 16'b0000_0000_0000_0000;
array[62650] <= 16'b0000_0000_0000_0000;
array[62651] <= 16'b0000_0000_0000_0000;
array[62652] <= 16'b0000_0000_0000_0000;
array[62653] <= 16'b0000_0000_0000_0000;
array[62654] <= 16'b0000_0000_0000_0000;
array[62655] <= 16'b0000_0000_0000_0000;
array[62656] <= 16'b0000_0000_0000_0000;
array[62657] <= 16'b0000_0000_0000_0000;
array[62658] <= 16'b0000_0000_0000_0000;
array[62659] <= 16'b0000_0000_0000_0000;
array[62660] <= 16'b0000_0000_0000_0000;
array[62661] <= 16'b0000_0000_0000_0000;
array[62662] <= 16'b0000_0000_0000_0000;
array[62663] <= 16'b0000_0000_0000_0000;
array[62664] <= 16'b0000_0000_0000_0000;
array[62665] <= 16'b0000_0000_0000_0000;
array[62666] <= 16'b0000_0000_0000_0000;
array[62667] <= 16'b0000_0000_0000_0000;
array[62668] <= 16'b0000_0000_0000_0000;
array[62669] <= 16'b0000_0000_0000_0000;
array[62670] <= 16'b0000_0000_0000_0000;
array[62671] <= 16'b0000_0000_0000_0000;
array[62672] <= 16'b0000_0000_0000_0000;
array[62673] <= 16'b0000_0000_0000_0000;
array[62674] <= 16'b0000_0000_0000_0000;
array[62675] <= 16'b0000_0000_0000_0000;
array[62676] <= 16'b0000_0000_0000_0000;
array[62677] <= 16'b0000_0000_0000_0000;
array[62678] <= 16'b0000_0000_0000_0000;
array[62679] <= 16'b0000_0000_0000_0000;
array[62680] <= 16'b0000_0000_0000_0000;
array[62681] <= 16'b0000_0000_0000_0000;
array[62682] <= 16'b0000_0000_0000_0000;
array[62683] <= 16'b0000_0000_0000_0000;
array[62684] <= 16'b0000_0000_0000_0000;
array[62685] <= 16'b0000_0000_0000_0000;
array[62686] <= 16'b0000_0000_0000_0000;
array[62687] <= 16'b0000_0000_0000_0000;
array[62688] <= 16'b0000_0000_0000_0000;
array[62689] <= 16'b0000_0000_0000_0000;
array[62690] <= 16'b0000_0000_0000_0000;
array[62691] <= 16'b0000_0000_0000_0000;
array[62692] <= 16'b0000_0000_0000_0000;
array[62693] <= 16'b0000_0000_0000_0000;
array[62694] <= 16'b0000_0000_0000_0000;
array[62695] <= 16'b0000_0000_0000_0000;
array[62696] <= 16'b0000_0000_0000_0000;
array[62697] <= 16'b0000_0000_0000_0000;
array[62698] <= 16'b0000_0000_0000_0000;
array[62699] <= 16'b0000_0000_0000_0000;
array[62700] <= 16'b0000_0000_0000_0000;
array[62701] <= 16'b0000_0000_0000_0000;
array[62702] <= 16'b0000_0000_0000_0000;
array[62703] <= 16'b0000_0000_0000_0000;
array[62704] <= 16'b0000_0000_0000_0000;
array[62705] <= 16'b0000_0000_0000_0000;
array[62706] <= 16'b0000_0000_0000_0000;
array[62707] <= 16'b0000_0000_0000_0000;
array[62708] <= 16'b0000_0000_0000_0000;
array[62709] <= 16'b0000_0000_0000_0000;
array[62710] <= 16'b0000_0000_0000_0000;
array[62711] <= 16'b0000_0000_0000_0000;
array[62712] <= 16'b0000_0000_0000_0000;
array[62713] <= 16'b0000_0000_0000_0000;
array[62714] <= 16'b0000_0000_0000_0000;
array[62715] <= 16'b0000_0000_0000_0000;
array[62716] <= 16'b0000_0000_0000_0000;
array[62717] <= 16'b0000_0000_0000_0000;
array[62718] <= 16'b0000_0000_0000_0000;
array[62719] <= 16'b0000_0000_0000_0000;
array[62720] <= 16'b0000_0000_0000_0000;
array[62721] <= 16'b0000_0000_0000_0000;
array[62722] <= 16'b0000_0000_0000_0000;
array[62723] <= 16'b0000_0000_0000_0000;
array[62724] <= 16'b0000_0000_0000_0000;
array[62725] <= 16'b0000_0000_0000_0000;
array[62726] <= 16'b0000_0000_0000_0000;
array[62727] <= 16'b0000_0000_0000_0000;
array[62728] <= 16'b0000_0000_0000_0000;
array[62729] <= 16'b0000_0000_0000_0000;
array[62730] <= 16'b0000_0000_0000_0000;
array[62731] <= 16'b0000_0000_0000_0000;
array[62732] <= 16'b0000_0000_0000_0000;
array[62733] <= 16'b0000_0000_0000_0000;
array[62734] <= 16'b0000_0000_0000_0000;
array[62735] <= 16'b0000_0000_0000_0000;
array[62736] <= 16'b0000_0000_0000_0000;
array[62737] <= 16'b0000_0000_0000_0000;
array[62738] <= 16'b0000_0000_0000_0000;
array[62739] <= 16'b0000_0000_0000_0000;
array[62740] <= 16'b0000_0000_0000_0000;
array[62741] <= 16'b0000_0000_0000_0000;
array[62742] <= 16'b0000_0000_0000_0000;
array[62743] <= 16'b0000_0000_0000_0000;
array[62744] <= 16'b0000_0000_0000_0000;
array[62745] <= 16'b0000_0000_0000_0000;
array[62746] <= 16'b0000_0000_0000_0000;
array[62747] <= 16'b0000_0000_0000_0000;
array[62748] <= 16'b0000_0000_0000_0000;
array[62749] <= 16'b0000_0000_0000_0000;
array[62750] <= 16'b0000_0000_0000_0000;
array[62751] <= 16'b0000_0000_0000_0000;
array[62752] <= 16'b0000_0000_0000_0000;
array[62753] <= 16'b0000_0000_0000_0000;
array[62754] <= 16'b0000_0000_0000_0000;
array[62755] <= 16'b0000_0000_0000_0000;
array[62756] <= 16'b0000_0000_0000_0000;
array[62757] <= 16'b0000_0000_0000_0000;
array[62758] <= 16'b0000_0000_0000_0000;
array[62759] <= 16'b0000_0000_0000_0000;
array[62760] <= 16'b0000_0000_0000_0000;
array[62761] <= 16'b0000_0000_0000_0000;
array[62762] <= 16'b0000_0000_0000_0000;
array[62763] <= 16'b0000_0000_0000_0000;
array[62764] <= 16'b0000_0000_0000_0000;
array[62765] <= 16'b0000_0000_0000_0000;
array[62766] <= 16'b0000_0000_0000_0000;
array[62767] <= 16'b0000_0000_0000_0000;
array[62768] <= 16'b0000_0000_0000_0000;
array[62769] <= 16'b0000_0000_0000_0000;
array[62770] <= 16'b0000_0000_0000_0000;
array[62771] <= 16'b0000_0000_0000_0000;
array[62772] <= 16'b0000_0000_0000_0000;
array[62773] <= 16'b0000_0000_0000_0000;
array[62774] <= 16'b0000_0000_0000_0000;
array[62775] <= 16'b0000_0000_0000_0000;
array[62776] <= 16'b0000_0000_0000_0000;
array[62777] <= 16'b0000_0000_0000_0000;
array[62778] <= 16'b0000_0000_0000_0000;
array[62779] <= 16'b0000_0000_0000_0000;
array[62780] <= 16'b0000_0000_0000_0000;
array[62781] <= 16'b0000_0000_0000_0000;
array[62782] <= 16'b0000_0000_0000_0000;
array[62783] <= 16'b0000_0000_0000_0000;
array[62784] <= 16'b0000_0000_0000_0000;
array[62785] <= 16'b0000_0000_0000_0000;
array[62786] <= 16'b0000_0000_0000_0000;
array[62787] <= 16'b0000_0000_0000_0000;
array[62788] <= 16'b0000_0000_0000_0000;
array[62789] <= 16'b0000_0000_0000_0000;
array[62790] <= 16'b0000_0000_0000_0000;
array[62791] <= 16'b0000_0000_0000_0000;
array[62792] <= 16'b0000_0000_0000_0000;
array[62793] <= 16'b0000_0000_0000_0000;
array[62794] <= 16'b0000_0000_0000_0000;
array[62795] <= 16'b0000_0000_0000_0000;
array[62796] <= 16'b0000_0000_0000_0000;
array[62797] <= 16'b0000_0000_0000_0000;
array[62798] <= 16'b0000_0000_0000_0000;
array[62799] <= 16'b0000_0000_0000_0000;
array[62800] <= 16'b0000_0000_0000_0000;
array[62801] <= 16'b0000_0000_0000_0000;
array[62802] <= 16'b0000_0000_0000_0000;
array[62803] <= 16'b0000_0000_0000_0000;
array[62804] <= 16'b0000_0000_0000_0000;
array[62805] <= 16'b0000_0000_0000_0000;
array[62806] <= 16'b0000_0000_0000_0000;
array[62807] <= 16'b0000_0000_0000_0000;
array[62808] <= 16'b0000_0000_0000_0000;
array[62809] <= 16'b0000_0000_0000_0000;
array[62810] <= 16'b0000_0000_0000_0000;
array[62811] <= 16'b0000_0000_0000_0000;
array[62812] <= 16'b0000_0000_0000_0000;
array[62813] <= 16'b0000_0000_0000_0000;
array[62814] <= 16'b0000_0000_0000_0000;
array[62815] <= 16'b0000_0000_0000_0000;
array[62816] <= 16'b0000_0000_0000_0000;
array[62817] <= 16'b0000_0000_0000_0000;
array[62818] <= 16'b0000_0000_0000_0000;
array[62819] <= 16'b0000_0000_0000_0000;
array[62820] <= 16'b0000_0000_0000_0000;
array[62821] <= 16'b0000_0000_0000_0000;
array[62822] <= 16'b0000_0000_0000_0000;
array[62823] <= 16'b0000_0000_0000_0000;
array[62824] <= 16'b0000_0000_0000_0000;
array[62825] <= 16'b0000_0000_0000_0000;
array[62826] <= 16'b0000_0000_0000_0000;
array[62827] <= 16'b0000_0000_0000_0000;
array[62828] <= 16'b0000_0000_0000_0000;
array[62829] <= 16'b0000_0000_0000_0000;
array[62830] <= 16'b0000_0000_0000_0000;
array[62831] <= 16'b0000_0000_0000_0000;
array[62832] <= 16'b0000_0000_0000_0000;
array[62833] <= 16'b0000_0000_0000_0000;
array[62834] <= 16'b0000_0000_0000_0000;
array[62835] <= 16'b0000_0000_0000_0000;
array[62836] <= 16'b0000_0000_0000_0000;
array[62837] <= 16'b0000_0000_0000_0000;
array[62838] <= 16'b0000_0000_0000_0000;
array[62839] <= 16'b0000_0000_0000_0000;
array[62840] <= 16'b0000_0000_0000_0000;
array[62841] <= 16'b0000_0000_0000_0000;
array[62842] <= 16'b0000_0000_0000_0000;
array[62843] <= 16'b0000_0000_0000_0000;
array[62844] <= 16'b0000_0000_0000_0000;
array[62845] <= 16'b0000_0000_0000_0000;
array[62846] <= 16'b0000_0000_0000_0000;
array[62847] <= 16'b0000_0000_0000_0000;
array[62848] <= 16'b0000_0000_0000_0000;
array[62849] <= 16'b0000_0000_0000_0000;
array[62850] <= 16'b0000_0000_0000_0000;
array[62851] <= 16'b0000_0000_0000_0000;
array[62852] <= 16'b0000_0000_0000_0000;
array[62853] <= 16'b0000_0000_0000_0000;
array[62854] <= 16'b0000_0000_0000_0000;
array[62855] <= 16'b0000_0000_0000_0000;
array[62856] <= 16'b0000_0000_0000_0000;
array[62857] <= 16'b0000_0000_0000_0000;
array[62858] <= 16'b0000_0000_0000_0000;
array[62859] <= 16'b0000_0000_0000_0000;
array[62860] <= 16'b0000_0000_0000_0000;
array[62861] <= 16'b0000_0000_0000_0000;
array[62862] <= 16'b0000_0000_0000_0000;
array[62863] <= 16'b0000_0000_0000_0000;
array[62864] <= 16'b0000_0000_0000_0000;
array[62865] <= 16'b0000_0000_0000_0000;
array[62866] <= 16'b0000_0000_0000_0000;
array[62867] <= 16'b0000_0000_0000_0000;
array[62868] <= 16'b0000_0000_0000_0000;
array[62869] <= 16'b0000_0000_0000_0000;
array[62870] <= 16'b0000_0000_0000_0000;
array[62871] <= 16'b0000_0000_0000_0000;
array[62872] <= 16'b0000_0000_0000_0000;
array[62873] <= 16'b0000_0000_0000_0000;
array[62874] <= 16'b0000_0000_0000_0000;
array[62875] <= 16'b0000_0000_0000_0000;
array[62876] <= 16'b0000_0000_0000_0000;
array[62877] <= 16'b0000_0000_0000_0000;
array[62878] <= 16'b0000_0000_0000_0000;
array[62879] <= 16'b0000_0000_0000_0000;
array[62880] <= 16'b0000_0000_0000_0000;
array[62881] <= 16'b0000_0000_0000_0000;
array[62882] <= 16'b0000_0000_0000_0000;
array[62883] <= 16'b0000_0000_0000_0000;
array[62884] <= 16'b0000_0000_0000_0000;
array[62885] <= 16'b0000_0000_0000_0000;
array[62886] <= 16'b0000_0000_0000_0000;
array[62887] <= 16'b0000_0000_0000_0000;
array[62888] <= 16'b0000_0000_0000_0000;
array[62889] <= 16'b0000_0000_0000_0000;
array[62890] <= 16'b0000_0000_0000_0000;
array[62891] <= 16'b0000_0000_0000_0000;
array[62892] <= 16'b0000_0000_0000_0000;
array[62893] <= 16'b0000_0000_0000_0000;
array[62894] <= 16'b0000_0000_0000_0000;
array[62895] <= 16'b0000_0000_0000_0000;
array[62896] <= 16'b0000_0000_0000_0000;
array[62897] <= 16'b0000_0000_0000_0000;
array[62898] <= 16'b0000_0000_0000_0000;
array[62899] <= 16'b0000_0000_0000_0000;
array[62900] <= 16'b0000_0000_0000_0000;
array[62901] <= 16'b0000_0000_0000_0000;
array[62902] <= 16'b0000_0000_0000_0000;
array[62903] <= 16'b0000_0000_0000_0000;
array[62904] <= 16'b0000_0000_0000_0000;
array[62905] <= 16'b0000_0000_0000_0000;
array[62906] <= 16'b0000_0000_0000_0000;
array[62907] <= 16'b0000_0000_0000_0000;
array[62908] <= 16'b0000_0000_0000_0000;
array[62909] <= 16'b0000_0000_0000_0000;
array[62910] <= 16'b0000_0000_0000_0000;
array[62911] <= 16'b0000_0000_0000_0000;
array[62912] <= 16'b0000_0000_0000_0000;
array[62913] <= 16'b0000_0000_0000_0000;
array[62914] <= 16'b0000_0000_0000_0000;
array[62915] <= 16'b0000_0000_0000_0000;
array[62916] <= 16'b0000_0000_0000_0000;
array[62917] <= 16'b0000_0000_0000_0000;
array[62918] <= 16'b0000_0000_0000_0000;
array[62919] <= 16'b0000_0000_0000_0000;
array[62920] <= 16'b0000_0000_0000_0000;
array[62921] <= 16'b0000_0000_0000_0000;
array[62922] <= 16'b0000_0000_0000_0000;
array[62923] <= 16'b0000_0000_0000_0000;
array[62924] <= 16'b0000_0000_0000_0000;
array[62925] <= 16'b0000_0000_0000_0000;
array[62926] <= 16'b0000_0000_0000_0000;
array[62927] <= 16'b0000_0000_0000_0000;
array[62928] <= 16'b0000_0000_0000_0000;
array[62929] <= 16'b0000_0000_0000_0000;
array[62930] <= 16'b0000_0000_0000_0000;
array[62931] <= 16'b0000_0000_0000_0000;
array[62932] <= 16'b0000_0000_0000_0000;
array[62933] <= 16'b0000_0000_0000_0000;
array[62934] <= 16'b0000_0000_0000_0000;
array[62935] <= 16'b0000_0000_0000_0000;
array[62936] <= 16'b0000_0000_0000_0000;
array[62937] <= 16'b0000_0000_0000_0000;
array[62938] <= 16'b0000_0000_0000_0000;
array[62939] <= 16'b0000_0000_0000_0000;
array[62940] <= 16'b0000_0000_0000_0000;
array[62941] <= 16'b0000_0000_0000_0000;
array[62942] <= 16'b0000_0000_0000_0000;
array[62943] <= 16'b0000_0000_0000_0000;
array[62944] <= 16'b0000_0000_0000_0000;
array[62945] <= 16'b0000_0000_0000_0000;
array[62946] <= 16'b0000_0000_0000_0000;
array[62947] <= 16'b0000_0000_0000_0000;
array[62948] <= 16'b0000_0000_0000_0000;
array[62949] <= 16'b0000_0000_0000_0000;
array[62950] <= 16'b0000_0000_0000_0000;
array[62951] <= 16'b0000_0000_0000_0000;
array[62952] <= 16'b0000_0000_0000_0000;
array[62953] <= 16'b0000_0000_0000_0000;
array[62954] <= 16'b0000_0000_0000_0000;
array[62955] <= 16'b0000_0000_0000_0000;
array[62956] <= 16'b0000_0000_0000_0000;
array[62957] <= 16'b0000_0000_0000_0000;
array[62958] <= 16'b0000_0000_0000_0000;
array[62959] <= 16'b0000_0000_0000_0000;
array[62960] <= 16'b0000_0000_0000_0000;
array[62961] <= 16'b0000_0000_0000_0000;
array[62962] <= 16'b0000_0000_0000_0000;
array[62963] <= 16'b0000_0000_0000_0000;
array[62964] <= 16'b0000_0000_0000_0000;
array[62965] <= 16'b0000_0000_0000_0000;
array[62966] <= 16'b0000_0000_0000_0000;
array[62967] <= 16'b0000_0000_0000_0000;
array[62968] <= 16'b0000_0000_0000_0000;
array[62969] <= 16'b0000_0000_0000_0000;
array[62970] <= 16'b0000_0000_0000_0000;
array[62971] <= 16'b0000_0000_0000_0000;
array[62972] <= 16'b0000_0000_0000_0000;
array[62973] <= 16'b0000_0000_0000_0000;
array[62974] <= 16'b0000_0000_0000_0000;
array[62975] <= 16'b0000_0000_0000_0000;
array[62976] <= 16'b0000_0000_0000_0000;
array[62977] <= 16'b0000_0000_0000_0000;
array[62978] <= 16'b0000_0000_0000_0000;
array[62979] <= 16'b0000_0000_0000_0000;
array[62980] <= 16'b0000_0000_0000_0000;
array[62981] <= 16'b0000_0000_0000_0000;
array[62982] <= 16'b0000_0000_0000_0000;
array[62983] <= 16'b0000_0000_0000_0000;
array[62984] <= 16'b0000_0000_0000_0000;
array[62985] <= 16'b0000_0000_0000_0000;
array[62986] <= 16'b0000_0000_0000_0000;
array[62987] <= 16'b0000_0000_0000_0000;
array[62988] <= 16'b0000_0000_0000_0000;
array[62989] <= 16'b0000_0000_0000_0000;
array[62990] <= 16'b0000_0000_0000_0000;
array[62991] <= 16'b0000_0000_0000_0000;
array[62992] <= 16'b0000_0000_0000_0000;
array[62993] <= 16'b0000_0000_0000_0000;
array[62994] <= 16'b0000_0000_0000_0000;
array[62995] <= 16'b0000_0000_0000_0000;
array[62996] <= 16'b0000_0000_0000_0000;
array[62997] <= 16'b0000_0000_0000_0000;
array[62998] <= 16'b0000_0000_0000_0000;
array[62999] <= 16'b0000_0000_0000_0000;
array[63000] <= 16'b0000_0000_0000_0000;
array[63001] <= 16'b0000_0000_0000_0000;
array[63002] <= 16'b0000_0000_0000_0000;
array[63003] <= 16'b0000_0000_0000_0000;
array[63004] <= 16'b0000_0000_0000_0000;
array[63005] <= 16'b0000_0000_0000_0000;
array[63006] <= 16'b0000_0000_0000_0000;
array[63007] <= 16'b0000_0000_0000_0000;
array[63008] <= 16'b0000_0000_0000_0000;
array[63009] <= 16'b0000_0000_0000_0000;
array[63010] <= 16'b0000_0000_0000_0000;
array[63011] <= 16'b0000_0000_0000_0000;
array[63012] <= 16'b0000_0000_0000_0000;
array[63013] <= 16'b0000_0000_0000_0000;
array[63014] <= 16'b0000_0000_0000_0000;
array[63015] <= 16'b0000_0000_0000_0000;
array[63016] <= 16'b0000_0000_0000_0000;
array[63017] <= 16'b0000_0000_0000_0000;
array[63018] <= 16'b0000_0000_0000_0000;
array[63019] <= 16'b0000_0000_0000_0000;
array[63020] <= 16'b0000_0000_0000_0000;
array[63021] <= 16'b0000_0000_0000_0000;
array[63022] <= 16'b0000_0000_0000_0000;
array[63023] <= 16'b0000_0000_0000_0000;
array[63024] <= 16'b0000_0000_0000_0000;
array[63025] <= 16'b0000_0000_0000_0000;
array[63026] <= 16'b0000_0000_0000_0000;
array[63027] <= 16'b0000_0000_0000_0000;
array[63028] <= 16'b0000_0000_0000_0000;
array[63029] <= 16'b0000_0000_0000_0000;
array[63030] <= 16'b0000_0000_0000_0000;
array[63031] <= 16'b0000_0000_0000_0000;
array[63032] <= 16'b0000_0000_0000_0000;
array[63033] <= 16'b0000_0000_0000_0000;
array[63034] <= 16'b0000_0000_0000_0000;
array[63035] <= 16'b0000_0000_0000_0000;
array[63036] <= 16'b0000_0000_0000_0000;
array[63037] <= 16'b0000_0000_0000_0000;
array[63038] <= 16'b0000_0000_0000_0000;
array[63039] <= 16'b0000_0000_0000_0000;
array[63040] <= 16'b0000_0000_0000_0000;
array[63041] <= 16'b0000_0000_0000_0000;
array[63042] <= 16'b0000_0000_0000_0000;
array[63043] <= 16'b0000_0000_0000_0000;
array[63044] <= 16'b0000_0000_0000_0000;
array[63045] <= 16'b0000_0000_0000_0000;
array[63046] <= 16'b0000_0000_0000_0000;
array[63047] <= 16'b0000_0000_0000_0000;
array[63048] <= 16'b0000_0000_0000_0000;
array[63049] <= 16'b0000_0000_0000_0000;
array[63050] <= 16'b0000_0000_0000_0000;
array[63051] <= 16'b0000_0000_0000_0000;
array[63052] <= 16'b0000_0000_0000_0000;
array[63053] <= 16'b0000_0000_0000_0000;
array[63054] <= 16'b0000_0000_0000_0000;
array[63055] <= 16'b0000_0000_0000_0000;
array[63056] <= 16'b0000_0000_0000_0000;
array[63057] <= 16'b0000_0000_0000_0000;
array[63058] <= 16'b0000_0000_0000_0000;
array[63059] <= 16'b0000_0000_0000_0000;
array[63060] <= 16'b0000_0000_0000_0000;
array[63061] <= 16'b0000_0000_0000_0000;
array[63062] <= 16'b0000_0000_0000_0000;
array[63063] <= 16'b0000_0000_0000_0000;
array[63064] <= 16'b0000_0000_0000_0000;
array[63065] <= 16'b0000_0000_0000_0000;
array[63066] <= 16'b0000_0000_0000_0000;
array[63067] <= 16'b0000_0000_0000_0000;
array[63068] <= 16'b0000_0000_0000_0000;
array[63069] <= 16'b0000_0000_0000_0000;
array[63070] <= 16'b0000_0000_0000_0000;
array[63071] <= 16'b0000_0000_0000_0000;
array[63072] <= 16'b0000_0000_0000_0000;
array[63073] <= 16'b0000_0000_0000_0000;
array[63074] <= 16'b0000_0000_0000_0000;
array[63075] <= 16'b0000_0000_0000_0000;
array[63076] <= 16'b0000_0000_0000_0000;
array[63077] <= 16'b0000_0000_0000_0000;
array[63078] <= 16'b0000_0000_0000_0000;
array[63079] <= 16'b0000_0000_0000_0000;
array[63080] <= 16'b0000_0000_0000_0000;
array[63081] <= 16'b0000_0000_0000_0000;
array[63082] <= 16'b0000_0000_0000_0000;
array[63083] <= 16'b0000_0000_0000_0000;
array[63084] <= 16'b0000_0000_0000_0000;
array[63085] <= 16'b0000_0000_0000_0000;
array[63086] <= 16'b0000_0000_0000_0000;
array[63087] <= 16'b0000_0000_0000_0000;
array[63088] <= 16'b0000_0000_0000_0000;
array[63089] <= 16'b0000_0000_0000_0000;
array[63090] <= 16'b0000_0000_0000_0000;
array[63091] <= 16'b0000_0000_0000_0000;
array[63092] <= 16'b0000_0000_0000_0000;
array[63093] <= 16'b0000_0000_0000_0000;
array[63094] <= 16'b0000_0000_0000_0000;
array[63095] <= 16'b0000_0000_0000_0000;
array[63096] <= 16'b0000_0000_0000_0000;
array[63097] <= 16'b0000_0000_0000_0000;
array[63098] <= 16'b0000_0000_0000_0000;
array[63099] <= 16'b0000_0000_0000_0000;
array[63100] <= 16'b0000_0000_0000_0000;
array[63101] <= 16'b0000_0000_0000_0000;
array[63102] <= 16'b0000_0000_0000_0000;
array[63103] <= 16'b0000_0000_0000_0000;
array[63104] <= 16'b0000_0000_0000_0000;
array[63105] <= 16'b0000_0000_0000_0000;
array[63106] <= 16'b0000_0000_0000_0000;
array[63107] <= 16'b0000_0000_0000_0000;
array[63108] <= 16'b0000_0000_0000_0000;
array[63109] <= 16'b0000_0000_0000_0000;
array[63110] <= 16'b0000_0000_0000_0000;
array[63111] <= 16'b0000_0000_0000_0000;
array[63112] <= 16'b0000_0000_0000_0000;
array[63113] <= 16'b0000_0000_0000_0000;
array[63114] <= 16'b0000_0000_0000_0000;
array[63115] <= 16'b0000_0000_0000_0000;
array[63116] <= 16'b0000_0000_0000_0000;
array[63117] <= 16'b0000_0000_0000_0000;
array[63118] <= 16'b0000_0000_0000_0000;
array[63119] <= 16'b0000_0000_0000_0000;
array[63120] <= 16'b0000_0000_0000_0000;
array[63121] <= 16'b0000_0000_0000_0000;
array[63122] <= 16'b0000_0000_0000_0000;
array[63123] <= 16'b0000_0000_0000_0000;
array[63124] <= 16'b0000_0000_0000_0000;
array[63125] <= 16'b0000_0000_0000_0000;
array[63126] <= 16'b0000_0000_0000_0000;
array[63127] <= 16'b0000_0000_0000_0000;
array[63128] <= 16'b0000_0000_0000_0000;
array[63129] <= 16'b0000_0000_0000_0000;
array[63130] <= 16'b0000_0000_0000_0000;
array[63131] <= 16'b0000_0000_0000_0000;
array[63132] <= 16'b0000_0000_0000_0000;
array[63133] <= 16'b0000_0000_0000_0000;
array[63134] <= 16'b0000_0000_0000_0000;
array[63135] <= 16'b0000_0000_0000_0000;
array[63136] <= 16'b0000_0000_0000_0000;
array[63137] <= 16'b0000_0000_0000_0000;
array[63138] <= 16'b0000_0000_0000_0000;
array[63139] <= 16'b0000_0000_0000_0000;
array[63140] <= 16'b0000_0000_0000_0000;
array[63141] <= 16'b0000_0000_0000_0000;
array[63142] <= 16'b0000_0000_0000_0000;
array[63143] <= 16'b0000_0000_0000_0000;
array[63144] <= 16'b0000_0000_0000_0000;
array[63145] <= 16'b0000_0000_0000_0000;
array[63146] <= 16'b0000_0000_0000_0000;
array[63147] <= 16'b0000_0000_0000_0000;
array[63148] <= 16'b0000_0000_0000_0000;
array[63149] <= 16'b0000_0000_0000_0000;
array[63150] <= 16'b0000_0000_0000_0000;
array[63151] <= 16'b0000_0000_0000_0000;
array[63152] <= 16'b0000_0000_0000_0000;
array[63153] <= 16'b0000_0000_0000_0000;
array[63154] <= 16'b0000_0000_0000_0000;
array[63155] <= 16'b0000_0000_0000_0000;
array[63156] <= 16'b0000_0000_0000_0000;
array[63157] <= 16'b0000_0000_0000_0000;
array[63158] <= 16'b0000_0000_0000_0000;
array[63159] <= 16'b0000_0000_0000_0000;
array[63160] <= 16'b0000_0000_0000_0000;
array[63161] <= 16'b0000_0000_0000_0000;
array[63162] <= 16'b0000_0000_0000_0000;
array[63163] <= 16'b0000_0000_0000_0000;
array[63164] <= 16'b0000_0000_0000_0000;
array[63165] <= 16'b0000_0000_0000_0000;
array[63166] <= 16'b0000_0000_0000_0000;
array[63167] <= 16'b0000_0000_0000_0000;
array[63168] <= 16'b0000_0000_0000_0000;
array[63169] <= 16'b0000_0000_0000_0000;
array[63170] <= 16'b0000_0000_0000_0000;
array[63171] <= 16'b0000_0000_0000_0000;
array[63172] <= 16'b0000_0000_0000_0000;
array[63173] <= 16'b0000_0000_0000_0000;
array[63174] <= 16'b0000_0000_0000_0000;
array[63175] <= 16'b0000_0000_0000_0000;
array[63176] <= 16'b0000_0000_0000_0000;
array[63177] <= 16'b0000_0000_0000_0000;
array[63178] <= 16'b0000_0000_0000_0000;
array[63179] <= 16'b0000_0000_0000_0000;
array[63180] <= 16'b0000_0000_0000_0000;
array[63181] <= 16'b0000_0000_0000_0000;
array[63182] <= 16'b0000_0000_0000_0000;
array[63183] <= 16'b0000_0000_0000_0000;
array[63184] <= 16'b0000_0000_0000_0000;
array[63185] <= 16'b0000_0000_0000_0000;
array[63186] <= 16'b0000_0000_0000_0000;
array[63187] <= 16'b0000_0000_0000_0000;
array[63188] <= 16'b0000_0000_0000_0000;
array[63189] <= 16'b0000_0000_0000_0000;
array[63190] <= 16'b0000_0000_0000_0000;
array[63191] <= 16'b0000_0000_0000_0000;
array[63192] <= 16'b0000_0000_0000_0000;
array[63193] <= 16'b0000_0000_0000_0000;
array[63194] <= 16'b0000_0000_0000_0000;
array[63195] <= 16'b0000_0000_0000_0000;
array[63196] <= 16'b0000_0000_0000_0000;
array[63197] <= 16'b0000_0000_0000_0000;
array[63198] <= 16'b0000_0000_0000_0000;
array[63199] <= 16'b0000_0000_0000_0000;
array[63200] <= 16'b0000_0000_0000_0000;
array[63201] <= 16'b0000_0000_0000_0000;
array[63202] <= 16'b0000_0000_0000_0000;
array[63203] <= 16'b0000_0000_0000_0000;
array[63204] <= 16'b0000_0000_0000_0000;
array[63205] <= 16'b0000_0000_0000_0000;
array[63206] <= 16'b0000_0000_0000_0000;
array[63207] <= 16'b0000_0000_0000_0000;
array[63208] <= 16'b0000_0000_0000_0000;
array[63209] <= 16'b0000_0000_0000_0000;
array[63210] <= 16'b0000_0000_0000_0000;
array[63211] <= 16'b0000_0000_0000_0000;
array[63212] <= 16'b0000_0000_0000_0000;
array[63213] <= 16'b0000_0000_0000_0000;
array[63214] <= 16'b0000_0000_0000_0000;
array[63215] <= 16'b0000_0000_0000_0000;
array[63216] <= 16'b0000_0000_0000_0000;
array[63217] <= 16'b0000_0000_0000_0000;
array[63218] <= 16'b0000_0000_0000_0000;
array[63219] <= 16'b0000_0000_0000_0000;
array[63220] <= 16'b0000_0000_0000_0000;
array[63221] <= 16'b0000_0000_0000_0000;
array[63222] <= 16'b0000_0000_0000_0000;
array[63223] <= 16'b0000_0000_0000_0000;
array[63224] <= 16'b0000_0000_0000_0000;
array[63225] <= 16'b0000_0000_0000_0000;
array[63226] <= 16'b0000_0000_0000_0000;
array[63227] <= 16'b0000_0000_0000_0000;
array[63228] <= 16'b0000_0000_0000_0000;
array[63229] <= 16'b0000_0000_0000_0000;
array[63230] <= 16'b0000_0000_0000_0000;
array[63231] <= 16'b0000_0000_0000_0000;
array[63232] <= 16'b0000_0000_0000_0000;
array[63233] <= 16'b0000_0000_0000_0000;
array[63234] <= 16'b0000_0000_0000_0000;
array[63235] <= 16'b0000_0000_0000_0000;
array[63236] <= 16'b0000_0000_0000_0000;
array[63237] <= 16'b0000_0000_0000_0000;
array[63238] <= 16'b0000_0000_0000_0000;
array[63239] <= 16'b0000_0000_0000_0000;
array[63240] <= 16'b0000_0000_0000_0000;
array[63241] <= 16'b0000_0000_0000_0000;
array[63242] <= 16'b0000_0000_0000_0000;
array[63243] <= 16'b0000_0000_0000_0000;
array[63244] <= 16'b0000_0000_0000_0000;
array[63245] <= 16'b0000_0000_0000_0000;
array[63246] <= 16'b0000_0000_0000_0000;
array[63247] <= 16'b0000_0000_0000_0000;
array[63248] <= 16'b0000_0000_0000_0000;
array[63249] <= 16'b0000_0000_0000_0000;
array[63250] <= 16'b0000_0000_0000_0000;
array[63251] <= 16'b0000_0000_0000_0000;
array[63252] <= 16'b0000_0000_0000_0000;
array[63253] <= 16'b0000_0000_0000_0000;
array[63254] <= 16'b0000_0000_0000_0000;
array[63255] <= 16'b0000_0000_0000_0000;
array[63256] <= 16'b0000_0000_0000_0000;
array[63257] <= 16'b0000_0000_0000_0000;
array[63258] <= 16'b0000_0000_0000_0000;
array[63259] <= 16'b0000_0000_0000_0000;
array[63260] <= 16'b0000_0000_0000_0000;
array[63261] <= 16'b0000_0000_0000_0000;
array[63262] <= 16'b0000_0000_0000_0000;
array[63263] <= 16'b0000_0000_0000_0000;
array[63264] <= 16'b0000_0000_0000_0000;
array[63265] <= 16'b0000_0000_0000_0000;
array[63266] <= 16'b0000_0000_0000_0000;
array[63267] <= 16'b0000_0000_0000_0000;
array[63268] <= 16'b0000_0000_0000_0000;
array[63269] <= 16'b0000_0000_0000_0000;
array[63270] <= 16'b0000_0000_0000_0000;
array[63271] <= 16'b0000_0000_0000_0000;
array[63272] <= 16'b0000_0000_0000_0000;
array[63273] <= 16'b0000_0000_0000_0000;
array[63274] <= 16'b0000_0000_0000_0000;
array[63275] <= 16'b0000_0000_0000_0000;
array[63276] <= 16'b0000_0000_0000_0000;
array[63277] <= 16'b0000_0000_0000_0000;
array[63278] <= 16'b0000_0000_0000_0000;
array[63279] <= 16'b0000_0000_0000_0000;
array[63280] <= 16'b0000_0000_0000_0000;
array[63281] <= 16'b0000_0000_0000_0000;
array[63282] <= 16'b0000_0000_0000_0000;
array[63283] <= 16'b0000_0000_0000_0000;
array[63284] <= 16'b0000_0000_0000_0000;
array[63285] <= 16'b0000_0000_0000_0000;
array[63286] <= 16'b0000_0000_0000_0000;
array[63287] <= 16'b0000_0000_0000_0000;
array[63288] <= 16'b0000_0000_0000_0000;
array[63289] <= 16'b0000_0000_0000_0000;
array[63290] <= 16'b0000_0000_0000_0000;
array[63291] <= 16'b0000_0000_0000_0000;
array[63292] <= 16'b0000_0000_0000_0000;
array[63293] <= 16'b0000_0000_0000_0000;
array[63294] <= 16'b0000_0000_0000_0000;
array[63295] <= 16'b0000_0000_0000_0000;
array[63296] <= 16'b0000_0000_0000_0000;
array[63297] <= 16'b0000_0000_0000_0000;
array[63298] <= 16'b0000_0000_0000_0000;
array[63299] <= 16'b0000_0000_0000_0000;
array[63300] <= 16'b0000_0000_0000_0000;
array[63301] <= 16'b0000_0000_0000_0000;
array[63302] <= 16'b0000_0000_0000_0000;
array[63303] <= 16'b0000_0000_0000_0000;
array[63304] <= 16'b0000_0000_0000_0000;
array[63305] <= 16'b0000_0000_0000_0000;
array[63306] <= 16'b0000_0000_0000_0000;
array[63307] <= 16'b0000_0000_0000_0000;
array[63308] <= 16'b0000_0000_0000_0000;
array[63309] <= 16'b0000_0000_0000_0000;
array[63310] <= 16'b0000_0000_0000_0000;
array[63311] <= 16'b0000_0000_0000_0000;
array[63312] <= 16'b0000_0000_0000_0000;
array[63313] <= 16'b0000_0000_0000_0000;
array[63314] <= 16'b0000_0000_0000_0000;
array[63315] <= 16'b0000_0000_0000_0000;
array[63316] <= 16'b0000_0000_0000_0000;
array[63317] <= 16'b0000_0000_0000_0000;
array[63318] <= 16'b0000_0000_0000_0000;
array[63319] <= 16'b0000_0000_0000_0000;
array[63320] <= 16'b0000_0000_0000_0000;
array[63321] <= 16'b0000_0000_0000_0000;
array[63322] <= 16'b0000_0000_0000_0000;
array[63323] <= 16'b0000_0000_0000_0000;
array[63324] <= 16'b0000_0000_0000_0000;
array[63325] <= 16'b0000_0000_0000_0000;
array[63326] <= 16'b0000_0000_0000_0000;
array[63327] <= 16'b0000_0000_0000_0000;
array[63328] <= 16'b0000_0000_0000_0000;
array[63329] <= 16'b0000_0000_0000_0000;
array[63330] <= 16'b0000_0000_0000_0000;
array[63331] <= 16'b0000_0000_0000_0000;
array[63332] <= 16'b0000_0000_0000_0000;
array[63333] <= 16'b0000_0000_0000_0000;
array[63334] <= 16'b0000_0000_0000_0000;
array[63335] <= 16'b0000_0000_0000_0000;
array[63336] <= 16'b0000_0000_0000_0000;
array[63337] <= 16'b0000_0000_0000_0000;
array[63338] <= 16'b0000_0000_0000_0000;
array[63339] <= 16'b0000_0000_0000_0000;
array[63340] <= 16'b0000_0000_0000_0000;
array[63341] <= 16'b0000_0000_0000_0000;
array[63342] <= 16'b0000_0000_0000_0000;
array[63343] <= 16'b0000_0000_0000_0000;
array[63344] <= 16'b0000_0000_0000_0000;
array[63345] <= 16'b0000_0000_0000_0000;
array[63346] <= 16'b0000_0000_0000_0000;
array[63347] <= 16'b0000_0000_0000_0000;
array[63348] <= 16'b0000_0000_0000_0000;
array[63349] <= 16'b0000_0000_0000_0000;
array[63350] <= 16'b0000_0000_0000_0000;
array[63351] <= 16'b0000_0000_0000_0000;
array[63352] <= 16'b0000_0000_0000_0000;
array[63353] <= 16'b0000_0000_0000_0000;
array[63354] <= 16'b0000_0000_0000_0000;
array[63355] <= 16'b0000_0000_0000_0000;
array[63356] <= 16'b0000_0000_0000_0000;
array[63357] <= 16'b0000_0000_0000_0000;
array[63358] <= 16'b0000_0000_0000_0000;
array[63359] <= 16'b0000_0000_0000_0000;
array[63360] <= 16'b0000_0000_0000_0000;
array[63361] <= 16'b0000_0000_0000_0000;
array[63362] <= 16'b0000_0000_0000_0000;
array[63363] <= 16'b0000_0000_0000_0000;
array[63364] <= 16'b0000_0000_0000_0000;
array[63365] <= 16'b0000_0000_0000_0000;
array[63366] <= 16'b0000_0000_0000_0000;
array[63367] <= 16'b0000_0000_0000_0000;
array[63368] <= 16'b0000_0000_0000_0000;
array[63369] <= 16'b0000_0000_0000_0000;
array[63370] <= 16'b0000_0000_0000_0000;
array[63371] <= 16'b0000_0000_0000_0000;
array[63372] <= 16'b0000_0000_0000_0000;
array[63373] <= 16'b0000_0000_0000_0000;
array[63374] <= 16'b0000_0000_0000_0000;
array[63375] <= 16'b0000_0000_0000_0000;
array[63376] <= 16'b0000_0000_0000_0000;
array[63377] <= 16'b0000_0000_0000_0000;
array[63378] <= 16'b0000_0000_0000_0000;
array[63379] <= 16'b0000_0000_0000_0000;
array[63380] <= 16'b0000_0000_0000_0000;
array[63381] <= 16'b0000_0000_0000_0000;
array[63382] <= 16'b0000_0000_0000_0000;
array[63383] <= 16'b0000_0000_0000_0000;
array[63384] <= 16'b0000_0000_0000_0000;
array[63385] <= 16'b0000_0000_0000_0000;
array[63386] <= 16'b0000_0000_0000_0000;
array[63387] <= 16'b0000_0000_0000_0000;
array[63388] <= 16'b0000_0000_0000_0000;
array[63389] <= 16'b0000_0000_0000_0000;
array[63390] <= 16'b0000_0000_0000_0000;
array[63391] <= 16'b0000_0000_0000_0000;
array[63392] <= 16'b0000_0000_0000_0000;
array[63393] <= 16'b0000_0000_0000_0000;
array[63394] <= 16'b0000_0000_0000_0000;
array[63395] <= 16'b0000_0000_0000_0000;
array[63396] <= 16'b0000_0000_0000_0000;
array[63397] <= 16'b0000_0000_0000_0000;
array[63398] <= 16'b0000_0000_0000_0000;
array[63399] <= 16'b0000_0000_0000_0000;
array[63400] <= 16'b0000_0000_0000_0000;
array[63401] <= 16'b0000_0000_0000_0000;
array[63402] <= 16'b0000_0000_0000_0000;
array[63403] <= 16'b0000_0000_0000_0000;
array[63404] <= 16'b0000_0000_0000_0000;
array[63405] <= 16'b0000_0000_0000_0000;
array[63406] <= 16'b0000_0000_0000_0000;
array[63407] <= 16'b0000_0000_0000_0000;
array[63408] <= 16'b0000_0000_0000_0000;
array[63409] <= 16'b0000_0000_0000_0000;
array[63410] <= 16'b0000_0000_0000_0000;
array[63411] <= 16'b0000_0000_0000_0000;
array[63412] <= 16'b0000_0000_0000_0000;
array[63413] <= 16'b0000_0000_0000_0000;
array[63414] <= 16'b0000_0000_0000_0000;
array[63415] <= 16'b0000_0000_0000_0000;
array[63416] <= 16'b0000_0000_0000_0000;
array[63417] <= 16'b0000_0000_0000_0000;
array[63418] <= 16'b0000_0000_0000_0000;
array[63419] <= 16'b0000_0000_0000_0000;
array[63420] <= 16'b0000_0000_0000_0000;
array[63421] <= 16'b0000_0000_0000_0000;
array[63422] <= 16'b0000_0000_0000_0000;
array[63423] <= 16'b0000_0000_0000_0000;
array[63424] <= 16'b0000_0000_0000_0000;
array[63425] <= 16'b0000_0000_0000_0000;
array[63426] <= 16'b0000_0000_0000_0000;
array[63427] <= 16'b0000_0000_0000_0000;
array[63428] <= 16'b0000_0000_0000_0000;
array[63429] <= 16'b0000_0000_0000_0000;
array[63430] <= 16'b0000_0000_0000_0000;
array[63431] <= 16'b0000_0000_0000_0000;
array[63432] <= 16'b0000_0000_0000_0000;
array[63433] <= 16'b0000_0000_0000_0000;
array[63434] <= 16'b0000_0000_0000_0000;
array[63435] <= 16'b0000_0000_0000_0000;
array[63436] <= 16'b0000_0000_0000_0000;
array[63437] <= 16'b0000_0000_0000_0000;
array[63438] <= 16'b0000_0000_0000_0000;
array[63439] <= 16'b0000_0000_0000_0000;
array[63440] <= 16'b0000_0000_0000_0000;
array[63441] <= 16'b0000_0000_0000_0000;
array[63442] <= 16'b0000_0000_0000_0000;
array[63443] <= 16'b0000_0000_0000_0000;
array[63444] <= 16'b0000_0000_0000_0000;
array[63445] <= 16'b0000_0000_0000_0000;
array[63446] <= 16'b0000_0000_0000_0000;
array[63447] <= 16'b0000_0000_0000_0000;
array[63448] <= 16'b0000_0000_0000_0000;
array[63449] <= 16'b0000_0000_0000_0000;
array[63450] <= 16'b0000_0000_0000_0000;
array[63451] <= 16'b0000_0000_0000_0000;
array[63452] <= 16'b0000_0000_0000_0000;
array[63453] <= 16'b0000_0000_0000_0000;
array[63454] <= 16'b0000_0000_0000_0000;
array[63455] <= 16'b0000_0000_0000_0000;
array[63456] <= 16'b0000_0000_0000_0000;
array[63457] <= 16'b0000_0000_0000_0000;
array[63458] <= 16'b0000_0000_0000_0000;
array[63459] <= 16'b0000_0000_0000_0000;
array[63460] <= 16'b0000_0000_0000_0000;
array[63461] <= 16'b0000_0000_0000_0000;
array[63462] <= 16'b0000_0000_0000_0000;
array[63463] <= 16'b0000_0000_0000_0000;
array[63464] <= 16'b0000_0000_0000_0000;
array[63465] <= 16'b0000_0000_0000_0000;
array[63466] <= 16'b0000_0000_0000_0000;
array[63467] <= 16'b0000_0000_0000_0000;
array[63468] <= 16'b0000_0000_0000_0000;
array[63469] <= 16'b0000_0000_0000_0000;
array[63470] <= 16'b0000_0000_0000_0000;
array[63471] <= 16'b0000_0000_0000_0000;
array[63472] <= 16'b0000_0000_0000_0000;
array[63473] <= 16'b0000_0000_0000_0000;
array[63474] <= 16'b0000_0000_0000_0000;
array[63475] <= 16'b0000_0000_0000_0000;
array[63476] <= 16'b0000_0000_0000_0000;
array[63477] <= 16'b0000_0000_0000_0000;
array[63478] <= 16'b0000_0000_0000_0000;
array[63479] <= 16'b0000_0000_0000_0000;
array[63480] <= 16'b0000_0000_0000_0000;
array[63481] <= 16'b0000_0000_0000_0000;
array[63482] <= 16'b0000_0000_0000_0000;
array[63483] <= 16'b0000_0000_0000_0000;
array[63484] <= 16'b0000_0000_0000_0000;
array[63485] <= 16'b0000_0000_0000_0000;
array[63486] <= 16'b0000_0000_0000_0000;
array[63487] <= 16'b0000_0000_0000_0000;
array[63488] <= 16'b0000_0000_0000_0000;
array[63489] <= 16'b0000_0000_0000_0000;
array[63490] <= 16'b0000_0000_0000_0000;
array[63491] <= 16'b0000_0000_0000_0000;
array[63492] <= 16'b0000_0000_0000_0000;
array[63493] <= 16'b0000_0000_0000_0000;
array[63494] <= 16'b0000_0000_0000_0000;
array[63495] <= 16'b0000_0000_0000_0000;
array[63496] <= 16'b0000_0000_0000_0000;
array[63497] <= 16'b0000_0000_0000_0000;
array[63498] <= 16'b0000_0000_0000_0000;
array[63499] <= 16'b0000_0000_0000_0000;
array[63500] <= 16'b0000_0000_0000_0000;
array[63501] <= 16'b0000_0000_0000_0000;
array[63502] <= 16'b0000_0000_0000_0000;
array[63503] <= 16'b0000_0000_0000_0000;
array[63504] <= 16'b0000_0000_0000_0000;
array[63505] <= 16'b0000_0000_0000_0000;
array[63506] <= 16'b0000_0000_0000_0000;
array[63507] <= 16'b0000_0000_0000_0000;
array[63508] <= 16'b0000_0000_0000_0000;
array[63509] <= 16'b0000_0000_0000_0000;
array[63510] <= 16'b0000_0000_0000_0000;
array[63511] <= 16'b0000_0000_0000_0000;
array[63512] <= 16'b0000_0000_0000_0000;
array[63513] <= 16'b0000_0000_0000_0000;
array[63514] <= 16'b0000_0000_0000_0000;
array[63515] <= 16'b0000_0000_0000_0000;
array[63516] <= 16'b0000_0000_0000_0000;
array[63517] <= 16'b0000_0000_0000_0000;
array[63518] <= 16'b0000_0000_0000_0000;
array[63519] <= 16'b0000_0000_0000_0000;
array[63520] <= 16'b0000_0000_0000_0000;
array[63521] <= 16'b0000_0000_0000_0000;
array[63522] <= 16'b0000_0000_0000_0000;
array[63523] <= 16'b0000_0000_0000_0000;
array[63524] <= 16'b0000_0000_0000_0000;
array[63525] <= 16'b0000_0000_0000_0000;
array[63526] <= 16'b0000_0000_0000_0000;
array[63527] <= 16'b0000_0000_0000_0000;
array[63528] <= 16'b0000_0000_0000_0000;
array[63529] <= 16'b0000_0000_0000_0000;
array[63530] <= 16'b0000_0000_0000_0000;
array[63531] <= 16'b0000_0000_0000_0000;
array[63532] <= 16'b0000_0000_0000_0000;
array[63533] <= 16'b0000_0000_0000_0000;
array[63534] <= 16'b0000_0000_0000_0000;
array[63535] <= 16'b0000_0000_0000_0000;
array[63536] <= 16'b0000_0000_0000_0000;
array[63537] <= 16'b0000_0000_0000_0000;
array[63538] <= 16'b0000_0000_0000_0000;
array[63539] <= 16'b0000_0000_0000_0000;
array[63540] <= 16'b0000_0000_0000_0000;
array[63541] <= 16'b0000_0000_0000_0000;
array[63542] <= 16'b0000_0000_0000_0000;
array[63543] <= 16'b0000_0000_0000_0000;
array[63544] <= 16'b0000_0000_0000_0000;
array[63545] <= 16'b0000_0000_0000_0000;
array[63546] <= 16'b0000_0000_0000_0000;
array[63547] <= 16'b0000_0000_0000_0000;
array[63548] <= 16'b0000_0000_0000_0000;
array[63549] <= 16'b0000_0000_0000_0000;
array[63550] <= 16'b0000_0000_0000_0000;
array[63551] <= 16'b0000_0000_0000_0000;
array[63552] <= 16'b0000_0000_0000_0000;
array[63553] <= 16'b0000_0000_0000_0000;
array[63554] <= 16'b0000_0000_0000_0000;
array[63555] <= 16'b0000_0000_0000_0000;
array[63556] <= 16'b0000_0000_0000_0000;
array[63557] <= 16'b0000_0000_0000_0000;
array[63558] <= 16'b0000_0000_0000_0000;
array[63559] <= 16'b0000_0000_0000_0000;
array[63560] <= 16'b0000_0000_0000_0000;
array[63561] <= 16'b0000_0000_0000_0000;
array[63562] <= 16'b0000_0000_0000_0000;
array[63563] <= 16'b0000_0000_0000_0000;
array[63564] <= 16'b0000_0000_0000_0000;
array[63565] <= 16'b0000_0000_0000_0000;
array[63566] <= 16'b0000_0000_0000_0000;
array[63567] <= 16'b0000_0000_0000_0000;
array[63568] <= 16'b0000_0000_0000_0000;
array[63569] <= 16'b0000_0000_0000_0000;
array[63570] <= 16'b0000_0000_0000_0000;
array[63571] <= 16'b0000_0000_0000_0000;
array[63572] <= 16'b0000_0000_0000_0000;
array[63573] <= 16'b0000_0000_0000_0000;
array[63574] <= 16'b0000_0000_0000_0000;
array[63575] <= 16'b0000_0000_0000_0000;
array[63576] <= 16'b0000_0000_0000_0000;
array[63577] <= 16'b0000_0000_0000_0000;
array[63578] <= 16'b0000_0000_0000_0000;
array[63579] <= 16'b0000_0000_0000_0000;
array[63580] <= 16'b0000_0000_0000_0000;
array[63581] <= 16'b0000_0000_0000_0000;
array[63582] <= 16'b0000_0000_0000_0000;
array[63583] <= 16'b0000_0000_0000_0000;
array[63584] <= 16'b0000_0000_0000_0000;
array[63585] <= 16'b0000_0000_0000_0000;
array[63586] <= 16'b0000_0000_0000_0000;
array[63587] <= 16'b0000_0000_0000_0000;
array[63588] <= 16'b0000_0000_0000_0000;
array[63589] <= 16'b0000_0000_0000_0000;
array[63590] <= 16'b0000_0000_0000_0000;
array[63591] <= 16'b0000_0000_0000_0000;
array[63592] <= 16'b0000_0000_0000_0000;
array[63593] <= 16'b0000_0000_0000_0000;
array[63594] <= 16'b0000_0000_0000_0000;
array[63595] <= 16'b0000_0000_0000_0000;
array[63596] <= 16'b0000_0000_0000_0000;
array[63597] <= 16'b0000_0000_0000_0000;
array[63598] <= 16'b0000_0000_0000_0000;
array[63599] <= 16'b0000_0000_0000_0000;
array[63600] <= 16'b0000_0000_0000_0000;
array[63601] <= 16'b0000_0000_0000_0000;
array[63602] <= 16'b0000_0000_0000_0000;
array[63603] <= 16'b0000_0000_0000_0000;
array[63604] <= 16'b0000_0000_0000_0000;
array[63605] <= 16'b0000_0000_0000_0000;
array[63606] <= 16'b0000_0000_0000_0000;
array[63607] <= 16'b0000_0000_0000_0000;
array[63608] <= 16'b0000_0000_0000_0000;
array[63609] <= 16'b0000_0000_0000_0000;
array[63610] <= 16'b0000_0000_0000_0000;
array[63611] <= 16'b0000_0000_0000_0000;
array[63612] <= 16'b0000_0000_0000_0000;
array[63613] <= 16'b0000_0000_0000_0000;
array[63614] <= 16'b0000_0000_0000_0000;
array[63615] <= 16'b0000_0000_0000_0000;
array[63616] <= 16'b0000_0000_0000_0000;
array[63617] <= 16'b0000_0000_0000_0000;
array[63618] <= 16'b0000_0000_0000_0000;
array[63619] <= 16'b0000_0000_0000_0000;
array[63620] <= 16'b0000_0000_0000_0000;
array[63621] <= 16'b0000_0000_0000_0000;
array[63622] <= 16'b0000_0000_0000_0000;
array[63623] <= 16'b0000_0000_0000_0000;
array[63624] <= 16'b0000_0000_0000_0000;
array[63625] <= 16'b0000_0000_0000_0000;
array[63626] <= 16'b0000_0000_0000_0000;
array[63627] <= 16'b0000_0000_0000_0000;
array[63628] <= 16'b0000_0000_0000_0000;
array[63629] <= 16'b0000_0000_0000_0000;
array[63630] <= 16'b0000_0000_0000_0000;
array[63631] <= 16'b0000_0000_0000_0000;
array[63632] <= 16'b0000_0000_0000_0000;
array[63633] <= 16'b0000_0000_0000_0000;
array[63634] <= 16'b0000_0000_0000_0000;
array[63635] <= 16'b0000_0000_0000_0000;
array[63636] <= 16'b0000_0000_0000_0000;
array[63637] <= 16'b0000_0000_0000_0000;
array[63638] <= 16'b0000_0000_0000_0000;
array[63639] <= 16'b0000_0000_0000_0000;
array[63640] <= 16'b0000_0000_0000_0000;
array[63641] <= 16'b0000_0000_0000_0000;
array[63642] <= 16'b0000_0000_0000_0000;
array[63643] <= 16'b0000_0000_0000_0000;
array[63644] <= 16'b0000_0000_0000_0000;
array[63645] <= 16'b0000_0000_0000_0000;
array[63646] <= 16'b0000_0000_0000_0000;
array[63647] <= 16'b0000_0000_0000_0000;
array[63648] <= 16'b0000_0000_0000_0000;
array[63649] <= 16'b0000_0000_0000_0000;
array[63650] <= 16'b0000_0000_0000_0000;
array[63651] <= 16'b0000_0000_0000_0000;
array[63652] <= 16'b0000_0000_0000_0000;
array[63653] <= 16'b0000_0000_0000_0000;
array[63654] <= 16'b0000_0000_0000_0000;
array[63655] <= 16'b0000_0000_0000_0000;
array[63656] <= 16'b0000_0000_0000_0000;
array[63657] <= 16'b0000_0000_0000_0000;
array[63658] <= 16'b0000_0000_0000_0000;
array[63659] <= 16'b0000_0000_0000_0000;
array[63660] <= 16'b0000_0000_0000_0000;
array[63661] <= 16'b0000_0000_0000_0000;
array[63662] <= 16'b0000_0000_0000_0000;
array[63663] <= 16'b0000_0000_0000_0000;
array[63664] <= 16'b0000_0000_0000_0000;
array[63665] <= 16'b0000_0000_0000_0000;
array[63666] <= 16'b0000_0000_0000_0000;
array[63667] <= 16'b0000_0000_0000_0000;
array[63668] <= 16'b0000_0000_0000_0000;
array[63669] <= 16'b0000_0000_0000_0000;
array[63670] <= 16'b0000_0000_0000_0000;
array[63671] <= 16'b0000_0000_0000_0000;
array[63672] <= 16'b0000_0000_0000_0000;
array[63673] <= 16'b0000_0000_0000_0000;
array[63674] <= 16'b0000_0000_0000_0000;
array[63675] <= 16'b0000_0000_0000_0000;
array[63676] <= 16'b0000_0000_0000_0000;
array[63677] <= 16'b0000_0000_0000_0000;
array[63678] <= 16'b0000_0000_0000_0000;
array[63679] <= 16'b0000_0000_0000_0000;
array[63680] <= 16'b0000_0000_0000_0000;
array[63681] <= 16'b0000_0000_0000_0000;
array[63682] <= 16'b0000_0000_0000_0000;
array[63683] <= 16'b0000_0000_0000_0000;
array[63684] <= 16'b0000_0000_0000_0000;
array[63685] <= 16'b0000_0000_0000_0000;
array[63686] <= 16'b0000_0000_0000_0000;
array[63687] <= 16'b0000_0000_0000_0000;
array[63688] <= 16'b0000_0000_0000_0000;
array[63689] <= 16'b0000_0000_0000_0000;
array[63690] <= 16'b0000_0000_0000_0000;
array[63691] <= 16'b0000_0000_0000_0000;
array[63692] <= 16'b0000_0000_0000_0000;
array[63693] <= 16'b0000_0000_0000_0000;
array[63694] <= 16'b0000_0000_0000_0000;
array[63695] <= 16'b0000_0000_0000_0000;
array[63696] <= 16'b0000_0000_0000_0000;
array[63697] <= 16'b0000_0000_0000_0000;
array[63698] <= 16'b0000_0000_0000_0000;
array[63699] <= 16'b0000_0000_0000_0000;
array[63700] <= 16'b0000_0000_0000_0000;
array[63701] <= 16'b0000_0000_0000_0000;
array[63702] <= 16'b0000_0000_0000_0000;
array[63703] <= 16'b0000_0000_0000_0000;
array[63704] <= 16'b0000_0000_0000_0000;
array[63705] <= 16'b0000_0000_0000_0000;
array[63706] <= 16'b0000_0000_0000_0000;
array[63707] <= 16'b0000_0000_0000_0000;
array[63708] <= 16'b0000_0000_0000_0000;
array[63709] <= 16'b0000_0000_0000_0000;
array[63710] <= 16'b0000_0000_0000_0000;
array[63711] <= 16'b0000_0000_0000_0000;
array[63712] <= 16'b0000_0000_0000_0000;
array[63713] <= 16'b0000_0000_0000_0000;
array[63714] <= 16'b0000_0000_0000_0000;
array[63715] <= 16'b0000_0000_0000_0000;
array[63716] <= 16'b0000_0000_0000_0000;
array[63717] <= 16'b0000_0000_0000_0000;
array[63718] <= 16'b0000_0000_0000_0000;
array[63719] <= 16'b0000_0000_0000_0000;
array[63720] <= 16'b0000_0000_0000_0000;
array[63721] <= 16'b0000_0000_0000_0000;
array[63722] <= 16'b0000_0000_0000_0000;
array[63723] <= 16'b0000_0000_0000_0000;
array[63724] <= 16'b0000_0000_0000_0000;
array[63725] <= 16'b0000_0000_0000_0000;
array[63726] <= 16'b0000_0000_0000_0000;
array[63727] <= 16'b0000_0000_0000_0000;
array[63728] <= 16'b0000_0000_0000_0000;
array[63729] <= 16'b0000_0000_0000_0000;
array[63730] <= 16'b0000_0000_0000_0000;
array[63731] <= 16'b0000_0000_0000_0000;
array[63732] <= 16'b0000_0000_0000_0000;
array[63733] <= 16'b0000_0000_0000_0000;
array[63734] <= 16'b0000_0000_0000_0000;
array[63735] <= 16'b0000_0000_0000_0000;
array[63736] <= 16'b0000_0000_0000_0000;
array[63737] <= 16'b0000_0000_0000_0000;
array[63738] <= 16'b0000_0000_0000_0000;
array[63739] <= 16'b0000_0000_0000_0000;
array[63740] <= 16'b0000_0000_0000_0000;
array[63741] <= 16'b0000_0000_0000_0000;
array[63742] <= 16'b0000_0000_0000_0000;
array[63743] <= 16'b0000_0000_0000_0000;
array[63744] <= 16'b0000_0000_0000_0000;
array[63745] <= 16'b0000_0000_0000_0000;
array[63746] <= 16'b0000_0000_0000_0000;
array[63747] <= 16'b0000_0000_0000_0000;
array[63748] <= 16'b0000_0000_0000_0000;
array[63749] <= 16'b0000_0000_0000_0000;
array[63750] <= 16'b0000_0000_0000_0000;
array[63751] <= 16'b0000_0000_0000_0000;
array[63752] <= 16'b0000_0000_0000_0000;
array[63753] <= 16'b0000_0000_0000_0000;
array[63754] <= 16'b0000_0000_0000_0000;
array[63755] <= 16'b0000_0000_0000_0000;
array[63756] <= 16'b0000_0000_0000_0000;
array[63757] <= 16'b0000_0000_0000_0000;
array[63758] <= 16'b0000_0000_0000_0000;
array[63759] <= 16'b0000_0000_0000_0000;
array[63760] <= 16'b0000_0000_0000_0000;
array[63761] <= 16'b0000_0000_0000_0000;
array[63762] <= 16'b0000_0000_0000_0000;
array[63763] <= 16'b0000_0000_0000_0000;
array[63764] <= 16'b0000_0000_0000_0000;
array[63765] <= 16'b0000_0000_0000_0000;
array[63766] <= 16'b0000_0000_0000_0000;
array[63767] <= 16'b0000_0000_0000_0000;
array[63768] <= 16'b0000_0000_0000_0000;
array[63769] <= 16'b0000_0000_0000_0000;
array[63770] <= 16'b0000_0000_0000_0000;
array[63771] <= 16'b0000_0000_0000_0000;
array[63772] <= 16'b0000_0000_0000_0000;
array[63773] <= 16'b0000_0000_0000_0000;
array[63774] <= 16'b0000_0000_0000_0000;
array[63775] <= 16'b0000_0000_0000_0000;
array[63776] <= 16'b0000_0000_0000_0000;
array[63777] <= 16'b0000_0000_0000_0000;
array[63778] <= 16'b0000_0000_0000_0000;
array[63779] <= 16'b0000_0000_0000_0000;
array[63780] <= 16'b0000_0000_0000_0000;
array[63781] <= 16'b0000_0000_0000_0000;
array[63782] <= 16'b0000_0000_0000_0000;
array[63783] <= 16'b0000_0000_0000_0000;
array[63784] <= 16'b0000_0000_0000_0000;
array[63785] <= 16'b0000_0000_0000_0000;
array[63786] <= 16'b0000_0000_0000_0000;
array[63787] <= 16'b0000_0000_0000_0000;
array[63788] <= 16'b0000_0000_0000_0000;
array[63789] <= 16'b0000_0000_0000_0000;
array[63790] <= 16'b0000_0000_0000_0000;
array[63791] <= 16'b0000_0000_0000_0000;
array[63792] <= 16'b0000_0000_0000_0000;
array[63793] <= 16'b0000_0000_0000_0000;
array[63794] <= 16'b0000_0000_0000_0000;
array[63795] <= 16'b0000_0000_0000_0000;
array[63796] <= 16'b0000_0000_0000_0000;
array[63797] <= 16'b0000_0000_0000_0000;
array[63798] <= 16'b0000_0000_0000_0000;
array[63799] <= 16'b0000_0000_0000_0000;
array[63800] <= 16'b0000_0000_0000_0000;
array[63801] <= 16'b0000_0000_0000_0000;
array[63802] <= 16'b0000_0000_0000_0000;
array[63803] <= 16'b0000_0000_0000_0000;
array[63804] <= 16'b0000_0000_0000_0000;
array[63805] <= 16'b0000_0000_0000_0000;
array[63806] <= 16'b0000_0000_0000_0000;
array[63807] <= 16'b0000_0000_0000_0000;
array[63808] <= 16'b0000_0000_0000_0000;
array[63809] <= 16'b0000_0000_0000_0000;
array[63810] <= 16'b0000_0000_0000_0000;
array[63811] <= 16'b0000_0000_0000_0000;
array[63812] <= 16'b0000_0000_0000_0000;
array[63813] <= 16'b0000_0000_0000_0000;
array[63814] <= 16'b0000_0000_0000_0000;
array[63815] <= 16'b0000_0000_0000_0000;
array[63816] <= 16'b0000_0000_0000_0000;
array[63817] <= 16'b0000_0000_0000_0000;
array[63818] <= 16'b0000_0000_0000_0000;
array[63819] <= 16'b0000_0000_0000_0000;
array[63820] <= 16'b0000_0000_0000_0000;
array[63821] <= 16'b0000_0000_0000_0000;
array[63822] <= 16'b0000_0000_0000_0000;
array[63823] <= 16'b0000_0000_0000_0000;
array[63824] <= 16'b0000_0000_0000_0000;
array[63825] <= 16'b0000_0000_0000_0000;
array[63826] <= 16'b0000_0000_0000_0000;
array[63827] <= 16'b0000_0000_0000_0000;
array[63828] <= 16'b0000_0000_0000_0000;
array[63829] <= 16'b0000_0000_0000_0000;
array[63830] <= 16'b0000_0000_0000_0000;
array[63831] <= 16'b0000_0000_0000_0000;
array[63832] <= 16'b0000_0000_0000_0000;
array[63833] <= 16'b0000_0000_0000_0000;
array[63834] <= 16'b0000_0000_0000_0000;
array[63835] <= 16'b0000_0000_0000_0000;
array[63836] <= 16'b0000_0000_0000_0000;
array[63837] <= 16'b0000_0000_0000_0000;
array[63838] <= 16'b0000_0000_0000_0000;
array[63839] <= 16'b0000_0000_0000_0000;
array[63840] <= 16'b0000_0000_0000_0000;
array[63841] <= 16'b0000_0000_0000_0000;
array[63842] <= 16'b0000_0000_0000_0000;
array[63843] <= 16'b0000_0000_0000_0000;
array[63844] <= 16'b0000_0000_0000_0000;
array[63845] <= 16'b0000_0000_0000_0000;
array[63846] <= 16'b0000_0000_0000_0000;
array[63847] <= 16'b0000_0000_0000_0000;
array[63848] <= 16'b0000_0000_0000_0000;
array[63849] <= 16'b0000_0000_0000_0000;
array[63850] <= 16'b0000_0000_0000_0000;
array[63851] <= 16'b0000_0000_0000_0000;
array[63852] <= 16'b0000_0000_0000_0000;
array[63853] <= 16'b0000_0000_0000_0000;
array[63854] <= 16'b0000_0000_0000_0000;
array[63855] <= 16'b0000_0000_0000_0000;
array[63856] <= 16'b0000_0000_0000_0000;
array[63857] <= 16'b0000_0000_0000_0000;
array[63858] <= 16'b0000_0000_0000_0000;
array[63859] <= 16'b0000_0000_0000_0000;
array[63860] <= 16'b0000_0000_0000_0000;
array[63861] <= 16'b0000_0000_0000_0000;
array[63862] <= 16'b0000_0000_0000_0000;
array[63863] <= 16'b0000_0000_0000_0000;
array[63864] <= 16'b0000_0000_0000_0000;
array[63865] <= 16'b0000_0000_0000_0000;
array[63866] <= 16'b0000_0000_0000_0000;
array[63867] <= 16'b0000_0000_0000_0000;
array[63868] <= 16'b0000_0000_0000_0000;
array[63869] <= 16'b0000_0000_0000_0000;
array[63870] <= 16'b0000_0000_0000_0000;
array[63871] <= 16'b0000_0000_0000_0000;
array[63872] <= 16'b0000_0000_0000_0000;
array[63873] <= 16'b0000_0000_0000_0000;
array[63874] <= 16'b0000_0000_0000_0000;
array[63875] <= 16'b0000_0000_0000_0000;
array[63876] <= 16'b0000_0000_0000_0000;
array[63877] <= 16'b0000_0000_0000_0000;
array[63878] <= 16'b0000_0000_0000_0000;
array[63879] <= 16'b0000_0000_0000_0000;
array[63880] <= 16'b0000_0000_0000_0000;
array[63881] <= 16'b0000_0000_0000_0000;
array[63882] <= 16'b0000_0000_0000_0000;
array[63883] <= 16'b0000_0000_0000_0000;
array[63884] <= 16'b0000_0000_0000_0000;
array[63885] <= 16'b0000_0000_0000_0000;
array[63886] <= 16'b0000_0000_0000_0000;
array[63887] <= 16'b0000_0000_0000_0000;
array[63888] <= 16'b0000_0000_0000_0000;
array[63889] <= 16'b0000_0000_0000_0000;
array[63890] <= 16'b0000_0000_0000_0000;
array[63891] <= 16'b0000_0000_0000_0000;
array[63892] <= 16'b0000_0000_0000_0000;
array[63893] <= 16'b0000_0000_0000_0000;
array[63894] <= 16'b0000_0000_0000_0000;
array[63895] <= 16'b0000_0000_0000_0000;
array[63896] <= 16'b0000_0000_0000_0000;
array[63897] <= 16'b0000_0000_0000_0000;
array[63898] <= 16'b0000_0000_0000_0000;
array[63899] <= 16'b0000_0000_0000_0000;
array[63900] <= 16'b0000_0000_0000_0000;
array[63901] <= 16'b0000_0000_0000_0000;
array[63902] <= 16'b0000_0000_0000_0000;
array[63903] <= 16'b0000_0000_0000_0000;
array[63904] <= 16'b0000_0000_0000_0000;
array[63905] <= 16'b0000_0000_0000_0000;
array[63906] <= 16'b0000_0000_0000_0000;
array[63907] <= 16'b0000_0000_0000_0000;
array[63908] <= 16'b0000_0000_0000_0000;
array[63909] <= 16'b0000_0000_0000_0000;
array[63910] <= 16'b0000_0000_0000_0000;
array[63911] <= 16'b0000_0000_0000_0000;
array[63912] <= 16'b0000_0000_0000_0000;
array[63913] <= 16'b0000_0000_0000_0000;
array[63914] <= 16'b0000_0000_0000_0000;
array[63915] <= 16'b0000_0000_0000_0000;
array[63916] <= 16'b0000_0000_0000_0000;
array[63917] <= 16'b0000_0000_0000_0000;
array[63918] <= 16'b0000_0000_0000_0000;
array[63919] <= 16'b0000_0000_0000_0000;
array[63920] <= 16'b0000_0000_0000_0000;
array[63921] <= 16'b0000_0000_0000_0000;
array[63922] <= 16'b0000_0000_0000_0000;
array[63923] <= 16'b0000_0000_0000_0000;
array[63924] <= 16'b0000_0000_0000_0000;
array[63925] <= 16'b0000_0000_0000_0000;
array[63926] <= 16'b0000_0000_0000_0000;
array[63927] <= 16'b0000_0000_0000_0000;
array[63928] <= 16'b0000_0000_0000_0000;
array[63929] <= 16'b0000_0000_0000_0000;
array[63930] <= 16'b0000_0000_0000_0000;
array[63931] <= 16'b0000_0000_0000_0000;
array[63932] <= 16'b0000_0000_0000_0000;
array[63933] <= 16'b0000_0000_0000_0000;
array[63934] <= 16'b0000_0000_0000_0000;
array[63935] <= 16'b0000_0000_0000_0000;
array[63936] <= 16'b0000_0000_0000_0000;
array[63937] <= 16'b0000_0000_0000_0000;
array[63938] <= 16'b0000_0000_0000_0000;
array[63939] <= 16'b0000_0000_0000_0000;
array[63940] <= 16'b0000_0000_0000_0000;
array[63941] <= 16'b0000_0000_0000_0000;
array[63942] <= 16'b0000_0000_0000_0000;
array[63943] <= 16'b0000_0000_0000_0000;
array[63944] <= 16'b0000_0000_0000_0000;
array[63945] <= 16'b0000_0000_0000_0000;
array[63946] <= 16'b0000_0000_0000_0000;
array[63947] <= 16'b0000_0000_0000_0000;
array[63948] <= 16'b0000_0000_0000_0000;
array[63949] <= 16'b0000_0000_0000_0000;
array[63950] <= 16'b0000_0000_0000_0000;
array[63951] <= 16'b0000_0000_0000_0000;
array[63952] <= 16'b0000_0000_0000_0000;
array[63953] <= 16'b0000_0000_0000_0000;
array[63954] <= 16'b0000_0000_0000_0000;
array[63955] <= 16'b0000_0000_0000_0000;
array[63956] <= 16'b0000_0000_0000_0000;
array[63957] <= 16'b0000_0000_0000_0000;
array[63958] <= 16'b0000_0000_0000_0000;
array[63959] <= 16'b0000_0000_0000_0000;
array[63960] <= 16'b0000_0000_0000_0000;
array[63961] <= 16'b0000_0000_0000_0000;
array[63962] <= 16'b0000_0000_0000_0000;
array[63963] <= 16'b0000_0000_0000_0000;
array[63964] <= 16'b0000_0000_0000_0000;
array[63965] <= 16'b0000_0000_0000_0000;
array[63966] <= 16'b0000_0000_0000_0000;
array[63967] <= 16'b0000_0000_0000_0000;
array[63968] <= 16'b0000_0000_0000_0000;
array[63969] <= 16'b0000_0000_0000_0000;
array[63970] <= 16'b0000_0000_0000_0000;
array[63971] <= 16'b0000_0000_0000_0000;
array[63972] <= 16'b0000_0000_0000_0000;
array[63973] <= 16'b0000_0000_0000_0000;
array[63974] <= 16'b0000_0000_0000_0000;
array[63975] <= 16'b0000_0000_0000_0000;
array[63976] <= 16'b0000_0000_0000_0000;
array[63977] <= 16'b0000_0000_0000_0000;
array[63978] <= 16'b0000_0000_0000_0000;
array[63979] <= 16'b0000_0000_0000_0000;
array[63980] <= 16'b0000_0000_0000_0000;
array[63981] <= 16'b0000_0000_0000_0000;
array[63982] <= 16'b0000_0000_0000_0000;
array[63983] <= 16'b0000_0000_0000_0000;
array[63984] <= 16'b0000_0000_0000_0000;
array[63985] <= 16'b0000_0000_0000_0000;
array[63986] <= 16'b0000_0000_0000_0000;
array[63987] <= 16'b0000_0000_0000_0000;
array[63988] <= 16'b0000_0000_0000_0000;
array[63989] <= 16'b0000_0000_0000_0000;
array[63990] <= 16'b0000_0000_0000_0000;
array[63991] <= 16'b0000_0000_0000_0000;
array[63992] <= 16'b0000_0000_0000_0000;
array[63993] <= 16'b0000_0000_0000_0000;
array[63994] <= 16'b0000_0000_0000_0000;
array[63995] <= 16'b0000_0000_0000_0000;
array[63996] <= 16'b0000_0000_0000_0000;
array[63997] <= 16'b0000_0000_0000_0000;
array[63998] <= 16'b0000_0000_0000_0000;
array[63999] <= 16'b0000_0000_0000_0000;
array[64000] <= 16'b0000_0000_0000_0000;
array[64001] <= 16'b0000_0000_0000_0000;
array[64002] <= 16'b0000_0000_0000_0000;
array[64003] <= 16'b0000_0000_0000_0000;
array[64004] <= 16'b0000_0000_0000_0000;
array[64005] <= 16'b0000_0000_0000_0000;
array[64006] <= 16'b0000_0000_0000_0000;
array[64007] <= 16'b0000_0000_0000_0000;
array[64008] <= 16'b0000_0000_0000_0000;
array[64009] <= 16'b0000_0000_0000_0000;
array[64010] <= 16'b0000_0000_0000_0000;
array[64011] <= 16'b0000_0000_0000_0000;
array[64012] <= 16'b0000_0000_0000_0000;
array[64013] <= 16'b0000_0000_0000_0000;
array[64014] <= 16'b0000_0000_0000_0000;
array[64015] <= 16'b0000_0000_0000_0000;
array[64016] <= 16'b0000_0000_0000_0000;
array[64017] <= 16'b0000_0000_0000_0000;
array[64018] <= 16'b0000_0000_0000_0000;
array[64019] <= 16'b0000_0000_0000_0000;
array[64020] <= 16'b0000_0000_0000_0000;
array[64021] <= 16'b0000_0000_0000_0000;
array[64022] <= 16'b0000_0000_0000_0000;
array[64023] <= 16'b0000_0000_0000_0000;
array[64024] <= 16'b0000_0000_0000_0000;
array[64025] <= 16'b0000_0000_0000_0000;
array[64026] <= 16'b0000_0000_0000_0000;
array[64027] <= 16'b0000_0000_0000_0000;
array[64028] <= 16'b0000_0000_0000_0000;
array[64029] <= 16'b0000_0000_0000_0000;
array[64030] <= 16'b0000_0000_0000_0000;
array[64031] <= 16'b0000_0000_0000_0000;
array[64032] <= 16'b0000_0000_0000_0000;
array[64033] <= 16'b0000_0000_0000_0000;
array[64034] <= 16'b0000_0000_0000_0000;
array[64035] <= 16'b0000_0000_0000_0000;
array[64036] <= 16'b0000_0000_0000_0000;
array[64037] <= 16'b0000_0000_0000_0000;
array[64038] <= 16'b0000_0000_0000_0000;
array[64039] <= 16'b0000_0000_0000_0000;
array[64040] <= 16'b0000_0000_0000_0000;
array[64041] <= 16'b0000_0000_0000_0000;
array[64042] <= 16'b0000_0000_0000_0000;
array[64043] <= 16'b0000_0000_0000_0000;
array[64044] <= 16'b0000_0000_0000_0000;
array[64045] <= 16'b0000_0000_0000_0000;
array[64046] <= 16'b0000_0000_0000_0000;
array[64047] <= 16'b0000_0000_0000_0000;
array[64048] <= 16'b0000_0000_0000_0000;
array[64049] <= 16'b0000_0000_0000_0000;
array[64050] <= 16'b0000_0000_0000_0000;
array[64051] <= 16'b0000_0000_0000_0000;
array[64052] <= 16'b0000_0000_0000_0000;
array[64053] <= 16'b0000_0000_0000_0000;
array[64054] <= 16'b0000_0000_0000_0000;
array[64055] <= 16'b0000_0000_0000_0000;
array[64056] <= 16'b0000_0000_0000_0000;
array[64057] <= 16'b0000_0000_0000_0000;
array[64058] <= 16'b0000_0000_0000_0000;
array[64059] <= 16'b0000_0000_0000_0000;
array[64060] <= 16'b0000_0000_0000_0000;
array[64061] <= 16'b0000_0000_0000_0000;
array[64062] <= 16'b0000_0000_0000_0000;
array[64063] <= 16'b0000_0000_0000_0000;
array[64064] <= 16'b0000_0000_0000_0000;
array[64065] <= 16'b0000_0000_0000_0000;
array[64066] <= 16'b0000_0000_0000_0000;
array[64067] <= 16'b0000_0000_0000_0000;
array[64068] <= 16'b0000_0000_0000_0000;
array[64069] <= 16'b0000_0000_0000_0000;
array[64070] <= 16'b0000_0000_0000_0000;
array[64071] <= 16'b0000_0000_0000_0000;
array[64072] <= 16'b0000_0000_0000_0000;
array[64073] <= 16'b0000_0000_0000_0000;
array[64074] <= 16'b0000_0000_0000_0000;
array[64075] <= 16'b0000_0000_0000_0000;
array[64076] <= 16'b0000_0000_0000_0000;
array[64077] <= 16'b0000_0000_0000_0000;
array[64078] <= 16'b0000_0000_0000_0000;
array[64079] <= 16'b0000_0000_0000_0000;
array[64080] <= 16'b0000_0000_0000_0000;
array[64081] <= 16'b0000_0000_0000_0000;
array[64082] <= 16'b0000_0000_0000_0000;
array[64083] <= 16'b0000_0000_0000_0000;
array[64084] <= 16'b0000_0000_0000_0000;
array[64085] <= 16'b0000_0000_0000_0000;
array[64086] <= 16'b0000_0000_0000_0000;
array[64087] <= 16'b0000_0000_0000_0000;
array[64088] <= 16'b0000_0000_0000_0000;
array[64089] <= 16'b0000_0000_0000_0000;
array[64090] <= 16'b0000_0000_0000_0000;
array[64091] <= 16'b0000_0000_0000_0000;
array[64092] <= 16'b0000_0000_0000_0000;
array[64093] <= 16'b0000_0000_0000_0000;
array[64094] <= 16'b0000_0000_0000_0000;
array[64095] <= 16'b0000_0000_0000_0000;
array[64096] <= 16'b0000_0000_0000_0000;
array[64097] <= 16'b0000_0000_0000_0000;
array[64098] <= 16'b0000_0000_0000_0000;
array[64099] <= 16'b0000_0000_0000_0000;
array[64100] <= 16'b0000_0000_0000_0000;
array[64101] <= 16'b0000_0000_0000_0000;
array[64102] <= 16'b0000_0000_0000_0000;
array[64103] <= 16'b0000_0000_0000_0000;
array[64104] <= 16'b0000_0000_0000_0000;
array[64105] <= 16'b0000_0000_0000_0000;
array[64106] <= 16'b0000_0000_0000_0000;
array[64107] <= 16'b0000_0000_0000_0000;
array[64108] <= 16'b0000_0000_0000_0000;
array[64109] <= 16'b0000_0000_0000_0000;
array[64110] <= 16'b0000_0000_0000_0000;
array[64111] <= 16'b0000_0000_0000_0000;
array[64112] <= 16'b0000_0000_0000_0000;
array[64113] <= 16'b0000_0000_0000_0000;
array[64114] <= 16'b0000_0000_0000_0000;
array[64115] <= 16'b0000_0000_0000_0000;
array[64116] <= 16'b0000_0000_0000_0000;
array[64117] <= 16'b0000_0000_0000_0000;
array[64118] <= 16'b0000_0000_0000_0000;
array[64119] <= 16'b0000_0000_0000_0000;
array[64120] <= 16'b0000_0000_0000_0000;
array[64121] <= 16'b0000_0000_0000_0000;
array[64122] <= 16'b0000_0000_0000_0000;
array[64123] <= 16'b0000_0000_0000_0000;
array[64124] <= 16'b0000_0000_0000_0000;
array[64125] <= 16'b0000_0000_0000_0000;
array[64126] <= 16'b0000_0000_0000_0000;
array[64127] <= 16'b0000_0000_0000_0000;
array[64128] <= 16'b0000_0000_0000_0000;
array[64129] <= 16'b0000_0000_0000_0000;
array[64130] <= 16'b0000_0000_0000_0000;
array[64131] <= 16'b0000_0000_0000_0000;
array[64132] <= 16'b0000_0000_0000_0000;
array[64133] <= 16'b0000_0000_0000_0000;
array[64134] <= 16'b0000_0000_0000_0000;
array[64135] <= 16'b0000_0000_0000_0000;
array[64136] <= 16'b0000_0000_0000_0000;
array[64137] <= 16'b0000_0000_0000_0000;
array[64138] <= 16'b0000_0000_0000_0000;
array[64139] <= 16'b0000_0000_0000_0000;
array[64140] <= 16'b0000_0000_0000_0000;
array[64141] <= 16'b0000_0000_0000_0000;
array[64142] <= 16'b0000_0000_0000_0000;
array[64143] <= 16'b0000_0000_0000_0000;
array[64144] <= 16'b0000_0000_0000_0000;
array[64145] <= 16'b0000_0000_0000_0000;
array[64146] <= 16'b0000_0000_0000_0000;
array[64147] <= 16'b0000_0000_0000_0000;
array[64148] <= 16'b0000_0000_0000_0000;
array[64149] <= 16'b0000_0000_0000_0000;
array[64150] <= 16'b0000_0000_0000_0000;
array[64151] <= 16'b0000_0000_0000_0000;
array[64152] <= 16'b0000_0000_0000_0000;
array[64153] <= 16'b0000_0000_0000_0000;
array[64154] <= 16'b0000_0000_0000_0000;
array[64155] <= 16'b0000_0000_0000_0000;
array[64156] <= 16'b0000_0000_0000_0000;
array[64157] <= 16'b0000_0000_0000_0000;
array[64158] <= 16'b0000_0000_0000_0000;
array[64159] <= 16'b0000_0000_0000_0000;
array[64160] <= 16'b0000_0000_0000_0000;
array[64161] <= 16'b0000_0000_0000_0000;
array[64162] <= 16'b0000_0000_0000_0000;
array[64163] <= 16'b0000_0000_0000_0000;
array[64164] <= 16'b0000_0000_0000_0000;
array[64165] <= 16'b0000_0000_0000_0000;
array[64166] <= 16'b0000_0000_0000_0000;
array[64167] <= 16'b0000_0000_0000_0000;
array[64168] <= 16'b0000_0000_0000_0000;
array[64169] <= 16'b0000_0000_0000_0000;
array[64170] <= 16'b0000_0000_0000_0000;
array[64171] <= 16'b0000_0000_0000_0000;
array[64172] <= 16'b0000_0000_0000_0000;
array[64173] <= 16'b0000_0000_0000_0000;
array[64174] <= 16'b0000_0000_0000_0000;
array[64175] <= 16'b0000_0000_0000_0000;
array[64176] <= 16'b0000_0000_0000_0000;
array[64177] <= 16'b0000_0000_0000_0000;
array[64178] <= 16'b0000_0000_0000_0000;
array[64179] <= 16'b0000_0000_0000_0000;
array[64180] <= 16'b0000_0000_0000_0000;
array[64181] <= 16'b0000_0000_0000_0000;
array[64182] <= 16'b0000_0000_0000_0000;
array[64183] <= 16'b0000_0000_0000_0000;
array[64184] <= 16'b0000_0000_0000_0000;
array[64185] <= 16'b0000_0000_0000_0000;
array[64186] <= 16'b0000_0000_0000_0000;
array[64187] <= 16'b0000_0000_0000_0000;
array[64188] <= 16'b0000_0000_0000_0000;
array[64189] <= 16'b0000_0000_0000_0000;
array[64190] <= 16'b0000_0000_0000_0000;
array[64191] <= 16'b0000_0000_0000_0000;
array[64192] <= 16'b0000_0000_0000_0000;
array[64193] <= 16'b0000_0000_0000_0000;
array[64194] <= 16'b0000_0000_0000_0000;
array[64195] <= 16'b0000_0000_0000_0000;
array[64196] <= 16'b0000_0000_0000_0000;
array[64197] <= 16'b0000_0000_0000_0000;
array[64198] <= 16'b0000_0000_0000_0000;
array[64199] <= 16'b0000_0000_0000_0000;
array[64200] <= 16'b0000_0000_0000_0000;
array[64201] <= 16'b0000_0000_0000_0000;
array[64202] <= 16'b0000_0000_0000_0000;
array[64203] <= 16'b0000_0000_0000_0000;
array[64204] <= 16'b0000_0000_0000_0000;
array[64205] <= 16'b0000_0000_0000_0000;
array[64206] <= 16'b0000_0000_0000_0000;
array[64207] <= 16'b0000_0000_0000_0000;
array[64208] <= 16'b0000_0000_0000_0000;
array[64209] <= 16'b0000_0000_0000_0000;
array[64210] <= 16'b0000_0000_0000_0000;
array[64211] <= 16'b0000_0000_0000_0000;
array[64212] <= 16'b0000_0000_0000_0000;
array[64213] <= 16'b0000_0000_0000_0000;
array[64214] <= 16'b0000_0000_0000_0000;
array[64215] <= 16'b0000_0000_0000_0000;
array[64216] <= 16'b0000_0000_0000_0000;
array[64217] <= 16'b0000_0000_0000_0000;
array[64218] <= 16'b0000_0000_0000_0000;
array[64219] <= 16'b0000_0000_0000_0000;
array[64220] <= 16'b0000_0000_0000_0000;
array[64221] <= 16'b0000_0000_0000_0000;
array[64222] <= 16'b0000_0000_0000_0000;
array[64223] <= 16'b0000_0000_0000_0000;
array[64224] <= 16'b0000_0000_0000_0000;
array[64225] <= 16'b0000_0000_0000_0000;
array[64226] <= 16'b0000_0000_0000_0000;
array[64227] <= 16'b0000_0000_0000_0000;
array[64228] <= 16'b0000_0000_0000_0000;
array[64229] <= 16'b0000_0000_0000_0000;
array[64230] <= 16'b0000_0000_0000_0000;
array[64231] <= 16'b0000_0000_0000_0000;
array[64232] <= 16'b0000_0000_0000_0000;
array[64233] <= 16'b0000_0000_0000_0000;
array[64234] <= 16'b0000_0000_0000_0000;
array[64235] <= 16'b0000_0000_0000_0000;
array[64236] <= 16'b0000_0000_0000_0000;
array[64237] <= 16'b0000_0000_0000_0000;
array[64238] <= 16'b0000_0000_0000_0000;
array[64239] <= 16'b0000_0000_0000_0000;
array[64240] <= 16'b0000_0000_0000_0000;
array[64241] <= 16'b0000_0000_0000_0000;
array[64242] <= 16'b0000_0000_0000_0000;
array[64243] <= 16'b0000_0000_0000_0000;
array[64244] <= 16'b0000_0000_0000_0000;
array[64245] <= 16'b0000_0000_0000_0000;
array[64246] <= 16'b0000_0000_0000_0000;
array[64247] <= 16'b0000_0000_0000_0000;
array[64248] <= 16'b0000_0000_0000_0000;
array[64249] <= 16'b0000_0000_0000_0000;
array[64250] <= 16'b0000_0000_0000_0000;
array[64251] <= 16'b0000_0000_0000_0000;
array[64252] <= 16'b0000_0000_0000_0000;
array[64253] <= 16'b0000_0000_0000_0000;
array[64254] <= 16'b0000_0000_0000_0000;
array[64255] <= 16'b0000_0000_0000_0000;
array[64256] <= 16'b0000_0000_0000_0000;
array[64257] <= 16'b0000_0000_0000_0000;
array[64258] <= 16'b0000_0000_0000_0000;
array[64259] <= 16'b0000_0000_0000_0000;
array[64260] <= 16'b0000_0000_0000_0000;
array[64261] <= 16'b0000_0000_0000_0000;
array[64262] <= 16'b0000_0000_0000_0000;
array[64263] <= 16'b0000_0000_0000_0000;
array[64264] <= 16'b0000_0000_0000_0000;
array[64265] <= 16'b0000_0000_0000_0000;
array[64266] <= 16'b0000_0000_0000_0000;
array[64267] <= 16'b0000_0000_0000_0000;
array[64268] <= 16'b0000_0000_0000_0000;
array[64269] <= 16'b0000_0000_0000_0000;
array[64270] <= 16'b0000_0000_0000_0000;
array[64271] <= 16'b0000_0000_0000_0000;
array[64272] <= 16'b0000_0000_0000_0000;
array[64273] <= 16'b0000_0000_0000_0000;
array[64274] <= 16'b0000_0000_0000_0000;
array[64275] <= 16'b0000_0000_0000_0000;
array[64276] <= 16'b0000_0000_0000_0000;
array[64277] <= 16'b0000_0000_0000_0000;
array[64278] <= 16'b0000_0000_0000_0000;
array[64279] <= 16'b0000_0000_0000_0000;
array[64280] <= 16'b0000_0000_0000_0000;
array[64281] <= 16'b0000_0000_0000_0000;
array[64282] <= 16'b0000_0000_0000_0000;
array[64283] <= 16'b0000_0000_0000_0000;
array[64284] <= 16'b0000_0000_0000_0000;
array[64285] <= 16'b0000_0000_0000_0000;
array[64286] <= 16'b0000_0000_0000_0000;
array[64287] <= 16'b0000_0000_0000_0000;
array[64288] <= 16'b0000_0000_0000_0000;
array[64289] <= 16'b0000_0000_0000_0000;
array[64290] <= 16'b0000_0000_0000_0000;
array[64291] <= 16'b0000_0000_0000_0000;
array[64292] <= 16'b0000_0000_0000_0000;
array[64293] <= 16'b0000_0000_0000_0000;
array[64294] <= 16'b0000_0000_0000_0000;
array[64295] <= 16'b0000_0000_0000_0000;
array[64296] <= 16'b0000_0000_0000_0000;
array[64297] <= 16'b0000_0000_0000_0000;
array[64298] <= 16'b0000_0000_0000_0000;
array[64299] <= 16'b0000_0000_0000_0000;
array[64300] <= 16'b0000_0000_0000_0000;
array[64301] <= 16'b0000_0000_0000_0000;
array[64302] <= 16'b0000_0000_0000_0000;
array[64303] <= 16'b0000_0000_0000_0000;
array[64304] <= 16'b0000_0000_0000_0000;
array[64305] <= 16'b0000_0000_0000_0000;
array[64306] <= 16'b0000_0000_0000_0000;
array[64307] <= 16'b0000_0000_0000_0000;
array[64308] <= 16'b0000_0000_0000_0000;
array[64309] <= 16'b0000_0000_0000_0000;
array[64310] <= 16'b0000_0000_0000_0000;
array[64311] <= 16'b0000_0000_0000_0000;
array[64312] <= 16'b0000_0000_0000_0000;
array[64313] <= 16'b0000_0000_0000_0000;
array[64314] <= 16'b0000_0000_0000_0000;
array[64315] <= 16'b0000_0000_0000_0000;
array[64316] <= 16'b0000_0000_0000_0000;
array[64317] <= 16'b0000_0000_0000_0000;
array[64318] <= 16'b0000_0000_0000_0000;
array[64319] <= 16'b0000_0000_0000_0000;
array[64320] <= 16'b0000_0000_0000_0000;
array[64321] <= 16'b0000_0000_0000_0000;
array[64322] <= 16'b0000_0000_0000_0000;
array[64323] <= 16'b0000_0000_0000_0000;
array[64324] <= 16'b0000_0000_0000_0000;
array[64325] <= 16'b0000_0000_0000_0000;
array[64326] <= 16'b0000_0000_0000_0000;
array[64327] <= 16'b0000_0000_0000_0000;
array[64328] <= 16'b0000_0000_0000_0000;
array[64329] <= 16'b0000_0000_0000_0000;
array[64330] <= 16'b0000_0000_0000_0000;
array[64331] <= 16'b0000_0000_0000_0000;
array[64332] <= 16'b0000_0000_0000_0000;
array[64333] <= 16'b0000_0000_0000_0000;
array[64334] <= 16'b0000_0000_0000_0000;
array[64335] <= 16'b0000_0000_0000_0000;
array[64336] <= 16'b0000_0000_0000_0000;
array[64337] <= 16'b0000_0000_0000_0000;
array[64338] <= 16'b0000_0000_0000_0000;
array[64339] <= 16'b0000_0000_0000_0000;
array[64340] <= 16'b0000_0000_0000_0000;
array[64341] <= 16'b0000_0000_0000_0000;
array[64342] <= 16'b0000_0000_0000_0000;
array[64343] <= 16'b0000_0000_0000_0000;
array[64344] <= 16'b0000_0000_0000_0000;
array[64345] <= 16'b0000_0000_0000_0000;
array[64346] <= 16'b0000_0000_0000_0000;
array[64347] <= 16'b0000_0000_0000_0000;
array[64348] <= 16'b0000_0000_0000_0000;
array[64349] <= 16'b0000_0000_0000_0000;
array[64350] <= 16'b0000_0000_0000_0000;
array[64351] <= 16'b0000_0000_0000_0000;
array[64352] <= 16'b0000_0000_0000_0000;
array[64353] <= 16'b0000_0000_0000_0000;
array[64354] <= 16'b0000_0000_0000_0000;
array[64355] <= 16'b0000_0000_0000_0000;
array[64356] <= 16'b0000_0000_0000_0000;
array[64357] <= 16'b0000_0000_0000_0000;
array[64358] <= 16'b0000_0000_0000_0000;
array[64359] <= 16'b0000_0000_0000_0000;
array[64360] <= 16'b0000_0000_0000_0000;
array[64361] <= 16'b0000_0000_0000_0000;
array[64362] <= 16'b0000_0000_0000_0000;
array[64363] <= 16'b0000_0000_0000_0000;
array[64364] <= 16'b0000_0000_0000_0000;
array[64365] <= 16'b0000_0000_0000_0000;
array[64366] <= 16'b0000_0000_0000_0000;
array[64367] <= 16'b0000_0000_0000_0000;
array[64368] <= 16'b0000_0000_0000_0000;
array[64369] <= 16'b0000_0000_0000_0000;
array[64370] <= 16'b0000_0000_0000_0000;
array[64371] <= 16'b0000_0000_0000_0000;
array[64372] <= 16'b0000_0000_0000_0000;
array[64373] <= 16'b0000_0000_0000_0000;
array[64374] <= 16'b0000_0000_0000_0000;
array[64375] <= 16'b0000_0000_0000_0000;
array[64376] <= 16'b0000_0000_0000_0000;
array[64377] <= 16'b0000_0000_0000_0000;
array[64378] <= 16'b0000_0000_0000_0000;
array[64379] <= 16'b0000_0000_0000_0000;
array[64380] <= 16'b0000_0000_0000_0000;
array[64381] <= 16'b0000_0000_0000_0000;
array[64382] <= 16'b0000_0000_0000_0000;
array[64383] <= 16'b0000_0000_0000_0000;
array[64384] <= 16'b0000_0000_0000_0000;
array[64385] <= 16'b0000_0000_0000_0000;
array[64386] <= 16'b0000_0000_0000_0000;
array[64387] <= 16'b0000_0000_0000_0000;
array[64388] <= 16'b0000_0000_0000_0000;
array[64389] <= 16'b0000_0000_0000_0000;
array[64390] <= 16'b0000_0000_0000_0000;
array[64391] <= 16'b0000_0000_0000_0000;
array[64392] <= 16'b0000_0000_0000_0000;
array[64393] <= 16'b0000_0000_0000_0000;
array[64394] <= 16'b0000_0000_0000_0000;
array[64395] <= 16'b0000_0000_0000_0000;
array[64396] <= 16'b0000_0000_0000_0000;
array[64397] <= 16'b0000_0000_0000_0000;
array[64398] <= 16'b0000_0000_0000_0000;
array[64399] <= 16'b0000_0000_0000_0000;
array[64400] <= 16'b0000_0000_0000_0000;
array[64401] <= 16'b0000_0000_0000_0000;
array[64402] <= 16'b0000_0000_0000_0000;
array[64403] <= 16'b0000_0000_0000_0000;
array[64404] <= 16'b0000_0000_0000_0000;
array[64405] <= 16'b0000_0000_0000_0000;
array[64406] <= 16'b0000_0000_0000_0000;
array[64407] <= 16'b0000_0000_0000_0000;
array[64408] <= 16'b0000_0000_0000_0000;
array[64409] <= 16'b0000_0000_0000_0000;
array[64410] <= 16'b0000_0000_0000_0000;
array[64411] <= 16'b0000_0000_0000_0000;
array[64412] <= 16'b0000_0000_0000_0000;
array[64413] <= 16'b0000_0000_0000_0000;
array[64414] <= 16'b0000_0000_0000_0000;
array[64415] <= 16'b0000_0000_0000_0000;
array[64416] <= 16'b0000_0000_0000_0000;
array[64417] <= 16'b0000_0000_0000_0000;
array[64418] <= 16'b0000_0000_0000_0000;
array[64419] <= 16'b0000_0000_0000_0000;
array[64420] <= 16'b0000_0000_0000_0000;
array[64421] <= 16'b0000_0000_0000_0000;
array[64422] <= 16'b0000_0000_0000_0000;
array[64423] <= 16'b0000_0000_0000_0000;
array[64424] <= 16'b0000_0000_0000_0000;
array[64425] <= 16'b0000_0000_0000_0000;
array[64426] <= 16'b0000_0000_0000_0000;
array[64427] <= 16'b0000_0000_0000_0000;
array[64428] <= 16'b0000_0000_0000_0000;
array[64429] <= 16'b0000_0000_0000_0000;
array[64430] <= 16'b0000_0000_0000_0000;
array[64431] <= 16'b0000_0000_0000_0000;
array[64432] <= 16'b0000_0000_0000_0000;
array[64433] <= 16'b0000_0000_0000_0000;
array[64434] <= 16'b0000_0000_0000_0000;
array[64435] <= 16'b0000_0000_0000_0000;
array[64436] <= 16'b0000_0000_0000_0000;
array[64437] <= 16'b0000_0000_0000_0000;
array[64438] <= 16'b0000_0000_0000_0000;
array[64439] <= 16'b0000_0000_0000_0000;
array[64440] <= 16'b0000_0000_0000_0000;
array[64441] <= 16'b0000_0000_0000_0000;
array[64442] <= 16'b0000_0000_0000_0000;
array[64443] <= 16'b0000_0000_0000_0000;
array[64444] <= 16'b0000_0000_0000_0000;
array[64445] <= 16'b0000_0000_0000_0000;
array[64446] <= 16'b0000_0000_0000_0000;
array[64447] <= 16'b0000_0000_0000_0000;
array[64448] <= 16'b0000_0000_0000_0000;
array[64449] <= 16'b0000_0000_0000_0000;
array[64450] <= 16'b0000_0000_0000_0000;
array[64451] <= 16'b0000_0000_0000_0000;
array[64452] <= 16'b0000_0000_0000_0000;
array[64453] <= 16'b0000_0000_0000_0000;
array[64454] <= 16'b0000_0000_0000_0000;
array[64455] <= 16'b0000_0000_0000_0000;
array[64456] <= 16'b0000_0000_0000_0000;
array[64457] <= 16'b0000_0000_0000_0000;
array[64458] <= 16'b0000_0000_0000_0000;
array[64459] <= 16'b0000_0000_0000_0000;
array[64460] <= 16'b0000_0000_0000_0000;
array[64461] <= 16'b0000_0000_0000_0000;
array[64462] <= 16'b0000_0000_0000_0000;
array[64463] <= 16'b0000_0000_0000_0000;
array[64464] <= 16'b0000_0000_0000_0000;
array[64465] <= 16'b0000_0000_0000_0000;
array[64466] <= 16'b0000_0000_0000_0000;
array[64467] <= 16'b0000_0000_0000_0000;
array[64468] <= 16'b0000_0000_0000_0000;
array[64469] <= 16'b0000_0000_0000_0000;
array[64470] <= 16'b0000_0000_0000_0000;
array[64471] <= 16'b0000_0000_0000_0000;
array[64472] <= 16'b0000_0000_0000_0000;
array[64473] <= 16'b0000_0000_0000_0000;
array[64474] <= 16'b0000_0000_0000_0000;
array[64475] <= 16'b0000_0000_0000_0000;
array[64476] <= 16'b0000_0000_0000_0000;
array[64477] <= 16'b0000_0000_0000_0000;
array[64478] <= 16'b0000_0000_0000_0000;
array[64479] <= 16'b0000_0000_0000_0000;
array[64480] <= 16'b0000_0000_0000_0000;
array[64481] <= 16'b0000_0000_0000_0000;
array[64482] <= 16'b0000_0000_0000_0000;
array[64483] <= 16'b0000_0000_0000_0000;
array[64484] <= 16'b0000_0000_0000_0000;
array[64485] <= 16'b0000_0000_0000_0000;
array[64486] <= 16'b0000_0000_0000_0000;
array[64487] <= 16'b0000_0000_0000_0000;
array[64488] <= 16'b0000_0000_0000_0000;
array[64489] <= 16'b0000_0000_0000_0000;
array[64490] <= 16'b0000_0000_0000_0000;
array[64491] <= 16'b0000_0000_0000_0000;
array[64492] <= 16'b0000_0000_0000_0000;
array[64493] <= 16'b0000_0000_0000_0000;
array[64494] <= 16'b0000_0000_0000_0000;
array[64495] <= 16'b0000_0000_0000_0000;
array[64496] <= 16'b0000_0000_0000_0000;
array[64497] <= 16'b0000_0000_0000_0000;
array[64498] <= 16'b0000_0000_0000_0000;
array[64499] <= 16'b0000_0000_0000_0000;
array[64500] <= 16'b0000_0000_0000_0000;
array[64501] <= 16'b0000_0000_0000_0000;
array[64502] <= 16'b0000_0000_0000_0000;
array[64503] <= 16'b0000_0000_0000_0000;
array[64504] <= 16'b0000_0000_0000_0000;
array[64505] <= 16'b0000_0000_0000_0000;
array[64506] <= 16'b0000_0000_0000_0000;
array[64507] <= 16'b0000_0000_0000_0000;
array[64508] <= 16'b0000_0000_0000_0000;
array[64509] <= 16'b0000_0000_0000_0000;
array[64510] <= 16'b0000_0000_0000_0000;
array[64511] <= 16'b0000_0000_0000_0000;
array[64512] <= 16'b0000_0000_0000_0000;
array[64513] <= 16'b0000_0000_0000_0000;
array[64514] <= 16'b0000_0000_0000_0000;
array[64515] <= 16'b0000_0000_0000_0000;
array[64516] <= 16'b0000_0000_0000_0000;
array[64517] <= 16'b0000_0000_0000_0000;
array[64518] <= 16'b0000_0000_0000_0000;
array[64519] <= 16'b0000_0000_0000_0000;
array[64520] <= 16'b0000_0000_0000_0000;
array[64521] <= 16'b0000_0000_0000_0000;
array[64522] <= 16'b0000_0000_0000_0000;
array[64523] <= 16'b0000_0000_0000_0000;
array[64524] <= 16'b0000_0000_0000_0000;
array[64525] <= 16'b0000_0000_0000_0000;
array[64526] <= 16'b0000_0000_0000_0000;
array[64527] <= 16'b0000_0000_0000_0000;
array[64528] <= 16'b0000_0000_0000_0000;
array[64529] <= 16'b0000_0000_0000_0000;
array[64530] <= 16'b0000_0000_0000_0000;
array[64531] <= 16'b0000_0000_0000_0000;
array[64532] <= 16'b0000_0000_0000_0000;
array[64533] <= 16'b0000_0000_0000_0000;
array[64534] <= 16'b0000_0000_0000_0000;
array[64535] <= 16'b0000_0000_0000_0000;
array[64536] <= 16'b0000_0000_0000_0000;
array[64537] <= 16'b0000_0000_0000_0000;
array[64538] <= 16'b0000_0000_0000_0000;
array[64539] <= 16'b0000_0000_0000_0000;
array[64540] <= 16'b0000_0000_0000_0000;
array[64541] <= 16'b0000_0000_0000_0000;
array[64542] <= 16'b0000_0000_0000_0000;
array[64543] <= 16'b0000_0000_0000_0000;
array[64544] <= 16'b0000_0000_0000_0000;
array[64545] <= 16'b0000_0000_0000_0000;
array[64546] <= 16'b0000_0000_0000_0000;
array[64547] <= 16'b0000_0000_0000_0000;
array[64548] <= 16'b0000_0000_0000_0000;
array[64549] <= 16'b0000_0000_0000_0000;
array[64550] <= 16'b0000_0000_0000_0000;
array[64551] <= 16'b0000_0000_0000_0000;
array[64552] <= 16'b0000_0000_0000_0000;
array[64553] <= 16'b0000_0000_0000_0000;
array[64554] <= 16'b0000_0000_0000_0000;
array[64555] <= 16'b0000_0000_0000_0000;
array[64556] <= 16'b0000_0000_0000_0000;
array[64557] <= 16'b0000_0000_0000_0000;
array[64558] <= 16'b0000_0000_0000_0000;
array[64559] <= 16'b0000_0000_0000_0000;
array[64560] <= 16'b0000_0000_0000_0000;
array[64561] <= 16'b0000_0000_0000_0000;
array[64562] <= 16'b0000_0000_0000_0000;
array[64563] <= 16'b0000_0000_0000_0000;
array[64564] <= 16'b0000_0000_0000_0000;
array[64565] <= 16'b0000_0000_0000_0000;
array[64566] <= 16'b0000_0000_0000_0000;
array[64567] <= 16'b0000_0000_0000_0000;
array[64568] <= 16'b0000_0000_0000_0000;
array[64569] <= 16'b0000_0000_0000_0000;
array[64570] <= 16'b0000_0000_0000_0000;
array[64571] <= 16'b0000_0000_0000_0000;
array[64572] <= 16'b0000_0000_0000_0000;
array[64573] <= 16'b0000_0000_0000_0000;
array[64574] <= 16'b0000_0000_0000_0000;
array[64575] <= 16'b0000_0000_0000_0000;
array[64576] <= 16'b0000_0000_0000_0000;
array[64577] <= 16'b0000_0000_0000_0000;
array[64578] <= 16'b0000_0000_0000_0000;
array[64579] <= 16'b0000_0000_0000_0000;
array[64580] <= 16'b0000_0000_0000_0000;
array[64581] <= 16'b0000_0000_0000_0000;
array[64582] <= 16'b0000_0000_0000_0000;
array[64583] <= 16'b0000_0000_0000_0000;
array[64584] <= 16'b0000_0000_0000_0000;
array[64585] <= 16'b0000_0000_0000_0000;
array[64586] <= 16'b0000_0000_0000_0000;
array[64587] <= 16'b0000_0000_0000_0000;
array[64588] <= 16'b0000_0000_0000_0000;
array[64589] <= 16'b0000_0000_0000_0000;
array[64590] <= 16'b0000_0000_0000_0000;
array[64591] <= 16'b0000_0000_0000_0000;
array[64592] <= 16'b0000_0000_0000_0000;
array[64593] <= 16'b0000_0000_0000_0000;
array[64594] <= 16'b0000_0000_0000_0000;
array[64595] <= 16'b0000_0000_0000_0000;
array[64596] <= 16'b0000_0000_0000_0000;
array[64597] <= 16'b0000_0000_0000_0000;
array[64598] <= 16'b0000_0000_0000_0000;
array[64599] <= 16'b0000_0000_0000_0000;
array[64600] <= 16'b0000_0000_0000_0000;
array[64601] <= 16'b0000_0000_0000_0000;
array[64602] <= 16'b0000_0000_0000_0000;
array[64603] <= 16'b0000_0000_0000_0000;
array[64604] <= 16'b0000_0000_0000_0000;
array[64605] <= 16'b0000_0000_0000_0000;
array[64606] <= 16'b0000_0000_0000_0000;
array[64607] <= 16'b0000_0000_0000_0000;
array[64608] <= 16'b0000_0000_0000_0000;
array[64609] <= 16'b0000_0000_0000_0000;
array[64610] <= 16'b0000_0000_0000_0000;
array[64611] <= 16'b0000_0000_0000_0000;
array[64612] <= 16'b0000_0000_0000_0000;
array[64613] <= 16'b0000_0000_0000_0000;
array[64614] <= 16'b0000_0000_0000_0000;
array[64615] <= 16'b0000_0000_0000_0000;
array[64616] <= 16'b0000_0000_0000_0000;
array[64617] <= 16'b0000_0000_0000_0000;
array[64618] <= 16'b0000_0000_0000_0000;
array[64619] <= 16'b0000_0000_0000_0000;
array[64620] <= 16'b0000_0000_0000_0000;
array[64621] <= 16'b0000_0000_0000_0000;
array[64622] <= 16'b0000_0000_0000_0000;
array[64623] <= 16'b0000_0000_0000_0000;
array[64624] <= 16'b0000_0000_0000_0000;
array[64625] <= 16'b0000_0000_0000_0000;
array[64626] <= 16'b0000_0000_0000_0000;
array[64627] <= 16'b0000_0000_0000_0000;
array[64628] <= 16'b0000_0000_0000_0000;
array[64629] <= 16'b0000_0000_0000_0000;
array[64630] <= 16'b0000_0000_0000_0000;
array[64631] <= 16'b0000_0000_0000_0000;
array[64632] <= 16'b0000_0000_0000_0000;
array[64633] <= 16'b0000_0000_0000_0000;
array[64634] <= 16'b0000_0000_0000_0000;
array[64635] <= 16'b0000_0000_0000_0000;
array[64636] <= 16'b0000_0000_0000_0000;
array[64637] <= 16'b0000_0000_0000_0000;
array[64638] <= 16'b0000_0000_0000_0000;
array[64639] <= 16'b0000_0000_0000_0000;
array[64640] <= 16'b0000_0000_0000_0000;
array[64641] <= 16'b0000_0000_0000_0000;
array[64642] <= 16'b0000_0000_0000_0000;
array[64643] <= 16'b0000_0000_0000_0000;
array[64644] <= 16'b0000_0000_0000_0000;
array[64645] <= 16'b0000_0000_0000_0000;
array[64646] <= 16'b0000_0000_0000_0000;
array[64647] <= 16'b0000_0000_0000_0000;
array[64648] <= 16'b0000_0000_0000_0000;
array[64649] <= 16'b0000_0000_0000_0000;
array[64650] <= 16'b0000_0000_0000_0000;
array[64651] <= 16'b0000_0000_0000_0000;
array[64652] <= 16'b0000_0000_0000_0000;
array[64653] <= 16'b0000_0000_0000_0000;
array[64654] <= 16'b0000_0000_0000_0000;
array[64655] <= 16'b0000_0000_0000_0000;
array[64656] <= 16'b0000_0000_0000_0000;
array[64657] <= 16'b0000_0000_0000_0000;
array[64658] <= 16'b0000_0000_0000_0000;
array[64659] <= 16'b0000_0000_0000_0000;
array[64660] <= 16'b0000_0000_0000_0000;
array[64661] <= 16'b0000_0000_0000_0000;
array[64662] <= 16'b0000_0000_0000_0000;
array[64663] <= 16'b0000_0000_0000_0000;
array[64664] <= 16'b0000_0000_0000_0000;
array[64665] <= 16'b0000_0000_0000_0000;
array[64666] <= 16'b0000_0000_0000_0000;
array[64667] <= 16'b0000_0000_0000_0000;
array[64668] <= 16'b0000_0000_0000_0000;
array[64669] <= 16'b0000_0000_0000_0000;
array[64670] <= 16'b0000_0000_0000_0000;
array[64671] <= 16'b0000_0000_0000_0000;
array[64672] <= 16'b0000_0000_0000_0000;
array[64673] <= 16'b0000_0000_0000_0000;
array[64674] <= 16'b0000_0000_0000_0000;
array[64675] <= 16'b0000_0000_0000_0000;
array[64676] <= 16'b0000_0000_0000_0000;
array[64677] <= 16'b0000_0000_0000_0000;
array[64678] <= 16'b0000_0000_0000_0000;
array[64679] <= 16'b0000_0000_0000_0000;
array[64680] <= 16'b0000_0000_0000_0000;
array[64681] <= 16'b0000_0000_0000_0000;
array[64682] <= 16'b0000_0000_0000_0000;
array[64683] <= 16'b0000_0000_0000_0000;
array[64684] <= 16'b0000_0000_0000_0000;
array[64685] <= 16'b0000_0000_0000_0000;
array[64686] <= 16'b0000_0000_0000_0000;
array[64687] <= 16'b0000_0000_0000_0000;
array[64688] <= 16'b0000_0000_0000_0000;
array[64689] <= 16'b0000_0000_0000_0000;
array[64690] <= 16'b0000_0000_0000_0000;
array[64691] <= 16'b0000_0000_0000_0000;
array[64692] <= 16'b0000_0000_0000_0000;
array[64693] <= 16'b0000_0000_0000_0000;
array[64694] <= 16'b0000_0000_0000_0000;
array[64695] <= 16'b0000_0000_0000_0000;
array[64696] <= 16'b0000_0000_0000_0000;
array[64697] <= 16'b0000_0000_0000_0000;
array[64698] <= 16'b0000_0000_0000_0000;
array[64699] <= 16'b0000_0000_0000_0000;
array[64700] <= 16'b0000_0000_0000_0000;
array[64701] <= 16'b0000_0000_0000_0000;
array[64702] <= 16'b0000_0000_0000_0000;
array[64703] <= 16'b0000_0000_0000_0000;
array[64704] <= 16'b0000_0000_0000_0000;
array[64705] <= 16'b0000_0000_0000_0000;
array[64706] <= 16'b0000_0000_0000_0000;
array[64707] <= 16'b0000_0000_0000_0000;
array[64708] <= 16'b0000_0000_0000_0000;
array[64709] <= 16'b0000_0000_0000_0000;
array[64710] <= 16'b0000_0000_0000_0000;
array[64711] <= 16'b0000_0000_0000_0000;
array[64712] <= 16'b0000_0000_0000_0000;
array[64713] <= 16'b0000_0000_0000_0000;
array[64714] <= 16'b0000_0000_0000_0000;
array[64715] <= 16'b0000_0000_0000_0000;
array[64716] <= 16'b0000_0000_0000_0000;
array[64717] <= 16'b0000_0000_0000_0000;
array[64718] <= 16'b0000_0000_0000_0000;
array[64719] <= 16'b0000_0000_0000_0000;
array[64720] <= 16'b0000_0000_0000_0000;
array[64721] <= 16'b0000_0000_0000_0000;
array[64722] <= 16'b0000_0000_0000_0000;
array[64723] <= 16'b0000_0000_0000_0000;
array[64724] <= 16'b0000_0000_0000_0000;
array[64725] <= 16'b0000_0000_0000_0000;
array[64726] <= 16'b0000_0000_0000_0000;
array[64727] <= 16'b0000_0000_0000_0000;
array[64728] <= 16'b0000_0000_0000_0000;
array[64729] <= 16'b0000_0000_0000_0000;
array[64730] <= 16'b0000_0000_0000_0000;
array[64731] <= 16'b0000_0000_0000_0000;
array[64732] <= 16'b0000_0000_0000_0000;
array[64733] <= 16'b0000_0000_0000_0000;
array[64734] <= 16'b0000_0000_0000_0000;
array[64735] <= 16'b0000_0000_0000_0000;
array[64736] <= 16'b0000_0000_0000_0000;
array[64737] <= 16'b0000_0000_0000_0000;
array[64738] <= 16'b0000_0000_0000_0000;
array[64739] <= 16'b0000_0000_0000_0000;
array[64740] <= 16'b0000_0000_0000_0000;
array[64741] <= 16'b0000_0000_0000_0000;
array[64742] <= 16'b0000_0000_0000_0000;
array[64743] <= 16'b0000_0000_0000_0000;
array[64744] <= 16'b0000_0000_0000_0000;
array[64745] <= 16'b0000_0000_0000_0000;
array[64746] <= 16'b0000_0000_0000_0000;
array[64747] <= 16'b0000_0000_0000_0000;
array[64748] <= 16'b0000_0000_0000_0000;
array[64749] <= 16'b0000_0000_0000_0000;
array[64750] <= 16'b0000_0000_0000_0000;
array[64751] <= 16'b0000_0000_0000_0000;
array[64752] <= 16'b0000_0000_0000_0000;
array[64753] <= 16'b0000_0000_0000_0000;
array[64754] <= 16'b0000_0000_0000_0000;
array[64755] <= 16'b0000_0000_0000_0000;
array[64756] <= 16'b0000_0000_0000_0000;
array[64757] <= 16'b0000_0000_0000_0000;
array[64758] <= 16'b0000_0000_0000_0000;
array[64759] <= 16'b0000_0000_0000_0000;
array[64760] <= 16'b0000_0000_0000_0000;
array[64761] <= 16'b0000_0000_0000_0000;
array[64762] <= 16'b0000_0000_0000_0000;
array[64763] <= 16'b0000_0000_0000_0000;
array[64764] <= 16'b0000_0000_0000_0000;
array[64765] <= 16'b0000_0000_0000_0000;
array[64766] <= 16'b0000_0000_0000_0000;
array[64767] <= 16'b0000_0000_0000_0000;
array[64768] <= 16'b0000_0000_0000_0000;
array[64769] <= 16'b0000_0000_0000_0000;
array[64770] <= 16'b0000_0000_0000_0000;
array[64771] <= 16'b0000_0000_0000_0000;
array[64772] <= 16'b0000_0000_0000_0000;
array[64773] <= 16'b0000_0000_0000_0000;
array[64774] <= 16'b0000_0000_0000_0000;
array[64775] <= 16'b0000_0000_0000_0000;
array[64776] <= 16'b0000_0000_0000_0000;
array[64777] <= 16'b0000_0000_0000_0000;
array[64778] <= 16'b0000_0000_0000_0000;
array[64779] <= 16'b0000_0000_0000_0000;
array[64780] <= 16'b0000_0000_0000_0000;
array[64781] <= 16'b0000_0000_0000_0000;
array[64782] <= 16'b0000_0000_0000_0000;
array[64783] <= 16'b0000_0000_0000_0000;
array[64784] <= 16'b0000_0000_0000_0000;
array[64785] <= 16'b0000_0000_0000_0000;
array[64786] <= 16'b0000_0000_0000_0000;
array[64787] <= 16'b0000_0000_0000_0000;
array[64788] <= 16'b0000_0000_0000_0000;
array[64789] <= 16'b0000_0000_0000_0000;
array[64790] <= 16'b0000_0000_0000_0000;
array[64791] <= 16'b0000_0000_0000_0000;
array[64792] <= 16'b0000_0000_0000_0000;
array[64793] <= 16'b0000_0000_0000_0000;
array[64794] <= 16'b0000_0000_0000_0000;
array[64795] <= 16'b0000_0000_0000_0000;
array[64796] <= 16'b0000_0000_0000_0000;
array[64797] <= 16'b0000_0000_0000_0000;
array[64798] <= 16'b0000_0000_0000_0000;
array[64799] <= 16'b0000_0000_0000_0000;
array[64800] <= 16'b0000_0000_0000_0000;
array[64801] <= 16'b0000_0000_0000_0000;
array[64802] <= 16'b0000_0000_0000_0000;
array[64803] <= 16'b0000_0000_0000_0000;
array[64804] <= 16'b0000_0000_0000_0000;
array[64805] <= 16'b0000_0000_0000_0000;
array[64806] <= 16'b0000_0000_0000_0000;
array[64807] <= 16'b0000_0000_0000_0000;
array[64808] <= 16'b0000_0000_0000_0000;
array[64809] <= 16'b0000_0000_0000_0000;
array[64810] <= 16'b0000_0000_0000_0000;
array[64811] <= 16'b0000_0000_0000_0000;
array[64812] <= 16'b0000_0000_0000_0000;
array[64813] <= 16'b0000_0000_0000_0000;
array[64814] <= 16'b0000_0000_0000_0000;
array[64815] <= 16'b0000_0000_0000_0000;
array[64816] <= 16'b0000_0000_0000_0000;
array[64817] <= 16'b0000_0000_0000_0000;
array[64818] <= 16'b0000_0000_0000_0000;
array[64819] <= 16'b0000_0000_0000_0000;
array[64820] <= 16'b0000_0000_0000_0000;
array[64821] <= 16'b0000_0000_0000_0000;
array[64822] <= 16'b0000_0000_0000_0000;
array[64823] <= 16'b0000_0000_0000_0000;
array[64824] <= 16'b0000_0000_0000_0000;
array[64825] <= 16'b0000_0000_0000_0000;
array[64826] <= 16'b0000_0000_0000_0000;
array[64827] <= 16'b0000_0000_0000_0000;
array[64828] <= 16'b0000_0000_0000_0000;
array[64829] <= 16'b0000_0000_0000_0000;
array[64830] <= 16'b0000_0000_0000_0000;
array[64831] <= 16'b0000_0000_0000_0000;
array[64832] <= 16'b0000_0000_0000_0000;
array[64833] <= 16'b0000_0000_0000_0000;
array[64834] <= 16'b0000_0000_0000_0000;
array[64835] <= 16'b0000_0000_0000_0000;
array[64836] <= 16'b0000_0000_0000_0000;
array[64837] <= 16'b0000_0000_0000_0000;
array[64838] <= 16'b0000_0000_0000_0000;
array[64839] <= 16'b0000_0000_0000_0000;
array[64840] <= 16'b0000_0000_0000_0000;
array[64841] <= 16'b0000_0000_0000_0000;
array[64842] <= 16'b0000_0000_0000_0000;
array[64843] <= 16'b0000_0000_0000_0000;
array[64844] <= 16'b0000_0000_0000_0000;
array[64845] <= 16'b0000_0000_0000_0000;
array[64846] <= 16'b0000_0000_0000_0000;
array[64847] <= 16'b0000_0000_0000_0000;
array[64848] <= 16'b0000_0000_0000_0000;
array[64849] <= 16'b0000_0000_0000_0000;
array[64850] <= 16'b0000_0000_0000_0000;
array[64851] <= 16'b0000_0000_0000_0000;
array[64852] <= 16'b0000_0000_0000_0000;
array[64853] <= 16'b0000_0000_0000_0000;
array[64854] <= 16'b0000_0000_0000_0000;
array[64855] <= 16'b0000_0000_0000_0000;
array[64856] <= 16'b0000_0000_0000_0000;
array[64857] <= 16'b0000_0000_0000_0000;
array[64858] <= 16'b0000_0000_0000_0000;
array[64859] <= 16'b0000_0000_0000_0000;
array[64860] <= 16'b0000_0000_0000_0000;
array[64861] <= 16'b0000_0000_0000_0000;
array[64862] <= 16'b0000_0000_0000_0000;
array[64863] <= 16'b0000_0000_0000_0000;
array[64864] <= 16'b0000_0000_0000_0000;
array[64865] <= 16'b0000_0000_0000_0000;
array[64866] <= 16'b0000_0000_0000_0000;
array[64867] <= 16'b0000_0000_0000_0000;
array[64868] <= 16'b0000_0000_0000_0000;
array[64869] <= 16'b0000_0000_0000_0000;
array[64870] <= 16'b0000_0000_0000_0000;
array[64871] <= 16'b0000_0000_0000_0000;
array[64872] <= 16'b0000_0000_0000_0000;
array[64873] <= 16'b0000_0000_0000_0000;
array[64874] <= 16'b0000_0000_0000_0000;
array[64875] <= 16'b0000_0000_0000_0000;
array[64876] <= 16'b0000_0000_0000_0000;
array[64877] <= 16'b0000_0000_0000_0000;
array[64878] <= 16'b0000_0000_0000_0000;
array[64879] <= 16'b0000_0000_0000_0000;
array[64880] <= 16'b0000_0000_0000_0000;
array[64881] <= 16'b0000_0000_0000_0000;
array[64882] <= 16'b0000_0000_0000_0000;
array[64883] <= 16'b0000_0000_0000_0000;
array[64884] <= 16'b0000_0000_0000_0000;
array[64885] <= 16'b0000_0000_0000_0000;
array[64886] <= 16'b0000_0000_0000_0000;
array[64887] <= 16'b0000_0000_0000_0000;
array[64888] <= 16'b0000_0000_0000_0000;
array[64889] <= 16'b0000_0000_0000_0000;
array[64890] <= 16'b0000_0000_0000_0000;
array[64891] <= 16'b0000_0000_0000_0000;
array[64892] <= 16'b0000_0000_0000_0000;
array[64893] <= 16'b0000_0000_0000_0000;
array[64894] <= 16'b0000_0000_0000_0000;
array[64895] <= 16'b0000_0000_0000_0000;
array[64896] <= 16'b0000_0000_0000_0000;
array[64897] <= 16'b0000_0000_0000_0000;
array[64898] <= 16'b0000_0000_0000_0000;
array[64899] <= 16'b0000_0000_0000_0000;
array[64900] <= 16'b0000_0000_0000_0000;
array[64901] <= 16'b0000_0000_0000_0000;
array[64902] <= 16'b0000_0000_0000_0000;
array[64903] <= 16'b0000_0000_0000_0000;
array[64904] <= 16'b0000_0000_0000_0000;
array[64905] <= 16'b0000_0000_0000_0000;
array[64906] <= 16'b0000_0000_0000_0000;
array[64907] <= 16'b0000_0000_0000_0000;
array[64908] <= 16'b0000_0000_0000_0000;
array[64909] <= 16'b0000_0000_0000_0000;
array[64910] <= 16'b0000_0000_0000_0000;
array[64911] <= 16'b0000_0000_0000_0000;
array[64912] <= 16'b0000_0000_0000_0000;
array[64913] <= 16'b0000_0000_0000_0000;
array[64914] <= 16'b0000_0000_0000_0000;
array[64915] <= 16'b0000_0000_0000_0000;
array[64916] <= 16'b0000_0000_0000_0000;
array[64917] <= 16'b0000_0000_0000_0000;
array[64918] <= 16'b0000_0000_0000_0000;
array[64919] <= 16'b0000_0000_0000_0000;
array[64920] <= 16'b0000_0000_0000_0000;
array[64921] <= 16'b0000_0000_0000_0000;
array[64922] <= 16'b0000_0000_0000_0000;
array[64923] <= 16'b0000_0000_0000_0000;
array[64924] <= 16'b0000_0000_0000_0000;
array[64925] <= 16'b0000_0000_0000_0000;
array[64926] <= 16'b0000_0000_0000_0000;
array[64927] <= 16'b0000_0000_0000_0000;
array[64928] <= 16'b0000_0000_0000_0000;
array[64929] <= 16'b0000_0000_0000_0000;
array[64930] <= 16'b0000_0000_0000_0000;
array[64931] <= 16'b0000_0000_0000_0000;
array[64932] <= 16'b0000_0000_0000_0000;
array[64933] <= 16'b0000_0000_0000_0000;
array[64934] <= 16'b0000_0000_0000_0000;
array[64935] <= 16'b0000_0000_0000_0000;
array[64936] <= 16'b0000_0000_0000_0000;
array[64937] <= 16'b0000_0000_0000_0000;
array[64938] <= 16'b0000_0000_0000_0000;
array[64939] <= 16'b0000_0000_0000_0000;
array[64940] <= 16'b0000_0000_0000_0000;
array[64941] <= 16'b0000_0000_0000_0000;
array[64942] <= 16'b0000_0000_0000_0000;
array[64943] <= 16'b0000_0000_0000_0000;
array[64944] <= 16'b0000_0000_0000_0000;
array[64945] <= 16'b0000_0000_0000_0000;
array[64946] <= 16'b0000_0000_0000_0000;
array[64947] <= 16'b0000_0000_0000_0000;
array[64948] <= 16'b0000_0000_0000_0000;
array[64949] <= 16'b0000_0000_0000_0000;
array[64950] <= 16'b0000_0000_0000_0000;
array[64951] <= 16'b0000_0000_0000_0000;
array[64952] <= 16'b0000_0000_0000_0000;
array[64953] <= 16'b0000_0000_0000_0000;
array[64954] <= 16'b0000_0000_0000_0000;
array[64955] <= 16'b0000_0000_0000_0000;
array[64956] <= 16'b0000_0000_0000_0000;
array[64957] <= 16'b0000_0000_0000_0000;
array[64958] <= 16'b0000_0000_0000_0000;
array[64959] <= 16'b0000_0000_0000_0000;
array[64960] <= 16'b0000_0000_0000_0000;
array[64961] <= 16'b0000_0000_0000_0000;
array[64962] <= 16'b0000_0000_0000_0000;
array[64963] <= 16'b0000_0000_0000_0000;
array[64964] <= 16'b0000_0000_0000_0000;
array[64965] <= 16'b0000_0000_0000_0000;
array[64966] <= 16'b0000_0000_0000_0000;
array[64967] <= 16'b0000_0000_0000_0000;
array[64968] <= 16'b0000_0000_0000_0000;
array[64969] <= 16'b0000_0000_0000_0000;
array[64970] <= 16'b0000_0000_0000_0000;
array[64971] <= 16'b0000_0000_0000_0000;
array[64972] <= 16'b0000_0000_0000_0000;
array[64973] <= 16'b0000_0000_0000_0000;
array[64974] <= 16'b0000_0000_0000_0000;
array[64975] <= 16'b0000_0000_0000_0000;
array[64976] <= 16'b0000_0000_0000_0000;
array[64977] <= 16'b0000_0000_0000_0000;
array[64978] <= 16'b0000_0000_0000_0000;
array[64979] <= 16'b0000_0000_0000_0000;
array[64980] <= 16'b0000_0000_0000_0000;
array[64981] <= 16'b0000_0000_0000_0000;
array[64982] <= 16'b0000_0000_0000_0000;
array[64983] <= 16'b0000_0000_0000_0000;
array[64984] <= 16'b0000_0000_0000_0000;
array[64985] <= 16'b0000_0000_0000_0000;
array[64986] <= 16'b0000_0000_0000_0000;
array[64987] <= 16'b0000_0000_0000_0000;
array[64988] <= 16'b0000_0000_0000_0000;
array[64989] <= 16'b0000_0000_0000_0000;
array[64990] <= 16'b0000_0000_0000_0000;
array[64991] <= 16'b0000_0000_0000_0000;
array[64992] <= 16'b0000_0000_0000_0000;
array[64993] <= 16'b0000_0000_0000_0000;
array[64994] <= 16'b0000_0000_0000_0000;
array[64995] <= 16'b0000_0000_0000_0000;
array[64996] <= 16'b0000_0000_0000_0000;
array[64997] <= 16'b0000_0000_0000_0000;
array[64998] <= 16'b0000_0000_0000_0000;
array[64999] <= 16'b0000_0000_0000_0000;
array[65000] <= 16'b0000_0000_0000_0000;
array[65001] <= 16'b0000_0000_0000_0000;
array[65002] <= 16'b0000_0000_0000_0000;
array[65003] <= 16'b0000_0000_0000_0000;
array[65004] <= 16'b0000_0000_0000_0000;
array[65005] <= 16'b0000_0000_0000_0000;
array[65006] <= 16'b0000_0000_0000_0000;
array[65007] <= 16'b0000_0000_0000_0000;
array[65008] <= 16'b0000_0000_0000_0000;
array[65009] <= 16'b0000_0000_0000_0000;
array[65010] <= 16'b0000_0000_0000_0000;
array[65011] <= 16'b0000_0000_0000_0000;
array[65012] <= 16'b0000_0000_0000_0000;
array[65013] <= 16'b0000_0000_0000_0000;
array[65014] <= 16'b0000_0000_0000_0000;
array[65015] <= 16'b0000_0000_0000_0000;
array[65016] <= 16'b0000_0000_0000_0000;
array[65017] <= 16'b0000_0000_0000_0000;
array[65018] <= 16'b0000_0000_0000_0000;
array[65019] <= 16'b0000_0000_0000_0000;
array[65020] <= 16'b0000_0000_0000_0000;
array[65021] <= 16'b0000_0000_0000_0000;
array[65022] <= 16'b0000_0000_0000_0000;
array[65023] <= 16'b0000_0000_0000_0000;
array[65024] <= 16'b0000_0000_0000_0000;
array[65025] <= 16'b0000_0000_0000_0000;
array[65026] <= 16'b0000_0000_0000_0000;
array[65027] <= 16'b0000_0000_0000_0000;
array[65028] <= 16'b0000_0000_0000_0000;
array[65029] <= 16'b0000_0000_0000_0000;
array[65030] <= 16'b0000_0000_0000_0000;
array[65031] <= 16'b0000_0000_0000_0000;
array[65032] <= 16'b0000_0000_0000_0000;
array[65033] <= 16'b0000_0000_0000_0000;
array[65034] <= 16'b0000_0000_0000_0000;
array[65035] <= 16'b0000_0000_0000_0000;
array[65036] <= 16'b0000_0000_0000_0000;
array[65037] <= 16'b0000_0000_0000_0000;
array[65038] <= 16'b0000_0000_0000_0000;
array[65039] <= 16'b0000_0000_0000_0000;
array[65040] <= 16'b0000_0000_0000_0000;
array[65041] <= 16'b0000_0000_0000_0000;
array[65042] <= 16'b0000_0000_0000_0000;
array[65043] <= 16'b0000_0000_0000_0000;
array[65044] <= 16'b0000_0000_0000_0000;
array[65045] <= 16'b0000_0000_0000_0000;
array[65046] <= 16'b0000_0000_0000_0000;
array[65047] <= 16'b0000_0000_0000_0000;
array[65048] <= 16'b0000_0000_0000_0000;
array[65049] <= 16'b0000_0000_0000_0000;
array[65050] <= 16'b0000_0000_0000_0000;
array[65051] <= 16'b0000_0000_0000_0000;
array[65052] <= 16'b0000_0000_0000_0000;
array[65053] <= 16'b0000_0000_0000_0000;
array[65054] <= 16'b0000_0000_0000_0000;
array[65055] <= 16'b0000_0000_0000_0000;
array[65056] <= 16'b0000_0000_0000_0000;
array[65057] <= 16'b0000_0000_0000_0000;
array[65058] <= 16'b0000_0000_0000_0000;
array[65059] <= 16'b0000_0000_0000_0000;
array[65060] <= 16'b0000_0000_0000_0000;
array[65061] <= 16'b0000_0000_0000_0000;
array[65062] <= 16'b0000_0000_0000_0000;
array[65063] <= 16'b0000_0000_0000_0000;
array[65064] <= 16'b0000_0000_0000_0000;
array[65065] <= 16'b0000_0000_0000_0000;
array[65066] <= 16'b0000_0000_0000_0000;
array[65067] <= 16'b0000_0000_0000_0000;
array[65068] <= 16'b0000_0000_0000_0000;
array[65069] <= 16'b0000_0000_0000_0000;
array[65070] <= 16'b0000_0000_0000_0000;
array[65071] <= 16'b0000_0000_0000_0000;
array[65072] <= 16'b0000_0000_0000_0000;
array[65073] <= 16'b0000_0000_0000_0000;
array[65074] <= 16'b0000_0000_0000_0000;
array[65075] <= 16'b0000_0000_0000_0000;
array[65076] <= 16'b0000_0000_0000_0000;
array[65077] <= 16'b0000_0000_0000_0000;
array[65078] <= 16'b0000_0000_0000_0000;
array[65079] <= 16'b0000_0000_0000_0000;
array[65080] <= 16'b0000_0000_0000_0000;
array[65081] <= 16'b0000_0000_0000_0000;
array[65082] <= 16'b0000_0000_0000_0000;
array[65083] <= 16'b0000_0000_0000_0000;
array[65084] <= 16'b0000_0000_0000_0000;
array[65085] <= 16'b0000_0000_0000_0000;
array[65086] <= 16'b0000_0000_0000_0000;
array[65087] <= 16'b0000_0000_0000_0000;
array[65088] <= 16'b0000_0000_0000_0000;
array[65089] <= 16'b0000_0000_0000_0000;
array[65090] <= 16'b0000_0000_0000_0000;
array[65091] <= 16'b0000_0000_0000_0000;
array[65092] <= 16'b0000_0000_0000_0000;
array[65093] <= 16'b0000_0000_0000_0000;
array[65094] <= 16'b0000_0000_0000_0000;
array[65095] <= 16'b0000_0000_0000_0000;
array[65096] <= 16'b0000_0000_0000_0000;
array[65097] <= 16'b0000_0000_0000_0000;
array[65098] <= 16'b0000_0000_0000_0000;
array[65099] <= 16'b0000_0000_0000_0000;
array[65100] <= 16'b0000_0000_0000_0000;
array[65101] <= 16'b0000_0000_0000_0000;
array[65102] <= 16'b0000_0000_0000_0000;
array[65103] <= 16'b0000_0000_0000_0000;
array[65104] <= 16'b0000_0000_0000_0000;
array[65105] <= 16'b0000_0000_0000_0000;
array[65106] <= 16'b0000_0000_0000_0000;
array[65107] <= 16'b0000_0000_0000_0000;
array[65108] <= 16'b0000_0000_0000_0000;
array[65109] <= 16'b0000_0000_0000_0000;
array[65110] <= 16'b0000_0000_0000_0000;
array[65111] <= 16'b0000_0000_0000_0000;
array[65112] <= 16'b0000_0000_0000_0000;
array[65113] <= 16'b0000_0000_0000_0000;
array[65114] <= 16'b0000_0000_0000_0000;
array[65115] <= 16'b0000_0000_0000_0000;
array[65116] <= 16'b0000_0000_0000_0000;
array[65117] <= 16'b0000_0000_0000_0000;
array[65118] <= 16'b0000_0000_0000_0000;
array[65119] <= 16'b0000_0000_0000_0000;
array[65120] <= 16'b0000_0000_0000_0000;
array[65121] <= 16'b0000_0000_0000_0000;
array[65122] <= 16'b0000_0000_0000_0000;
array[65123] <= 16'b0000_0000_0000_0000;
array[65124] <= 16'b0000_0000_0000_0000;
array[65125] <= 16'b0000_0000_0000_0000;
array[65126] <= 16'b0000_0000_0000_0000;
array[65127] <= 16'b0000_0000_0000_0000;
array[65128] <= 16'b0000_0000_0000_0000;
array[65129] <= 16'b0000_0000_0000_0000;
array[65130] <= 16'b0000_0000_0000_0000;
array[65131] <= 16'b0000_0000_0000_0000;
array[65132] <= 16'b0000_0000_0000_0000;
array[65133] <= 16'b0000_0000_0000_0000;
array[65134] <= 16'b0000_0000_0000_0000;
array[65135] <= 16'b0000_0000_0000_0000;
array[65136] <= 16'b0000_0000_0000_0000;
array[65137] <= 16'b0000_0000_0000_0000;
array[65138] <= 16'b0000_0000_0000_0000;
array[65139] <= 16'b0000_0000_0000_0000;
array[65140] <= 16'b0000_0000_0000_0000;
array[65141] <= 16'b0000_0000_0000_0000;
array[65142] <= 16'b0000_0000_0000_0000;
array[65143] <= 16'b0000_0000_0000_0000;
array[65144] <= 16'b0000_0000_0000_0000;
array[65145] <= 16'b0000_0000_0000_0000;
array[65146] <= 16'b0000_0000_0000_0000;
array[65147] <= 16'b0000_0000_0000_0000;
array[65148] <= 16'b0000_0000_0000_0000;
array[65149] <= 16'b0000_0000_0000_0000;
array[65150] <= 16'b0000_0000_0000_0000;
array[65151] <= 16'b0000_0000_0000_0000;
array[65152] <= 16'b0000_0000_0000_0000;
array[65153] <= 16'b0000_0000_0000_0000;
array[65154] <= 16'b0000_0000_0000_0000;
array[65155] <= 16'b0000_0000_0000_0000;
array[65156] <= 16'b0000_0000_0000_0000;
array[65157] <= 16'b0000_0000_0000_0000;
array[65158] <= 16'b0000_0000_0000_0000;
array[65159] <= 16'b0000_0000_0000_0000;
array[65160] <= 16'b0000_0000_0000_0000;
array[65161] <= 16'b0000_0000_0000_0000;
array[65162] <= 16'b0000_0000_0000_0000;
array[65163] <= 16'b0000_0000_0000_0000;
array[65164] <= 16'b0000_0000_0000_0000;
array[65165] <= 16'b0000_0000_0000_0000;
array[65166] <= 16'b0000_0000_0000_0000;
array[65167] <= 16'b0000_0000_0000_0000;
array[65168] <= 16'b0000_0000_0000_0000;
array[65169] <= 16'b0000_0000_0000_0000;
array[65170] <= 16'b0000_0000_0000_0000;
array[65171] <= 16'b0000_0000_0000_0000;
array[65172] <= 16'b0000_0000_0000_0000;
array[65173] <= 16'b0000_0000_0000_0000;
array[65174] <= 16'b0000_0000_0000_0000;
array[65175] <= 16'b0000_0000_0000_0000;
array[65176] <= 16'b0000_0000_0000_0000;
array[65177] <= 16'b0000_0000_0000_0000;
array[65178] <= 16'b0000_0000_0000_0000;
array[65179] <= 16'b0000_0000_0000_0000;
array[65180] <= 16'b0000_0000_0000_0000;
array[65181] <= 16'b0000_0000_0000_0000;
array[65182] <= 16'b0000_0000_0000_0000;
array[65183] <= 16'b0000_0000_0000_0000;
array[65184] <= 16'b0000_0000_0000_0000;
array[65185] <= 16'b0000_0000_0000_0000;
array[65186] <= 16'b0000_0000_0000_0000;
array[65187] <= 16'b0000_0000_0000_0000;
array[65188] <= 16'b0000_0000_0000_0000;
array[65189] <= 16'b0000_0000_0000_0000;
array[65190] <= 16'b0000_0000_0000_0000;
array[65191] <= 16'b0000_0000_0000_0000;
array[65192] <= 16'b0000_0000_0000_0000;
array[65193] <= 16'b0000_0000_0000_0000;
array[65194] <= 16'b0000_0000_0000_0000;
array[65195] <= 16'b0000_0000_0000_0000;
array[65196] <= 16'b0000_0000_0000_0000;
array[65197] <= 16'b0000_0000_0000_0000;
array[65198] <= 16'b0000_0000_0000_0000;
array[65199] <= 16'b0000_0000_0000_0000;
array[65200] <= 16'b0000_0000_0000_0000;
array[65201] <= 16'b0000_0000_0000_0000;
array[65202] <= 16'b0000_0000_0000_0000;
array[65203] <= 16'b0000_0000_0000_0000;
array[65204] <= 16'b0000_0000_0000_0000;
array[65205] <= 16'b0000_0000_0000_0000;
array[65206] <= 16'b0000_0000_0000_0000;
array[65207] <= 16'b0000_0000_0000_0000;
array[65208] <= 16'b0000_0000_0000_0000;
array[65209] <= 16'b0000_0000_0000_0000;
array[65210] <= 16'b0000_0000_0000_0000;
array[65211] <= 16'b0000_0000_0000_0000;
array[65212] <= 16'b0000_0000_0000_0000;
array[65213] <= 16'b0000_0000_0000_0000;
array[65214] <= 16'b0000_0000_0000_0000;
array[65215] <= 16'b0000_0000_0000_0000;
array[65216] <= 16'b0000_0000_0000_0000;
array[65217] <= 16'b0000_0000_0000_0000;
array[65218] <= 16'b0000_0000_0000_0000;
array[65219] <= 16'b0000_0000_0000_0000;
array[65220] <= 16'b0000_0000_0000_0000;
array[65221] <= 16'b0000_0000_0000_0000;
array[65222] <= 16'b0000_0000_0000_0000;
array[65223] <= 16'b0000_0000_0000_0000;
array[65224] <= 16'b0000_0000_0000_0000;
array[65225] <= 16'b0000_0000_0000_0000;
array[65226] <= 16'b0000_0000_0000_0000;
array[65227] <= 16'b0000_0000_0000_0000;
array[65228] <= 16'b0000_0000_0000_0000;
array[65229] <= 16'b0000_0000_0000_0000;
array[65230] <= 16'b0000_0000_0000_0000;
array[65231] <= 16'b0000_0000_0000_0000;
array[65232] <= 16'b0000_0000_0000_0000;
array[65233] <= 16'b0000_0000_0000_0000;
array[65234] <= 16'b0000_0000_0000_0000;
array[65235] <= 16'b0000_0000_0000_0000;
array[65236] <= 16'b0000_0000_0000_0000;
array[65237] <= 16'b0000_0000_0000_0000;
array[65238] <= 16'b0000_0000_0000_0000;
array[65239] <= 16'b0000_0000_0000_0000;
array[65240] <= 16'b0000_0000_0000_0000;
array[65241] <= 16'b0000_0000_0000_0000;
array[65242] <= 16'b0000_0000_0000_0000;
array[65243] <= 16'b0000_0000_0000_0000;
array[65244] <= 16'b0000_0000_0000_0000;
array[65245] <= 16'b0000_0000_0000_0000;
array[65246] <= 16'b0000_0000_0000_0000;
array[65247] <= 16'b0000_0000_0000_0000;
array[65248] <= 16'b0000_0000_0000_0000;
array[65249] <= 16'b0000_0000_0000_0000;
array[65250] <= 16'b0000_0000_0000_0000;
array[65251] <= 16'b0000_0000_0000_0000;
array[65252] <= 16'b0000_0000_0000_0000;
array[65253] <= 16'b0000_0000_0000_0000;
array[65254] <= 16'b0000_0000_0000_0000;
array[65255] <= 16'b0000_0000_0000_0000;
array[65256] <= 16'b0000_0000_0000_0000;
array[65257] <= 16'b0000_0000_0000_0000;
array[65258] <= 16'b0000_0000_0000_0000;
array[65259] <= 16'b0000_0000_0000_0000;
array[65260] <= 16'b0000_0000_0000_0000;
array[65261] <= 16'b0000_0000_0000_0000;
array[65262] <= 16'b0000_0000_0000_0000;
array[65263] <= 16'b0000_0000_0000_0000;
array[65264] <= 16'b0000_0000_0000_0000;
array[65265] <= 16'b0000_0000_0000_0000;
array[65266] <= 16'b0000_0000_0000_0000;
array[65267] <= 16'b0000_0000_0000_0000;
array[65268] <= 16'b0000_0000_0000_0000;
array[65269] <= 16'b0000_0000_0000_0000;
array[65270] <= 16'b0000_0000_0000_0000;
array[65271] <= 16'b0000_0000_0000_0000;
array[65272] <= 16'b0000_0000_0000_0000;
array[65273] <= 16'b0000_0000_0000_0000;
array[65274] <= 16'b0000_0000_0000_0000;
array[65275] <= 16'b0000_0000_0000_0000;
array[65276] <= 16'b0000_0000_0000_0000;
array[65277] <= 16'b0000_0000_0000_0000;
array[65278] <= 16'b0000_0000_0000_0000;
array[65279] <= 16'b0000_0000_0000_0000;
array[65280] <= 16'b0000_0000_0000_0000;
array[65281] <= 16'b0000_0000_0000_0000;
array[65282] <= 16'b0000_0000_0000_0000;
array[65283] <= 16'b0000_0000_0000_0000;
array[65284] <= 16'b0000_0000_0000_0000;
array[65285] <= 16'b0000_0000_0000_0000;
array[65286] <= 16'b0000_0000_0000_0000;
array[65287] <= 16'b0000_0000_0000_0000;
array[65288] <= 16'b0000_0000_0000_0000;
array[65289] <= 16'b0000_0000_0000_0000;
array[65290] <= 16'b0000_0000_0000_0000;
array[65291] <= 16'b0000_0000_0000_0000;
array[65292] <= 16'b0000_0000_0000_0000;
array[65293] <= 16'b0000_0000_0000_0000;
array[65294] <= 16'b0000_0000_0000_0000;
array[65295] <= 16'b0000_0000_0000_0000;
array[65296] <= 16'b0000_0000_0000_0000;
array[65297] <= 16'b0000_0000_0000_0000;
array[65298] <= 16'b0000_0000_0000_0000;
array[65299] <= 16'b0000_0000_0000_0000;
array[65300] <= 16'b0000_0000_0000_0000;
array[65301] <= 16'b0000_0000_0000_0000;
array[65302] <= 16'b0000_0000_0000_0000;
array[65303] <= 16'b0000_0000_0000_0000;
array[65304] <= 16'b0000_0000_0000_0000;
array[65305] <= 16'b0000_0000_0000_0000;
array[65306] <= 16'b0000_0000_0000_0000;
array[65307] <= 16'b0000_0000_0000_0000;
array[65308] <= 16'b0000_0000_0000_0000;
array[65309] <= 16'b0000_0000_0000_0000;
array[65310] <= 16'b0000_0000_0000_0000;
array[65311] <= 16'b0000_0000_0000_0000;
array[65312] <= 16'b0000_0000_0000_0000;
array[65313] <= 16'b0000_0000_0000_0000;
array[65314] <= 16'b0000_0000_0000_0000;
array[65315] <= 16'b0000_0000_0000_0000;
array[65316] <= 16'b0000_0000_0000_0000;
array[65317] <= 16'b0000_0000_0000_0000;
array[65318] <= 16'b0000_0000_0000_0000;
array[65319] <= 16'b0000_0000_0000_0000;
array[65320] <= 16'b0000_0000_0000_0000;
array[65321] <= 16'b0000_0000_0000_0000;
array[65322] <= 16'b0000_0000_0000_0000;
array[65323] <= 16'b0000_0000_0000_0000;
array[65324] <= 16'b0000_0000_0000_0000;
array[65325] <= 16'b0000_0000_0000_0000;
array[65326] <= 16'b0000_0000_0000_0000;
array[65327] <= 16'b0000_0000_0000_0000;
array[65328] <= 16'b0000_0000_0000_0000;
array[65329] <= 16'b0000_0000_0000_0000;
array[65330] <= 16'b0000_0000_0000_0000;
array[65331] <= 16'b0000_0000_0000_0000;
array[65332] <= 16'b0000_0000_0000_0000;
array[65333] <= 16'b0000_0000_0000_0000;
array[65334] <= 16'b0000_0000_0000_0000;
array[65335] <= 16'b0000_0000_0000_0000;
array[65336] <= 16'b0000_0000_0000_0000;
array[65337] <= 16'b0000_0000_0000_0000;
array[65338] <= 16'b0000_0000_0000_0000;
array[65339] <= 16'b0000_0000_0000_0000;
array[65340] <= 16'b0000_0000_0000_0000;
array[65341] <= 16'b0000_0000_0000_0000;
array[65342] <= 16'b0000_0000_0000_0000;
array[65343] <= 16'b0000_0000_0000_0000;
array[65344] <= 16'b0000_0000_0000_0000;
array[65345] <= 16'b0000_0000_0000_0000;
array[65346] <= 16'b0000_0000_0000_0000;
array[65347] <= 16'b0000_0000_0000_0000;
array[65348] <= 16'b0000_0000_0000_0000;
array[65349] <= 16'b0000_0000_0000_0000;
array[65350] <= 16'b0000_0000_0000_0000;
array[65351] <= 16'b0000_0000_0000_0000;
array[65352] <= 16'b0000_0000_0000_0000;
array[65353] <= 16'b0000_0000_0000_0000;
array[65354] <= 16'b0000_0000_0000_0000;
array[65355] <= 16'b0000_0000_0000_0000;
array[65356] <= 16'b0000_0000_0000_0000;
array[65357] <= 16'b0000_0000_0000_0000;
array[65358] <= 16'b0000_0000_0000_0000;
array[65359] <= 16'b0000_0000_0000_0000;
array[65360] <= 16'b0000_0000_0000_0000;
array[65361] <= 16'b0000_0000_0000_0000;
array[65362] <= 16'b0000_0000_0000_0000;
array[65363] <= 16'b0000_0000_0000_0000;
array[65364] <= 16'b0000_0000_0000_0000;
array[65365] <= 16'b0000_0000_0000_0000;
array[65366] <= 16'b0000_0000_0000_0000;
array[65367] <= 16'b0000_0000_0000_0000;
array[65368] <= 16'b0000_0000_0000_0000;
array[65369] <= 16'b0000_0000_0000_0000;
array[65370] <= 16'b0000_0000_0000_0000;
array[65371] <= 16'b0000_0000_0000_0000;
array[65372] <= 16'b0000_0000_0000_0000;
array[65373] <= 16'b0000_0000_0000_0000;
array[65374] <= 16'b0000_0000_0000_0000;
array[65375] <= 16'b0000_0000_0000_0000;
array[65376] <= 16'b0000_0000_0000_0000;
array[65377] <= 16'b0000_0000_0000_0000;
array[65378] <= 16'b0000_0000_0000_0000;
array[65379] <= 16'b0000_0000_0000_0000;
array[65380] <= 16'b0000_0000_0000_0000;
array[65381] <= 16'b0000_0000_0000_0000;
array[65382] <= 16'b0000_0000_0000_0000;
array[65383] <= 16'b0000_0000_0000_0000;
array[65384] <= 16'b0000_0000_0000_0000;
array[65385] <= 16'b0000_0000_0000_0000;
array[65386] <= 16'b0000_0000_0000_0000;
array[65387] <= 16'b0000_0000_0000_0000;
array[65388] <= 16'b0000_0000_0000_0000;
array[65389] <= 16'b0000_0000_0000_0000;
array[65390] <= 16'b0000_0000_0000_0000;
array[65391] <= 16'b0000_0000_0000_0000;
array[65392] <= 16'b0000_0000_0000_0000;
array[65393] <= 16'b0000_0000_0000_0000;
array[65394] <= 16'b0000_0000_0000_0000;
array[65395] <= 16'b0000_0000_0000_0000;
array[65396] <= 16'b0000_0000_0000_0000;
array[65397] <= 16'b0000_0000_0000_0000;
array[65398] <= 16'b0000_0000_0000_0000;
array[65399] <= 16'b0000_0000_0000_0000;
array[65400] <= 16'b0000_0000_0000_0000;
array[65401] <= 16'b0000_0000_0000_0000;
array[65402] <= 16'b0000_0000_0000_0000;
array[65403] <= 16'b0000_0000_0000_0000;
array[65404] <= 16'b0000_0000_0000_0000;
array[65405] <= 16'b0000_0000_0000_0000;
array[65406] <= 16'b0000_0000_0000_0000;
array[65407] <= 16'b0000_0000_0000_0000;
array[65408] <= 16'b0000_0000_0000_0000;
array[65409] <= 16'b0000_0000_0000_0000;
array[65410] <= 16'b0000_0000_0000_0000;
array[65411] <= 16'b0000_0000_0000_0000;
array[65412] <= 16'b0000_0000_0000_0000;
array[65413] <= 16'b0000_0000_0000_0000;
array[65414] <= 16'b0000_0000_0000_0000;
array[65415] <= 16'b0000_0000_0000_0000;
array[65416] <= 16'b0000_0000_0000_0000;
array[65417] <= 16'b0000_0000_0000_0000;
array[65418] <= 16'b0000_0000_0000_0000;
array[65419] <= 16'b0000_0000_0000_0000;
array[65420] <= 16'b0000_0000_0000_0000;
array[65421] <= 16'b0000_0000_0000_0000;
array[65422] <= 16'b0000_0000_0000_0000;
array[65423] <= 16'b0000_0000_0000_0000;
array[65424] <= 16'b0000_0000_0000_0000;
array[65425] <= 16'b0000_0000_0000_0000;
array[65426] <= 16'b0000_0000_0000_0000;
array[65427] <= 16'b0000_0000_0000_0000;
array[65428] <= 16'b0000_0000_0000_0000;
array[65429] <= 16'b0000_0000_0000_0000;
array[65430] <= 16'b0000_0000_0000_0000;
array[65431] <= 16'b0000_0000_0000_0000;
array[65432] <= 16'b0000_0000_0000_0000;
array[65433] <= 16'b0000_0000_0000_0000;
array[65434] <= 16'b0000_0000_0000_0000;
array[65435] <= 16'b0000_0000_0000_0000;
array[65436] <= 16'b0000_0000_0000_0000;
array[65437] <= 16'b0000_0000_0000_0000;
array[65438] <= 16'b0000_0000_0000_0000;
array[65439] <= 16'b0000_0000_0000_0000;
array[65440] <= 16'b0000_0000_0000_0000;
array[65441] <= 16'b0000_0000_0000_0000;
array[65442] <= 16'b0000_0000_0000_0000;
array[65443] <= 16'b0000_0000_0000_0000;
array[65444] <= 16'b0000_0000_0000_0000;
array[65445] <= 16'b0000_0000_0000_0000;
array[65446] <= 16'b0000_0000_0000_0000;
array[65447] <= 16'b0000_0000_0000_0000;
array[65448] <= 16'b0000_0000_0000_0000;
array[65449] <= 16'b0000_0000_0000_0000;
array[65450] <= 16'b0000_0000_0000_0000;
array[65451] <= 16'b0000_0000_0000_0000;
array[65452] <= 16'b0000_0000_0000_0000;
array[65453] <= 16'b0000_0000_0000_0000;
array[65454] <= 16'b0000_0000_0000_0000;
array[65455] <= 16'b0000_0000_0000_0000;
array[65456] <= 16'b0000_0000_0000_0000;
array[65457] <= 16'b0000_0000_0000_0000;
array[65458] <= 16'b0000_0000_0000_0000;
array[65459] <= 16'b0000_0000_0000_0000;
array[65460] <= 16'b0000_0000_0000_0000;
array[65461] <= 16'b0000_0000_0000_0000;
array[65462] <= 16'b0000_0000_0000_0000;
array[65463] <= 16'b0000_0000_0000_0000;
array[65464] <= 16'b0000_0000_0000_0000;
array[65465] <= 16'b0000_0000_0000_0000;
array[65466] <= 16'b0000_0000_0000_0000;
array[65467] <= 16'b0000_0000_0000_0000;
array[65468] <= 16'b0000_0000_0000_0000;
array[65469] <= 16'b0000_0000_0000_0000;
array[65470] <= 16'b0000_0000_0000_0000;
array[65471] <= 16'b0000_0000_0000_0000;
array[65472] <= 16'b0000_0000_0000_0000;
array[65473] <= 16'b0000_0000_0000_0000;
array[65474] <= 16'b0000_0000_0000_0000;
array[65475] <= 16'b0000_0000_0000_0000;
array[65476] <= 16'b0000_0000_0000_0000;
array[65477] <= 16'b0000_0000_0000_0000;
array[65478] <= 16'b0000_0000_0000_0000;
array[65479] <= 16'b0000_0000_0000_0000;
array[65480] <= 16'b0000_0000_0000_0000;
array[65481] <= 16'b0000_0000_0000_0000;
array[65482] <= 16'b0000_0000_0000_0000;
array[65483] <= 16'b0000_0000_0000_0000;
array[65484] <= 16'b0000_0000_0000_0000;
array[65485] <= 16'b0000_0000_0000_0000;
array[65486] <= 16'b0000_0000_0000_0000;
array[65487] <= 16'b0000_0000_0000_0000;
array[65488] <= 16'b0000_0000_0000_0000;
array[65489] <= 16'b0000_0000_0000_0000;
array[65490] <= 16'b0000_0000_0000_0000;
array[65491] <= 16'b0000_0000_0000_0000;
array[65492] <= 16'b0000_0000_0000_0000;
array[65493] <= 16'b0000_0000_0000_0000;
array[65494] <= 16'b0000_0000_0000_0000;
array[65495] <= 16'b0000_0000_0000_0000;
array[65496] <= 16'b0000_0000_0000_0000;
array[65497] <= 16'b0000_0000_0000_0000;
array[65498] <= 16'b0000_0000_0000_0000;
array[65499] <= 16'b0000_0000_0000_0000;
array[65500] <= 16'b0000_0000_0000_0000;
array[65501] <= 16'b0000_0000_0000_0000;
array[65502] <= 16'b0000_0000_0000_0000;
array[65503] <= 16'b0000_0000_0000_0000;
array[65504] <= 16'b0000_0000_0000_0000;
array[65505] <= 16'b0000_0000_0000_0000;
array[65506] <= 16'b0000_0000_0000_0000;
array[65507] <= 16'b0000_0000_0000_0000;
array[65508] <= 16'b0000_0000_0000_0000;
array[65509] <= 16'b0000_0000_0000_0000;
array[65510] <= 16'b0000_0000_0000_0000;
array[65511] <= 16'b0000_0000_0000_0000;
array[65512] <= 16'b0000_0000_0000_0000;
array[65513] <= 16'b0000_0000_0000_0000;
array[65514] <= 16'b0000_0000_0000_0000;
array[65515] <= 16'b0000_0000_0000_0000;
array[65516] <= 16'b0000_0000_0000_0000;
array[65517] <= 16'b0000_0000_0000_0000;
array[65518] <= 16'b0000_0000_0000_0000;
array[65519] <= 16'b0000_0000_0000_0000;
array[65520] <= 16'b0000_0000_0000_0000;
array[65521] <= 16'b0000_0000_0000_0000;
array[65522] <= 16'b0000_0000_0000_0000;
array[65523] <= 16'b0000_0000_0000_0000;
array[65524] <= 16'b0000_0000_0000_0000;
array[65525] <= 16'b0000_0000_0000_0000;
array[65526] <= 16'b0000_0000_0000_0000;
array[65527] <= 16'b0000_0000_0000_0000;
array[65528] <= 16'b0000_0000_0000_0000;
array[65529] <= 16'b0000_0000_0000_0000;
array[65530] <= 16'b0000_0000_0000_0000;
array[65531] <= 16'b0000_0000_0000_0000;
array[65532] <= 16'b0000_0000_0000_0000;
array[65533] <= 16'b0000_0000_0000_0000;
array[65534] <= 16'b0000_0000_0000_0000;
array[65535] <= 16'b0000_0000_0000_0000;
state=0;
end
else if(start & ~state)
begin
ad_t=address;
rwn_t=rwn;
data_t=data_in;
counter=address[1:0];
state=1;
end
else if(|counter && state)
counter=counter-1;
else if(state)
begin
if(rwn_t)
data_out=array[ad_t];
else
array[ad_t]=data_t;
state=0;
end
end
endmodule
